/* modified netlist. Source: module sbox in file Designs/AESSbox/lookup/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 34 time(s)  */

module sbox_HPC1_ClockGating_d3 (SI_s0, clk, SI_s1, SI_s2, SI_s3, Fresh, rst, SO_s0, SO_s1, SO_s2, SO_s3, Synch);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input [7:0] SI_s2 ;
    input [7:0] SI_s3 ;
    input rst ;
    input [8679:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    output [7:0] SO_s2 ;
    output [7:0] SO_s3 ;
    output Synch ;
    wire N169 ;
    wire N277 ;
    wire N379 ;
    wire N470 ;
    wire N563 ;
    wire N639 ;
    wire N723 ;
    wire N789 ;
    wire n1922 ;
    wire n1923 ;
    wire n1924 ;
    wire n1925 ;
    wire n1926 ;
    wire n1927 ;
    wire n1928 ;
    wire n1929 ;
    wire n1930 ;
    wire n1931 ;
    wire n1932 ;
    wire n1933 ;
    wire n1934 ;
    wire n1935 ;
    wire n1936 ;
    wire n1937 ;
    wire n1938 ;
    wire n1939 ;
    wire n1940 ;
    wire n1941 ;
    wire n1942 ;
    wire n1943 ;
    wire n1944 ;
    wire n1945 ;
    wire n1946 ;
    wire n1947 ;
    wire n1948 ;
    wire n1949 ;
    wire n1950 ;
    wire n1951 ;
    wire n1952 ;
    wire n1953 ;
    wire n1954 ;
    wire n1955 ;
    wire n1956 ;
    wire n1957 ;
    wire n1958 ;
    wire n1959 ;
    wire n1960 ;
    wire n1961 ;
    wire n1962 ;
    wire n1963 ;
    wire n1964 ;
    wire n1965 ;
    wire n1966 ;
    wire n1967 ;
    wire n1968 ;
    wire n1969 ;
    wire n1970 ;
    wire n1971 ;
    wire n1972 ;
    wire n1973 ;
    wire n1974 ;
    wire n1975 ;
    wire n1976 ;
    wire n1977 ;
    wire n1978 ;
    wire n1979 ;
    wire n1980 ;
    wire n1981 ;
    wire n1982 ;
    wire n1983 ;
    wire n1984 ;
    wire n1985 ;
    wire n1986 ;
    wire n1987 ;
    wire n1988 ;
    wire n1989 ;
    wire n1990 ;
    wire n1991 ;
    wire n1992 ;
    wire n1993 ;
    wire n1994 ;
    wire n1995 ;
    wire n1996 ;
    wire n1997 ;
    wire n1998 ;
    wire n1999 ;
    wire n2000 ;
    wire n2001 ;
    wire n2002 ;
    wire n2003 ;
    wire n2004 ;
    wire n2005 ;
    wire n2006 ;
    wire n2007 ;
    wire n2008 ;
    wire n2009 ;
    wire n2010 ;
    wire n2011 ;
    wire n2012 ;
    wire n2013 ;
    wire n2014 ;
    wire n2015 ;
    wire n2016 ;
    wire n2017 ;
    wire n2018 ;
    wire n2019 ;
    wire n2020 ;
    wire n2021 ;
    wire n2022 ;
    wire n2023 ;
    wire n2024 ;
    wire n2025 ;
    wire n2026 ;
    wire n2027 ;
    wire n2028 ;
    wire n2029 ;
    wire n2030 ;
    wire n2031 ;
    wire n2032 ;
    wire n2033 ;
    wire n2034 ;
    wire n2035 ;
    wire n2036 ;
    wire n2037 ;
    wire n2038 ;
    wire n2039 ;
    wire n2040 ;
    wire n2041 ;
    wire n2042 ;
    wire n2043 ;
    wire n2044 ;
    wire n2045 ;
    wire n2046 ;
    wire n2047 ;
    wire n2048 ;
    wire n2049 ;
    wire n2050 ;
    wire n2051 ;
    wire n2052 ;
    wire n2053 ;
    wire n2054 ;
    wire n2055 ;
    wire n2056 ;
    wire n2057 ;
    wire n2058 ;
    wire n2059 ;
    wire n2060 ;
    wire n2061 ;
    wire n2062 ;
    wire n2063 ;
    wire n2064 ;
    wire n2065 ;
    wire n2066 ;
    wire n2067 ;
    wire n2068 ;
    wire n2069 ;
    wire n2070 ;
    wire n2071 ;
    wire n2072 ;
    wire n2073 ;
    wire n2074 ;
    wire n2075 ;
    wire n2076 ;
    wire n2077 ;
    wire n2078 ;
    wire n2079 ;
    wire n2080 ;
    wire n2081 ;
    wire n2082 ;
    wire n2083 ;
    wire n2084 ;
    wire n2085 ;
    wire n2086 ;
    wire n2087 ;
    wire n2088 ;
    wire n2089 ;
    wire n2090 ;
    wire n2091 ;
    wire n2092 ;
    wire n2093 ;
    wire n2094 ;
    wire n2095 ;
    wire n2096 ;
    wire n2097 ;
    wire n2098 ;
    wire n2099 ;
    wire n2100 ;
    wire n2101 ;
    wire n2102 ;
    wire n2103 ;
    wire n2104 ;
    wire n2105 ;
    wire n2106 ;
    wire n2107 ;
    wire n2108 ;
    wire n2109 ;
    wire n2110 ;
    wire n2111 ;
    wire n2112 ;
    wire n2113 ;
    wire n2114 ;
    wire n2115 ;
    wire n2116 ;
    wire n2117 ;
    wire n2118 ;
    wire n2119 ;
    wire n2120 ;
    wire n2121 ;
    wire n2122 ;
    wire n2123 ;
    wire n2124 ;
    wire n2125 ;
    wire n2126 ;
    wire n2127 ;
    wire n2128 ;
    wire n2129 ;
    wire n2130 ;
    wire n2131 ;
    wire n2132 ;
    wire n2133 ;
    wire n2134 ;
    wire n2135 ;
    wire n2136 ;
    wire n2137 ;
    wire n2138 ;
    wire n2139 ;
    wire n2140 ;
    wire n2141 ;
    wire n2142 ;
    wire n2143 ;
    wire n2144 ;
    wire n2145 ;
    wire n2146 ;
    wire n2147 ;
    wire n2148 ;
    wire n2149 ;
    wire n2150 ;
    wire n2151 ;
    wire n2152 ;
    wire n2153 ;
    wire n2154 ;
    wire n2155 ;
    wire n2156 ;
    wire n2157 ;
    wire n2158 ;
    wire n2159 ;
    wire n2160 ;
    wire n2161 ;
    wire n2162 ;
    wire n2163 ;
    wire n2164 ;
    wire n2165 ;
    wire n2166 ;
    wire n2167 ;
    wire n2168 ;
    wire n2169 ;
    wire n2170 ;
    wire n2171 ;
    wire n2172 ;
    wire n2173 ;
    wire n2174 ;
    wire n2175 ;
    wire n2176 ;
    wire n2177 ;
    wire n2178 ;
    wire n2179 ;
    wire n2180 ;
    wire n2181 ;
    wire n2182 ;
    wire n2183 ;
    wire n2184 ;
    wire n2185 ;
    wire n2186 ;
    wire n2187 ;
    wire n2188 ;
    wire n2189 ;
    wire n2190 ;
    wire n2191 ;
    wire n2192 ;
    wire n2193 ;
    wire n2194 ;
    wire n2195 ;
    wire n2196 ;
    wire n2197 ;
    wire n2198 ;
    wire n2199 ;
    wire n2200 ;
    wire n2201 ;
    wire n2202 ;
    wire n2203 ;
    wire n2204 ;
    wire n2205 ;
    wire n2206 ;
    wire n2207 ;
    wire n2208 ;
    wire n2209 ;
    wire n2210 ;
    wire n2211 ;
    wire n2212 ;
    wire n2213 ;
    wire n2214 ;
    wire n2215 ;
    wire n2216 ;
    wire n2217 ;
    wire n2218 ;
    wire n2219 ;
    wire n2220 ;
    wire n2221 ;
    wire n2222 ;
    wire n2223 ;
    wire n2224 ;
    wire n2225 ;
    wire n2226 ;
    wire n2227 ;
    wire n2228 ;
    wire n2229 ;
    wire n2230 ;
    wire n2231 ;
    wire n2232 ;
    wire n2233 ;
    wire n2234 ;
    wire n2235 ;
    wire n2236 ;
    wire n2237 ;
    wire n2238 ;
    wire n2239 ;
    wire n2240 ;
    wire n2241 ;
    wire n2242 ;
    wire n2243 ;
    wire n2244 ;
    wire n2245 ;
    wire n2246 ;
    wire n2247 ;
    wire n2248 ;
    wire n2249 ;
    wire n2250 ;
    wire n2251 ;
    wire n2252 ;
    wire n2253 ;
    wire n2254 ;
    wire n2255 ;
    wire n2256 ;
    wire n2257 ;
    wire n2258 ;
    wire n2259 ;
    wire n2260 ;
    wire n2261 ;
    wire n2262 ;
    wire n2263 ;
    wire n2264 ;
    wire n2265 ;
    wire n2266 ;
    wire n2267 ;
    wire n2268 ;
    wire n2269 ;
    wire n2270 ;
    wire n2271 ;
    wire n2272 ;
    wire n2273 ;
    wire n2274 ;
    wire n2275 ;
    wire n2276 ;
    wire n2277 ;
    wire n2278 ;
    wire n2279 ;
    wire n2280 ;
    wire n2281 ;
    wire n2282 ;
    wire n2283 ;
    wire n2284 ;
    wire n2285 ;
    wire n2286 ;
    wire n2287 ;
    wire n2288 ;
    wire n2289 ;
    wire n2290 ;
    wire n2291 ;
    wire n2292 ;
    wire n2293 ;
    wire n2294 ;
    wire n2295 ;
    wire n2296 ;
    wire n2297 ;
    wire n2298 ;
    wire n2299 ;
    wire n2300 ;
    wire n2301 ;
    wire n2302 ;
    wire n2303 ;
    wire n2304 ;
    wire n2305 ;
    wire n2306 ;
    wire n2307 ;
    wire n2308 ;
    wire n2309 ;
    wire n2310 ;
    wire n2311 ;
    wire n2312 ;
    wire n2313 ;
    wire n2314 ;
    wire n2315 ;
    wire n2316 ;
    wire n2317 ;
    wire n2318 ;
    wire n2319 ;
    wire n2320 ;
    wire n2321 ;
    wire n2322 ;
    wire n2323 ;
    wire n2324 ;
    wire n2325 ;
    wire n2326 ;
    wire n2327 ;
    wire n2328 ;
    wire n2329 ;
    wire n2330 ;
    wire n2331 ;
    wire n2332 ;
    wire n2333 ;
    wire n2334 ;
    wire n2335 ;
    wire n2336 ;
    wire n2337 ;
    wire n2338 ;
    wire n2339 ;
    wire n2340 ;
    wire n2341 ;
    wire n2342 ;
    wire n2343 ;
    wire n2344 ;
    wire n2345 ;
    wire n2346 ;
    wire n2347 ;
    wire n2348 ;
    wire n2349 ;
    wire n2350 ;
    wire n2351 ;
    wire n2352 ;
    wire n2353 ;
    wire n2354 ;
    wire n2355 ;
    wire n2356 ;
    wire n2357 ;
    wire n2358 ;
    wire n2359 ;
    wire n2360 ;
    wire n2361 ;
    wire n2362 ;
    wire n2363 ;
    wire n2364 ;
    wire n2365 ;
    wire n2366 ;
    wire n2367 ;
    wire n2368 ;
    wire n2369 ;
    wire n2370 ;
    wire n2371 ;
    wire n2372 ;
    wire n2373 ;
    wire n2374 ;
    wire n2375 ;
    wire n2376 ;
    wire n2377 ;
    wire n2378 ;
    wire n2379 ;
    wire n2380 ;
    wire n2381 ;
    wire n2382 ;
    wire n2383 ;
    wire n2384 ;
    wire n2385 ;
    wire n2386 ;
    wire n2387 ;
    wire n2388 ;
    wire n2389 ;
    wire n2390 ;
    wire n2391 ;
    wire n2392 ;
    wire n2393 ;
    wire n2394 ;
    wire n2395 ;
    wire n2396 ;
    wire n2397 ;
    wire n2398 ;
    wire n2399 ;
    wire n2400 ;
    wire n2401 ;
    wire n2402 ;
    wire n2403 ;
    wire n2404 ;
    wire n2405 ;
    wire n2406 ;
    wire n2407 ;
    wire n2408 ;
    wire n2409 ;
    wire n2410 ;
    wire n2411 ;
    wire n2412 ;
    wire n2413 ;
    wire n2414 ;
    wire n2415 ;
    wire n2416 ;
    wire n2417 ;
    wire n2418 ;
    wire n2419 ;
    wire n2420 ;
    wire n2421 ;
    wire n2422 ;
    wire n2423 ;
    wire n2424 ;
    wire n2425 ;
    wire n2426 ;
    wire n2427 ;
    wire n2428 ;
    wire n2429 ;
    wire n2430 ;
    wire n2431 ;
    wire n2432 ;
    wire n2433 ;
    wire n2434 ;
    wire n2435 ;
    wire n2436 ;
    wire n2437 ;
    wire n2438 ;
    wire n2439 ;
    wire n2440 ;
    wire n2441 ;
    wire n2442 ;
    wire n2443 ;
    wire n2444 ;
    wire n2445 ;
    wire n2446 ;
    wire n2447 ;
    wire n2448 ;
    wire n2449 ;
    wire n2450 ;
    wire n2451 ;
    wire n2452 ;
    wire n2453 ;
    wire n2454 ;
    wire n2455 ;
    wire n2456 ;
    wire n2457 ;
    wire n2458 ;
    wire n2459 ;
    wire n2460 ;
    wire n2461 ;
    wire n2462 ;
    wire n2463 ;
    wire n2464 ;
    wire n2465 ;
    wire n2466 ;
    wire n2467 ;
    wire n2468 ;
    wire n2469 ;
    wire n2470 ;
    wire n2471 ;
    wire n2472 ;
    wire n2473 ;
    wire n2474 ;
    wire n2475 ;
    wire n2476 ;
    wire n2477 ;
    wire n2478 ;
    wire n2479 ;
    wire n2480 ;
    wire n2481 ;
    wire n2482 ;
    wire n2483 ;
    wire n2484 ;
    wire n2485 ;
    wire n2486 ;
    wire n2487 ;
    wire n2488 ;
    wire n2489 ;
    wire n2490 ;
    wire n2491 ;
    wire n2492 ;
    wire n2493 ;
    wire n2494 ;
    wire n2495 ;
    wire n2496 ;
    wire n2497 ;
    wire n2498 ;
    wire n2499 ;
    wire n2500 ;
    wire n2501 ;
    wire n2502 ;
    wire n2503 ;
    wire n2504 ;
    wire n2505 ;
    wire n2506 ;
    wire n2507 ;
    wire n2508 ;
    wire n2509 ;
    wire n2510 ;
    wire n2511 ;
    wire n2512 ;
    wire n2513 ;
    wire n2514 ;
    wire n2515 ;
    wire n2516 ;
    wire n2517 ;
    wire n2518 ;
    wire n2519 ;
    wire n2520 ;
    wire n2521 ;
    wire n2522 ;
    wire n2523 ;
    wire n2524 ;
    wire n2525 ;
    wire n2526 ;
    wire n2527 ;
    wire n2528 ;
    wire n2529 ;
    wire n2530 ;
    wire n2531 ;
    wire n2532 ;
    wire n2533 ;
    wire n2534 ;
    wire n2535 ;
    wire n2536 ;
    wire n2537 ;
    wire n2538 ;
    wire n2539 ;
    wire n2540 ;
    wire n2541 ;
    wire n2542 ;
    wire n2543 ;
    wire n2544 ;
    wire n2545 ;
    wire n2546 ;
    wire n2547 ;
    wire n2548 ;
    wire n2549 ;
    wire n2550 ;
    wire n2551 ;
    wire n2552 ;
    wire n2553 ;
    wire n2554 ;
    wire n2555 ;
    wire n2556 ;
    wire n2557 ;
    wire n2558 ;
    wire n2559 ;
    wire n2560 ;
    wire n2561 ;
    wire n2562 ;
    wire n2563 ;
    wire n2564 ;
    wire n2565 ;
    wire n2566 ;
    wire n2567 ;
    wire n2568 ;
    wire n2569 ;
    wire n2570 ;
    wire n2571 ;
    wire n2572 ;
    wire n2573 ;
    wire n2574 ;
    wire n2575 ;
    wire n2576 ;
    wire n2577 ;
    wire n2578 ;
    wire n2579 ;
    wire n2580 ;
    wire n2581 ;
    wire n2582 ;
    wire n2583 ;
    wire n2584 ;
    wire n2585 ;
    wire n2586 ;
    wire n2587 ;
    wire n2588 ;
    wire n2589 ;
    wire n2590 ;
    wire n2591 ;
    wire n2592 ;
    wire n2593 ;
    wire n2594 ;
    wire n2595 ;
    wire n2596 ;
    wire n2597 ;
    wire n2598 ;
    wire n2599 ;
    wire n2600 ;
    wire n2601 ;
    wire n2602 ;
    wire n2603 ;
    wire n2604 ;
    wire n2605 ;
    wire n2606 ;
    wire n2607 ;
    wire n2608 ;
    wire n2609 ;
    wire n2610 ;
    wire n2611 ;
    wire n2612 ;
    wire n2613 ;
    wire n2614 ;
    wire n2615 ;
    wire n2616 ;
    wire n2617 ;
    wire n2618 ;
    wire n2619 ;
    wire n2620 ;
    wire n2621 ;
    wire n2622 ;
    wire n2623 ;
    wire n2624 ;
    wire n2625 ;
    wire n2626 ;
    wire n2627 ;
    wire n2628 ;
    wire n2629 ;
    wire n2630 ;
    wire n2631 ;
    wire n2632 ;
    wire n2633 ;
    wire n2634 ;
    wire n2635 ;
    wire n2636 ;
    wire n2637 ;
    wire n2638 ;
    wire n2639 ;
    wire n2640 ;
    wire n2641 ;
    wire n2642 ;
    wire n2643 ;
    wire n2644 ;
    wire n2645 ;
    wire n2646 ;
    wire n2647 ;
    wire n2648 ;
    wire n2649 ;
    wire n2650 ;
    wire n2651 ;
    wire n2652 ;
    wire n2653 ;
    wire n2654 ;
    wire n2655 ;
    wire n2656 ;
    wire n2657 ;
    wire n2658 ;
    wire n2659 ;
    wire n2660 ;
    wire n2661 ;
    wire n2662 ;
    wire n2663 ;
    wire n2664 ;
    wire n2665 ;
    wire n2666 ;
    wire n2667 ;
    wire n2668 ;
    wire n2669 ;
    wire n2670 ;
    wire n2671 ;
    wire n2672 ;
    wire n2673 ;
    wire n2674 ;
    wire n2675 ;
    wire n2676 ;
    wire n2677 ;
    wire n2678 ;
    wire n2679 ;
    wire n2680 ;
    wire n2681 ;
    wire n2682 ;
    wire n2683 ;
    wire n2684 ;
    wire n2685 ;
    wire n2686 ;
    wire n2687 ;
    wire n2688 ;
    wire n2689 ;
    wire n2690 ;
    wire n2691 ;
    wire n2692 ;
    wire n2693 ;
    wire n2694 ;
    wire n2695 ;
    wire n2696 ;
    wire n2697 ;
    wire n2698 ;
    wire n2699 ;
    wire n2700 ;
    wire n2701 ;
    wire n2702 ;
    wire n2703 ;
    wire n2704 ;
    wire n2705 ;
    wire n2706 ;
    wire n2707 ;
    wire n2708 ;
    wire n2709 ;
    wire n2710 ;
    wire n2711 ;
    wire n2712 ;
    wire n2713 ;
    wire n2714 ;
    wire n2715 ;
    wire n2716 ;
    wire n2717 ;
    wire n2718 ;
    wire n2719 ;
    wire n2720 ;
    wire n2721 ;
    wire n2722 ;
    wire n2723 ;
    wire n2724 ;
    wire n2725 ;
    wire n2726 ;
    wire n2727 ;
    wire n2728 ;
    wire n2729 ;
    wire n2730 ;
    wire n2731 ;
    wire n2732 ;
    wire n2733 ;
    wire n2734 ;
    wire n2735 ;
    wire n2736 ;
    wire n2737 ;
    wire n2738 ;
    wire n2739 ;
    wire n2740 ;
    wire n2741 ;
    wire n2742 ;
    wire n2743 ;
    wire n2744 ;
    wire n2745 ;
    wire n2746 ;
    wire n2747 ;
    wire n2748 ;
    wire n2749 ;
    wire n2750 ;
    wire n2751 ;
    wire n2752 ;
    wire n2753 ;
    wire n2754 ;
    wire n2755 ;
    wire n2756 ;
    wire n2757 ;
    wire n2758 ;
    wire n2759 ;
    wire n2760 ;
    wire n2761 ;
    wire n2762 ;
    wire n2763 ;
    wire n2764 ;
    wire n2765 ;
    wire n2766 ;
    wire n2767 ;
    wire n2768 ;
    wire n2769 ;
    wire n2770 ;
    wire n2771 ;
    wire n2772 ;
    wire n2773 ;
    wire n2774 ;
    wire n2775 ;
    wire n2776 ;
    wire n2777 ;
    wire n2778 ;
    wire n2779 ;
    wire n2780 ;
    wire n2781 ;
    wire n2782 ;
    wire n2783 ;
    wire n2784 ;
    wire n2785 ;
    wire n2786 ;
    wire n2787 ;
    wire n2788 ;
    wire n2789 ;
    wire n2790 ;
    wire n2791 ;
    wire n2792 ;
    wire n2793 ;
    wire n2794 ;
    wire n2795 ;
    wire n2796 ;
    wire n2797 ;
    wire n2798 ;
    wire n2799 ;
    wire n2800 ;
    wire n2801 ;
    wire n2802 ;
    wire n2803 ;
    wire n2804 ;
    wire n2805 ;
    wire n2806 ;
    wire n2807 ;
    wire n2808 ;
    wire n2809 ;
    wire n2810 ;
    wire n2811 ;
    wire n2812 ;
    wire n2813 ;
    wire n2814 ;
    wire n2815 ;
    wire n2816 ;
    wire n2817 ;
    wire n2818 ;
    wire n2819 ;
    wire n2820 ;
    wire n2821 ;
    wire n2822 ;
    wire n2823 ;
    wire n2824 ;
    wire n2825 ;
    wire n2826 ;
    wire n2827 ;
    wire n2828 ;
    wire n2829 ;
    wire n2830 ;
    wire n2831 ;
    wire n2832 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_946 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_952 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_958 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_992 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire clk_gated ;

    /* cells in depth 0 */
    not_masked #(.security_order(3), .pipeline(0)) U1938 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1939 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1940 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1941 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1942 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1944 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1945 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1946 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}) ) ;
    ClockGatingController #(35) ClockGatingInst ( .clk ( clk ), .rst ( rst ), .GatedClk ( clk_gated ), .Synch ( Synch ) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1937 ( .ina ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .inb ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .clk ( clk ), .rnd ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .outt ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1943 ( .a ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, new_AGEMA_signal_1125, n2624}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1947 ( .ina ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .outt ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1948 ( .ina ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}), .inb ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .clk ( clk ), .rnd ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .outt ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1949 ( .ina ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .outt ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1950 ( .ina ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .inb ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .clk ( clk ), .rnd ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .outt ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1951 ( .a ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .b ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1952 ( .ina ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .outt ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1953 ( .a ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}), .b ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2640}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1955 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .outt ({new_AGEMA_signal_1040, new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2699}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1956 ( .a ({new_AGEMA_signal_1040, new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2699}), .b ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1957 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .rnd ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .outt ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1958 ( .a ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .b ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1961 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .outt ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1962 ( .a ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .b ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1963 ( .ina ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .inb ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .clk ( clk ), .rnd ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .outt ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1965 ( .ina ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .inb ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .clk ( clk ), .rnd ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .outt ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1966 ( .a ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .b ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1969 ( .ina ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .inb ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .rnd ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .outt ({new_AGEMA_signal_1055, new_AGEMA_signal_1054, new_AGEMA_signal_1053, n2073}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1970 ( .a ({new_AGEMA_signal_1055, new_AGEMA_signal_1054, new_AGEMA_signal_1053, n2073}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1971 ( .ina ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .outt ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1972 ( .ina ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .inb ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130]}), .outt ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1973 ( .a ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}), .b ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1975 ( .ina ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .inb ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .outt ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1976 ( .a ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .b ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1978 ( .ina ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .inb ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .clk ( clk ), .rnd ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .outt ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1979 ( .a ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .b ({new_AGEMA_signal_1214, new_AGEMA_signal_1213, new_AGEMA_signal_1212, n2541}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1984 ( .ina ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .inb ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .rnd ({Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .outt ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1985 ( .a ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .b ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, n2086}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1987 ( .ina ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .inb ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .rnd ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170]}), .outt ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2600}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1990 ( .ina ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .outt ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, new_AGEMA_signal_1071, n2538}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1991 ( .a ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, new_AGEMA_signal_1071, n2538}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1995 ( .ina ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .inb ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190]}), .outt ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, new_AGEMA_signal_1005, n2595}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1996 ( .a ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, new_AGEMA_signal_1005, n2595}), .b ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1999 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200]}), .outt ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2000 ( .a ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}), .b ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, n2577}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2004 ( .ina ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .inb ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .rnd ({Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .outt ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2400}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2008 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220]}), .outt ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, n2785}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2009 ( .a ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, n2785}), .b ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2013 ( .ina ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .inb ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230]}), .outt ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2014 ( .a ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .b ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2017 ( .ina ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .inb ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .rnd ({Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .outt ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2018 ( .a ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}), .b ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, n2174}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2020 ( .ina ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250]}), .outt ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2021 ( .a ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .b ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2493}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2025 ( .ina ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260]}), .outt ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, n2587}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2028 ( .a ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .b ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2570}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2029 ( .ina ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .inb ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .outt ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2035 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280]}), .outt ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2036 ( .a ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .b ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2038 ( .a ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .b ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, new_AGEMA_signal_1101, n2739}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2044 ( .ina ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}), .inb ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .clk ( clk ), .rnd ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290]}), .outt ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2045 ( .ina ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .inb ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .rnd ({Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .outt ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2046 ( .a ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}), .b ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2052 ( .ina ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .inb ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .rnd ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310]}), .outt ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2452}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2055 ( .a ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .b ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2068 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .outt ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2772}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2070 ( .ina ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .outt ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2071 ( .a ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2074 ( .a ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2400}), .b ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2313}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2089 ( .ina ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .inb ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .clk ( clk ), .rnd ({Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340]}), .outt ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2395}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2090 ( .a ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2395}), .b ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2094 ( .ina ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350]}), .outt ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, new_AGEMA_signal_1017, n2779}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2096 ( .ina ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .inb ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .rnd ({Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .outt ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, new_AGEMA_signal_1125, n2624}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2097 ( .ina ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .inb ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .rnd ({Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370]}), .outt ({new_AGEMA_signal_1022, new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2242}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2100 ( .ina ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .rnd ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384], Fresh[383], Fresh[382], Fresh[381], Fresh[380]}), .outt ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2356}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2119 ( .a ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2772}), .b ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2122 ( .ina ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .outt ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2131 ( .a ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .b ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, n2828}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2133 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400]}), .outt ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2134 ( .a ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}), .b ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2679}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2138 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .clk ( clk ), .rnd ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410]}), .outt ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2139 ( .a ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}), .b ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, n2809}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2150 ( .a ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .b ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, new_AGEMA_signal_1320, n2709}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2163 ( .ina ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .inb ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .clk ( clk ), .rnd ({Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .outt ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2401}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2211 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432], Fresh[431], Fresh[430]}), .outt ({new_AGEMA_signal_1148, new_AGEMA_signal_1147, new_AGEMA_signal_1146, n2061}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2232 ( .ina ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .inb ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .rnd ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440]}), .outt ({new_AGEMA_signal_1151, new_AGEMA_signal_1150, new_AGEMA_signal_1149, n2721}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2276 ( .ina ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .inb ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .clk ( clk ), .rnd ({Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .outt ({new_AGEMA_signal_1154, new_AGEMA_signal_1153, new_AGEMA_signal_1152, n2298}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2278 ( .a ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2401}), .b ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, new_AGEMA_signal_1356, n2118}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2307 ( .ina ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462], Fresh[461], Fresh[460]}), .outt ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, new_AGEMA_signal_1155, n2346}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2341 ( .ina ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .rnd ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470]}), .outt ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, new_AGEMA_signal_1161, n2430}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2383 ( .ina ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .inb ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .rnd ({Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .outt ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, n2712}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2402 ( .ina ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .rnd ({Fresh[499], Fresh[498], Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490]}), .outt ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, n2777}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2615 ( .ina ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}), .clk ( clk ), .rnd ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500]}), .outt ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, new_AGEMA_signal_1173, n2463}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2627 ( .ina ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .inb ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[519], Fresh[518], Fresh[517], Fresh[516], Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .outt ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, new_AGEMA_signal_1176, n2474}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1954 ( .ina ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .inb ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2640}), .clk ( clk ), .rnd ({Fresh[529], Fresh[528], Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520]}), .outt ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, new_AGEMA_signal_1497, n2575}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1959 ( .ina ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}), .inb ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .clk ( clk ), .rnd ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530]}), .outt ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, new_AGEMA_signal_1500, n1962}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1964 ( .ina ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .inb ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}), .clk ( clk ), .rnd ({Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .outt ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, new_AGEMA_signal_1503, n1922}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1974 ( .ina ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .inb ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .rnd ({Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552], Fresh[551], Fresh[550]}), .outt ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, new_AGEMA_signal_1206, n2755}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1977 ( .ina ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}), .inb ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .clk ( clk ), .rnd ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564], Fresh[563], Fresh[562], Fresh[561], Fresh[560]}), .outt ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, new_AGEMA_signal_1506, n1926}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1980 ( .ina ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .inb ({new_AGEMA_signal_1214, new_AGEMA_signal_1213, new_AGEMA_signal_1212, n2541}), .clk ( clk ), .rnd ({Fresh[579], Fresh[578], Fresh[577], Fresh[576], Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .outt ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, new_AGEMA_signal_1509, n1925}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1986 ( .ina ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, n2086}), .inb ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}), .clk ( clk ), .rnd ({Fresh[589], Fresh[588], Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580]}), .outt ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, new_AGEMA_signal_1512, n2151}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1988 ( .ina ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .inb ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2600}), .clk ( clk ), .rnd ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592], Fresh[591], Fresh[590]}), .outt ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2631}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U1989 ( .a ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2631}), .b ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, n2734}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1992 ( .ina ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .inb ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .clk ( clk ), .rnd ({Fresh[609], Fresh[608], Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .outt ({new_AGEMA_signal_1520, new_AGEMA_signal_1519, new_AGEMA_signal_1518, n2763}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1997 ( .ina ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .inb ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .clk ( clk ), .rnd ({Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612], Fresh[611], Fresh[610]}), .outt ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, new_AGEMA_signal_1224, n1930}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2005 ( .ina ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2400}), .inb ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .clk ( clk ), .rnd ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624], Fresh[623], Fresh[622], Fresh[621], Fresh[620]}), .outt ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2006 ( .a ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}), .b ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2010 ( .ina ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .inb ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .clk ( clk ), .rnd ({Fresh[639], Fresh[638], Fresh[637], Fresh[636], Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .outt ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, new_AGEMA_signal_1524, n1937}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2022 ( .ina ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .inb ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2493}), .clk ( clk ), .rnd ({Fresh[649], Fresh[648], Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640]}), .outt ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, new_AGEMA_signal_1242, n1942}) ) ;
    or_HPC1 #(.security_order(3), .pipeline(0)) U2026 ( .ina ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, n2587}), .inb ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .clk ( clk ), .rnd ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650]}), .outt ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, new_AGEMA_signal_1245, n2676}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2030 ( .ina ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .inb ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}), .clk ( clk ), .rnd ({Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .outt ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, new_AGEMA_signal_1533, n1944}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2037 ( .ina ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .inb ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .clk ( clk ), .rnd ({Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672], Fresh[671], Fresh[670]}), .outt ({new_AGEMA_signal_1538, new_AGEMA_signal_1537, new_AGEMA_signal_1536, n1950}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2039 ( .ina ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .inb ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, new_AGEMA_signal_1101, n2739}), .clk ( clk ), .rnd ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684], Fresh[683], Fresh[682], Fresh[681], Fresh[680]}), .outt ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, new_AGEMA_signal_1254, n1949}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2042 ( .ina ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .inb ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2600}), .clk ( clk ), .rnd ({Fresh[699], Fresh[698], Fresh[697], Fresh[696], Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .outt ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, n2677}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2043 ( .a ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, n2677}), .b ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1539, n2662}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2047 ( .ina ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .inb ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .clk ( clk ), .rnd ({Fresh[709], Fresh[708], Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702], Fresh[701], Fresh[700]}), .outt ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2053 ( .ina ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .inb ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2452}), .clk ( clk ), .rnd ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710]}), .outt ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, new_AGEMA_signal_1263, n1957}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2056 ( .ina ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .inb ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2600}), .clk ( clk ), .rnd ({Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .outt ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, new_AGEMA_signal_1542, n2088}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2062 ( .ina ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .inb ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .clk ( clk ), .rnd ({Fresh[739], Fresh[738], Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732], Fresh[731], Fresh[730]}), .outt ({new_AGEMA_signal_1115, new_AGEMA_signal_1114, new_AGEMA_signal_1113, n1964}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2063 ( .ina ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .clk ( clk ), .rnd ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744], Fresh[743], Fresh[742], Fresh[741], Fresh[740]}), .outt ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, n2736}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2069 ( .ina ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2772}), .inb ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[759], Fresh[758], Fresh[757], Fresh[756], Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .outt ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, new_AGEMA_signal_1272, n2673}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2072 ( .ina ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .inb ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .clk ( clk ), .rnd ({Fresh[769], Fresh[768], Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760]}), .outt ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2073 ( .a ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, n2720}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2075 ( .ina ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2313}), .inb ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .clk ( clk ), .rnd ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770]}), .outt ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, new_AGEMA_signal_1551, n2412}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2076 ( .a ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, new_AGEMA_signal_1551, n2412}), .b ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2079 ( .ina ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .inb ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}), .clk ( clk ), .rnd ({Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .outt ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, n2571}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2080 ( .a ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, n2571}), .b ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2505}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2081 ( .ina ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .inb ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}), .clk ( clk ), .rnd ({Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792], Fresh[791], Fresh[790]}), .outt ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2083 ( .ina ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .inb ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804], Fresh[803], Fresh[802], Fresh[801], Fresh[800]}), .outt ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, new_AGEMA_signal_1557, n2359}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2086 ( .ina ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .inb ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .clk ( clk ), .rnd ({Fresh[819], Fresh[818], Fresh[817], Fresh[816], Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .outt ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, n2101}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2087 ( .a ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, n2101}), .b ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2625}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2091 ( .ina ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .inb ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .clk ( clk ), .rnd ({Fresh[829], Fresh[828], Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820]}), .outt ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, n2190}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2095 ( .ina ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, new_AGEMA_signal_1101, n2739}), .inb ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, new_AGEMA_signal_1017, n2779}), .clk ( clk ), .rnd ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832], Fresh[831], Fresh[830]}), .outt ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, new_AGEMA_signal_1296, n1976}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2098 ( .ina ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .inb ({new_AGEMA_signal_1022, new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2242}), .clk ( clk ), .rnd ({Fresh[849], Fresh[848], Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .outt ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, new_AGEMA_signal_1566, n2535}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2101 ( .ina ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .inb ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2356}), .clk ( clk ), .rnd ({Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852], Fresh[851], Fresh[850]}), .outt ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, new_AGEMA_signal_1569, n1973}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2105 ( .ina ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .inb ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .clk ( clk ), .rnd ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864], Fresh[863], Fresh[862], Fresh[861], Fresh[860]}), .outt ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, n2690}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2111 ( .ina ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2493}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[879], Fresh[878], Fresh[877], Fresh[876], Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .outt ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2113 ( .ina ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .inb ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, new_AGEMA_signal_1017, n2779}), .clk ( clk ), .rnd ({Fresh[889], Fresh[888], Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880]}), .outt ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, new_AGEMA_signal_1575, n2741}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2118 ( .ina ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .inb ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .clk ( clk ), .rnd ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890]}), .outt ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, new_AGEMA_signal_1578, n1992}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2120 ( .ina ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .outt ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, new_AGEMA_signal_1581, n1991}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2123 ( .ina ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .inb ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .clk ( clk ), .rnd ({Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912], Fresh[911], Fresh[910]}), .outt ({new_AGEMA_signal_1310, new_AGEMA_signal_1309, new_AGEMA_signal_1308, n1993}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2125 ( .ina ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}), .inb ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .clk ( clk ), .rnd ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924], Fresh[923], Fresh[922], Fresh[921], Fresh[920]}), .outt ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, new_AGEMA_signal_1584, n1995}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2132 ( .ina ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .inb ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .clk ( clk ), .rnd ({Fresh[939], Fresh[938], Fresh[937], Fresh[936], Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .outt ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, new_AGEMA_signal_1587, n2241}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2135 ( .ina ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .inb ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2679}), .clk ( clk ), .rnd ({Fresh[949], Fresh[948], Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942], Fresh[941], Fresh[940]}), .outt ({new_AGEMA_signal_1592, new_AGEMA_signal_1591, new_AGEMA_signal_1590, n2003}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2140 ( .ina ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .inb ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, n2809}), .clk ( clk ), .rnd ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950]}), .outt ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, new_AGEMA_signal_1593, n2008}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2141 ( .ina ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2679}), .inb ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .clk ( clk ), .rnd ({Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .outt ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, n2572}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2143 ( .ina ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, n2809}), .inb ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2356}), .clk ( clk ), .rnd ({Fresh[979], Fresh[978], Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972], Fresh[971], Fresh[970]}), .outt ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, new_AGEMA_signal_1599, n2004}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2147 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984], Fresh[983], Fresh[982], Fresh[981], Fresh[980]}), .outt ({new_AGEMA_signal_1604, new_AGEMA_signal_1603, new_AGEMA_signal_1602, n2009}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2151 ( .ina ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[999], Fresh[998], Fresh[997], Fresh[996], Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .outt ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2157 ( .ina ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .inb ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}), .clk ( clk ), .rnd ({Fresh[1009], Fresh[1008], Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000]}), .outt ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, new_AGEMA_signal_1323, n2026}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2158 ( .ina ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .inb ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2493}), .clk ( clk ), .rnd ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010]}), .outt ({new_AGEMA_signal_1610, new_AGEMA_signal_1609, new_AGEMA_signal_1608, n2022}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2159 ( .ina ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}), .inb ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .clk ( clk ), .rnd ({Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026], Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .outt ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2227}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2167 ( .ina ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[1039], Fresh[1038], Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032], Fresh[1031], Fresh[1030]}), .outt ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, new_AGEMA_signal_1143, n2027}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2171 ( .ina ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .inb ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .clk ( clk ), .rnd ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044], Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040]}), .outt ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, new_AGEMA_signal_1617, n2214}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2173 ( .ina ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .inb ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .rnd ({Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056], Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .outt ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, new_AGEMA_signal_1620, n2290}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2174 ( .ina ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .clk ( clk ), .rnd ({Fresh[1069], Fresh[1068], Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062], Fresh[1061], Fresh[1060]}), .outt ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2178 ( .ina ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .inb ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2400}), .clk ( clk ), .rnd ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074], Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070]}), .outt ({new_AGEMA_signal_1334, new_AGEMA_signal_1333, new_AGEMA_signal_1332, n2034}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2182 ( .ina ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .inb ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .clk ( clk ), .rnd ({Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086], Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .outt ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335, n2171}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2183 ( .ina ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, n2828}), .inb ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .clk ( clk ), .rnd ({Fresh[1099], Fresh[1098], Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092], Fresh[1091], Fresh[1090]}), .outt ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, new_AGEMA_signal_1626, n2039}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2188 ( .ina ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .inb ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .rnd ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104], Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100]}), .outt ({new_AGEMA_signal_1634, new_AGEMA_signal_1633, new_AGEMA_signal_1632, n2042}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2191 ( .ina ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .inb ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .clk ( clk ), .rnd ({Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116], Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .outt ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, new_AGEMA_signal_1635, n2754}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2192 ( .ina ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2313}), .inb ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .clk ( clk ), .rnd ({Fresh[1129], Fresh[1128], Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122], Fresh[1121], Fresh[1120]}), .outt ({new_AGEMA_signal_1640, new_AGEMA_signal_1639, new_AGEMA_signal_1638, n2044}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2198 ( .ina ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2313}), .inb ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .clk ( clk ), .rnd ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134], Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130]}), .outt ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, n2654}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2202 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, n2577}), .clk ( clk ), .rnd ({Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146], Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .outt ({new_AGEMA_signal_1646, new_AGEMA_signal_1645, new_AGEMA_signal_1644, n2055}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2205 ( .ina ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2395}), .inb ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .clk ( clk ), .rnd ({Fresh[1159], Fresh[1158], Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152], Fresh[1151], Fresh[1150]}), .outt ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, new_AGEMA_signal_1647, n2057}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2208 ( .ina ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2679}), .inb ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}), .clk ( clk ), .rnd ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164], Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160]}), .outt ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, new_AGEMA_signal_1650, n2407}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2212 ( .ina ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .inb ({new_AGEMA_signal_1148, new_AGEMA_signal_1147, new_AGEMA_signal_1146, n2061}), .clk ( clk ), .rnd ({Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176], Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .outt ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, new_AGEMA_signal_1653, n2062}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2216 ( .ina ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .inb ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}), .clk ( clk ), .rnd ({Fresh[1189], Fresh[1188], Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182], Fresh[1181], Fresh[1180]}), .outt ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, new_AGEMA_signal_1656, n2731}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2220 ( .a ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, n2690}), .b ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, new_AGEMA_signal_1659, n2068}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2224 ( .ina ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .inb ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .clk ( clk ), .rnd ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194], Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190]}), .outt ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, new_AGEMA_signal_1338, n2642}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2225 ( .ina ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .inb ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .clk ( clk ), .rnd ({Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206], Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .outt ({new_AGEMA_signal_1664, new_AGEMA_signal_1663, new_AGEMA_signal_1662, n2252}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2228 ( .ina ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, new_AGEMA_signal_1101, n2739}), .inb ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .clk ( clk ), .rnd ({Fresh[1219], Fresh[1218], Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212], Fresh[1211], Fresh[1210]}), .outt ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, new_AGEMA_signal_1341, n2075}) ) ;
    or_HPC1 #(.security_order(3), .pipeline(0)) U2233 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .clk ( clk ), .rnd ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224], Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220]}), .outt ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, new_AGEMA_signal_1344, n2081}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2234 ( .ina ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .inb ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}), .clk ( clk ), .rnd ({Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236], Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .outt ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, new_AGEMA_signal_1665, n2080}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2237 ( .ina ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2600}), .inb ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .clk ( clk ), .rnd ({Fresh[1249], Fresh[1248], Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242], Fresh[1241], Fresh[1240]}), .outt ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2238 ( .a ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .b ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, new_AGEMA_signal_1668, n2773}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2239 ( .ina ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .inb ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .clk ( clk ), .rnd ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254], Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250]}), .outt ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, new_AGEMA_signal_1671, n2083}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2244 ( .ina ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .inb ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, n2086}), .clk ( clk ), .rnd ({Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266], Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .outt ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, new_AGEMA_signal_1674, n2562}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2247 ( .ina ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}), .clk ( clk ), .rnd ({Fresh[1279], Fresh[1278], Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272], Fresh[1271], Fresh[1270]}), .outt ({new_AGEMA_signal_1352, new_AGEMA_signal_1351, new_AGEMA_signal_1350, n2087}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2251 ( .ina ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}), .inb ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, n2174}), .clk ( clk ), .rnd ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284], Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280]}), .outt ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, new_AGEMA_signal_1677, n2156}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2260 ( .ina ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .inb ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2401}), .clk ( clk ), .rnd ({Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296], Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .outt ({new_AGEMA_signal_1682, new_AGEMA_signal_1681, new_AGEMA_signal_1680, n2100}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2277 ( .ina ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, new_AGEMA_signal_1101, n2739}), .inb ({new_AGEMA_signal_1154, new_AGEMA_signal_1153, new_AGEMA_signal_1152, n2298}), .clk ( clk ), .rnd ({Fresh[1309], Fresh[1308], Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302], Fresh[1301], Fresh[1300]}), .outt ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, new_AGEMA_signal_1353, n2544}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2279 ( .ina ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2356}), .inb ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, new_AGEMA_signal_1356, n2118}), .clk ( clk ), .rnd ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314], Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310]}), .outt ({new_AGEMA_signal_1691, new_AGEMA_signal_1690, new_AGEMA_signal_1689, n2121}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2284 ( .ina ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .inb ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2570}), .clk ( clk ), .rnd ({Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326], Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .outt ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, new_AGEMA_signal_1695, n2122}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2286 ( .ina ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .inb ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .clk ( clk ), .rnd ({Fresh[1339], Fresh[1338], Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332], Fresh[1331], Fresh[1330]}), .outt ({new_AGEMA_signal_1700, new_AGEMA_signal_1699, new_AGEMA_signal_1698, n2811}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2294 ( .ina ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .inb ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .clk ( clk ), .rnd ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344], Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340]}), .outt ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, n2647}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2297 ( .ina ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .inb ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .clk ( clk ), .rnd ({Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356], Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .outt ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, new_AGEMA_signal_1362, n2132}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2304 ( .ina ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}), .inb ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .rnd ({Fresh[1369], Fresh[1368], Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362], Fresh[1361], Fresh[1360]}), .outt ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, new_AGEMA_signal_1713, n2220}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2305 ( .ina ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .inb ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .clk ( clk ), .rnd ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374], Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370]}), .outt ({new_AGEMA_signal_1718, new_AGEMA_signal_1717, new_AGEMA_signal_1716, n2138}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2312 ( .ina ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .inb ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .clk ( clk ), .rnd ({Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386], Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .outt ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, new_AGEMA_signal_1719, n2555}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2322 ( .ina ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .inb ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .clk ( clk ), .rnd ({Fresh[1399], Fresh[1398], Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392], Fresh[1391], Fresh[1390]}), .outt ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, n2429}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2328 ( .ina ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404], Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400]}), .outt ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, n2162}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2337 ( .ina ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .inb ({new_AGEMA_signal_1022, new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2242}), .clk ( clk ), .rnd ({Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416], Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .outt ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2545}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2340 ( .ina ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}), .inb ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .clk ( clk ), .rnd ({Fresh[1429], Fresh[1428], Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422], Fresh[1421], Fresh[1420]}), .outt ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, new_AGEMA_signal_1371, n2178}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2342 ( .ina ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, new_AGEMA_signal_1161, n2430}), .inb ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .rnd ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434], Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430]}), .outt ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, new_AGEMA_signal_1728, n2176}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2343 ( .ina ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, n2174}), .inb ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .rnd ({Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446], Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .outt ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, new_AGEMA_signal_1731, n2175}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2348 ( .ina ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}), .inb ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .clk ( clk ), .rnd ({Fresh[1459], Fresh[1458], Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452], Fresh[1451], Fresh[1450]}), .outt ({new_AGEMA_signal_1166, new_AGEMA_signal_1165, new_AGEMA_signal_1164, n2182}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2353 ( .ina ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .inb ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, new_AGEMA_signal_1161, n2430}), .clk ( clk ), .rnd ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464], Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460]}), .outt ({new_AGEMA_signal_1736, new_AGEMA_signal_1735, new_AGEMA_signal_1734, n2188}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2355 ( .ina ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .inb ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .clk ( clk ), .rnd ({Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476], Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .outt ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, new_AGEMA_signal_1737, n2189}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2357 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .clk ( clk ), .rnd ({Fresh[1489], Fresh[1488], Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482], Fresh[1481], Fresh[1480]}), .outt ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, new_AGEMA_signal_1740, n2446}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2362 ( .ina ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .inb ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}), .clk ( clk ), .rnd ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494], Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490]}), .outt ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, n2576}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2363 ( .ina ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .inb ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .clk ( clk ), .rnd ({Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506], Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .outt ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, new_AGEMA_signal_1380, n2748}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) U2368 ( .a ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, n2654}), .b ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, n2674}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2378 ( .ina ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .inb ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .clk ( clk ), .rnd ({Fresh[1519], Fresh[1518], Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512], Fresh[1511], Fresh[1510]}), .outt ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, n2213}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2380 ( .ina ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .inb ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524], Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520]}), .outt ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, new_AGEMA_signal_1386, n2215}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2384 ( .ina ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, n2712}), .inb ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .clk ( clk ), .rnd ({Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536], Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .outt ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, new_AGEMA_signal_1749, n2218}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2386 ( .ina ({new_AGEMA_signal_1154, new_AGEMA_signal_1153, new_AGEMA_signal_1152, n2298}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[1549], Fresh[1548], Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542], Fresh[1541], Fresh[1540]}), .outt ({new_AGEMA_signal_1754, new_AGEMA_signal_1753, new_AGEMA_signal_1752, n2219}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2405 ( .ina ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .inb ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .rnd ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554], Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550]}), .outt ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, new_AGEMA_signal_1767, n2240}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2407 ( .ina ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, new_AGEMA_signal_1320, n2709}), .inb ({new_AGEMA_signal_1022, new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2242}), .clk ( clk ), .rnd ({Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566], Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .outt ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, new_AGEMA_signal_1770, n2561}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2408 ( .ina ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .inb ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .clk ( clk ), .rnd ({Fresh[1579], Fresh[1578], Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572], Fresh[1571], Fresh[1570]}), .outt ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, new_AGEMA_signal_1773, n2243}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2411 ( .ina ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}), .inb ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .clk ( clk ), .rnd ({Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584], Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580]}), .outt ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, new_AGEMA_signal_1776, n2245}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2422 ( .ina ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .inb ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, new_AGEMA_signal_1161, n2430}), .clk ( clk ), .rnd ({Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596], Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590]}), .outt ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, new_AGEMA_signal_1779, n2540}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2423 ( .ina ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}), .inb ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2640}), .clk ( clk ), .rnd ({Fresh[1609], Fresh[1608], Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602], Fresh[1601], Fresh[1600]}), .outt ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, new_AGEMA_signal_1782, n2259}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2426 ( .ina ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}), .inb ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}), .clk ( clk ), .rnd ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614], Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610]}), .outt ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, new_AGEMA_signal_1389, n2262}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2431 ( .ina ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .inb ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, n2777}), .clk ( clk ), .rnd ({Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626], Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .outt ({new_AGEMA_signal_1394, new_AGEMA_signal_1393, new_AGEMA_signal_1392, n2266}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2432 ( .ina ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2772}), .inb ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .clk ( clk ), .rnd ({Fresh[1639], Fresh[1638], Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632], Fresh[1631], Fresh[1630]}), .outt ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, n2645}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2436 ( .ina ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .inb ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .clk ( clk ), .rnd ({Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644], Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640]}), .outt ({new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2268}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2443 ( .ina ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .inb ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .clk ( clk ), .rnd ({Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656], Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650]}), .outt ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, new_AGEMA_signal_1791, n2278}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2448 ( .ina ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .inb ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .rnd ({Fresh[1669], Fresh[1668], Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662], Fresh[1661], Fresh[1660]}), .outt ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, n2383}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2455 ( .ina ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .inb ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2570}), .clk ( clk ), .rnd ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674], Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670]}), .outt ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, new_AGEMA_signal_1800, n2774}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2458 ( .ina ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}), .inb ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .clk ( clk ), .rnd ({Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686], Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680]}), .outt ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, new_AGEMA_signal_1803, n2287}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2470 ( .ina ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .inb ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .rnd ({Fresh[1699], Fresh[1698], Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692], Fresh[1691], Fresh[1690]}), .outt ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, new_AGEMA_signal_1809, n2438}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2471 ( .ina ({new_AGEMA_signal_1154, new_AGEMA_signal_1153, new_AGEMA_signal_1152, n2298}), .inb ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .clk ( clk ), .rnd ({Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704], Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700]}), .outt ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, new_AGEMA_signal_1404, n2299}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2481 ( .ina ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .inb ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2313}), .clk ( clk ), .rnd ({Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716], Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710]}), .outt ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, new_AGEMA_signal_1812, n2371}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2484 ( .ina ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .inb ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .clk ( clk ), .rnd ({Fresh[1729], Fresh[1728], Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722], Fresh[1721], Fresh[1720]}), .outt ({new_AGEMA_signal_1172, new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2316}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2486 ( .ina ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, new_AGEMA_signal_1125, n2624}), .inb ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}), .clk ( clk ), .rnd ({Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734], Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730]}), .outt ({new_AGEMA_signal_1412, new_AGEMA_signal_1411, new_AGEMA_signal_1410, n2318}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2492 ( .ina ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746], Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740]}), .outt ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, new_AGEMA_signal_1821, n2325}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2494 ( .ina ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .inb ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .rnd ({Fresh[1759], Fresh[1758], Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752], Fresh[1751], Fresh[1750]}), .outt ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, new_AGEMA_signal_1824, n2328}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2495 ( .ina ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .inb ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .clk ( clk ), .rnd ({Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764], Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760]}), .outt ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, new_AGEMA_signal_1413, n2327}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2505 ( .ina ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}), .inb ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .clk ( clk ), .rnd ({Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776], Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770]}), .outt ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, new_AGEMA_signal_1827, n2343}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2510 ( .ina ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[1789], Fresh[1788], Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782], Fresh[1781], Fresh[1780]}), .outt ({new_AGEMA_signal_1835, new_AGEMA_signal_1834, new_AGEMA_signal_1833, n2344}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(0)) U2512 ( .ina ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2395}), .inb ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, new_AGEMA_signal_1155, n2346}), .clk ( clk ), .rnd ({Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794], Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790]}), .outt ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, new_AGEMA_signal_1416, n2348}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2513 ( .ina ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .inb ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .clk ( clk ), .rnd ({Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806], Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800]}), .outt ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, n2347}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2520 ( .ina ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .inb ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}), .clk ( clk ), .rnd ({Fresh[1819], Fresh[1818], Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812], Fresh[1811], Fresh[1810]}), .outt ({new_AGEMA_signal_1424, new_AGEMA_signal_1423, new_AGEMA_signal_1422, n2363}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2521 ( .ina ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, n2809}), .inb ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824], Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820]}), .outt ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, new_AGEMA_signal_1845, n2353}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2524 ( .ina ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .inb ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .rnd ({Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836], Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830]}), .outt ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, new_AGEMA_signal_1848, n2355}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2530 ( .ina ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, n2712}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[1849], Fresh[1848], Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842], Fresh[1841], Fresh[1840]}), .outt ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, new_AGEMA_signal_1851, n2364}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2543 ( .ina ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .inb ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2401}), .clk ( clk ), .rnd ({Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854], Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850]}), .outt ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, new_AGEMA_signal_1425, n2415}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2558 ( .ina ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2395}), .inb ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .clk ( clk ), .rnd ({Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866], Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860]}), .outt ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, new_AGEMA_signal_1428, n2700}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2563 ( .ina ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2400}), .clk ( clk ), .rnd ({Fresh[1879], Fresh[1878], Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872], Fresh[1871], Fresh[1870]}), .outt ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, n2594}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2564 ( .ina ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2401}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884], Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880]}), .outt ({new_AGEMA_signal_1436, new_AGEMA_signal_1435, new_AGEMA_signal_1434, n2402}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2585 ( .ina ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, n2712}), .inb ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}), .clk ( clk ), .rnd ({Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896], Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890]}), .outt ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, new_AGEMA_signal_1881, n2428}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2588 ( .ina ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, new_AGEMA_signal_1161, n2430}), .inb ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2570}), .clk ( clk ), .rnd ({Fresh[1909], Fresh[1908], Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902], Fresh[1901], Fresh[1900]}), .outt ({new_AGEMA_signal_1886, new_AGEMA_signal_1885, new_AGEMA_signal_1884, n2431}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2594 ( .ina ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .inb ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}), .clk ( clk ), .rnd ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914], Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910]}), .outt ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, n2483}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2599 ( .ina ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .inb ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .rnd ({Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926], Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .outt ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, new_AGEMA_signal_1890, n2443}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2606 ( .ina ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .inb ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .clk ( clk ), .rnd ({Fresh[1939], Fresh[1938], Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932], Fresh[1931], Fresh[1930]}), .outt ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, new_AGEMA_signal_1893, n2693}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2608 ( .ina ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2452}), .inb ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .rnd ({Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944], Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940]}), .outt ({new_AGEMA_signal_1442, new_AGEMA_signal_1441, new_AGEMA_signal_1440, n2453}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2616 ( .ina ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .inb ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, new_AGEMA_signal_1173, n2463}), .clk ( clk ), .rnd ({Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956], Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950]}), .outt ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443, n2464}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2620 ( .ina ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .inb ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .clk ( clk ), .rnd ({Fresh[1969], Fresh[1968], Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962], Fresh[1961], Fresh[1960]}), .outt ({new_AGEMA_signal_1448, new_AGEMA_signal_1447, new_AGEMA_signal_1446, n2468}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2624 ( .ina ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .inb ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974], Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970]}), .outt ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, new_AGEMA_signal_1449, n2473}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2625 ( .ina ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .inb ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .clk ( clk ), .rnd ({Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986], Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980]}), .outt ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, new_AGEMA_signal_1452, n2472}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2628 ( .ina ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}), .inb ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, new_AGEMA_signal_1176, n2474}), .clk ( clk ), .rnd ({Fresh[1999], Fresh[1998], Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992], Fresh[1991], Fresh[1990]}), .outt ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, new_AGEMA_signal_1455, n2475}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2632 ( .ina ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .inb ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, n2828}), .clk ( clk ), .rnd ({Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004], Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000]}), .outt ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, new_AGEMA_signal_1905, n2480}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2638 ( .ina ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, n2577}), .inb ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}), .clk ( clk ), .rnd ({Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016], Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010]}), .outt ({new_AGEMA_signal_1910, new_AGEMA_signal_1909, new_AGEMA_signal_1908, n2487}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2641 ( .ina ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}), .inb ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}), .clk ( clk ), .rnd ({Fresh[2029], Fresh[2028], Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022], Fresh[2021], Fresh[2020]}), .outt ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, new_AGEMA_signal_1458, n2488}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2665 ( .ina ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .inb ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .clk ( clk ), .rnd ({Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034], Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030]}), .outt ({new_AGEMA_signal_1928, new_AGEMA_signal_1927, new_AGEMA_signal_1926, n2520}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2667 ( .ina ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .inb ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, n2587}), .clk ( clk ), .rnd ({Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046], Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040]}), .outt ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, new_AGEMA_signal_1461, n2521}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2674 ( .ina ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}), .inb ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, new_AGEMA_signal_1005, n2595}), .clk ( clk ), .rnd ({Fresh[2059], Fresh[2058], Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052], Fresh[2051], Fresh[2050]}), .outt ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, new_AGEMA_signal_1929, n2531}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2689 ( .ina ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}), .inb ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .clk ( clk ), .rnd ({Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064], Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060]}), .outt ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, new_AGEMA_signal_1935, n2553}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2691 ( .ina ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .inb ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .clk ( clk ), .rnd ({Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076], Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070]}), .outt ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, new_AGEMA_signal_1938, n2554}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(0)) U2695 ( .ina ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}), .inb ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .clk ( clk ), .rnd ({Fresh[2089], Fresh[2088], Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082], Fresh[2081], Fresh[2080]}), .outt ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, new_AGEMA_signal_1464, n2560}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2698 ( .ina ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}), .inb ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}), .clk ( clk ), .rnd ({Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094], Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090]}), .outt ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, new_AGEMA_signal_1941, n2564}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2714 ( .ina ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .inb ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .clk ( clk ), .rnd ({Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106], Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100]}), .outt ({new_AGEMA_signal_1952, new_AGEMA_signal_1951, new_AGEMA_signal_1950, n2586}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2720 ( .ina ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, new_AGEMA_signal_1005, n2595}), .inb ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .clk ( clk ), .rnd ({Fresh[2119], Fresh[2118], Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112], Fresh[2111], Fresh[2110]}), .outt ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, new_AGEMA_signal_1467, n2597}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2721 ( .ina ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2640}), .inb ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .clk ( clk ), .rnd ({Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124], Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120]}), .outt ({new_AGEMA_signal_1958, new_AGEMA_signal_1957, new_AGEMA_signal_1956, n2596}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2723 ( .ina ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}), .inb ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .clk ( clk ), .rnd ({Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136], Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130]}), .outt ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, new_AGEMA_signal_1959, n2598}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2725 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[2149], Fresh[2148], Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142], Fresh[2141], Fresh[2140]}), .outt ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, n2599}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2732 ( .ina ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .inb ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .clk ( clk ), .rnd ({Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154], Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150]}), .outt ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, new_AGEMA_signal_1965, n2610}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2734 ( .ina ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .inb ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .clk ( clk ), .rnd ({Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166], Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160]}), .outt ({new_AGEMA_signal_1970, new_AGEMA_signal_1969, new_AGEMA_signal_1968, n2614}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2735 ( .ina ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .inb ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .clk ( clk ), .rnd ({Fresh[2179], Fresh[2178], Fresh[2177], Fresh[2176], Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172], Fresh[2171], Fresh[2170]}), .outt ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, new_AGEMA_signal_1971, n2613}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2737 ( .ina ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}), .inb ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}), .clk ( clk ), .rnd ({Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184], Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180]}), .outt ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, new_AGEMA_signal_1473, n2617}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2742 ( .ina ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, new_AGEMA_signal_1125, n2624}), .inb ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .clk ( clk ), .rnd ({Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196], Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190]}), .outt ({new_AGEMA_signal_1478, new_AGEMA_signal_1477, new_AGEMA_signal_1476, n2629}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2751 ( .ina ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .inb ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2640}), .clk ( clk ), .rnd ({Fresh[2209], Fresh[2208], Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202], Fresh[2201], Fresh[2200]}), .outt ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, new_AGEMA_signal_1977, n2784}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2757 ( .ina ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, n2785}), .inb ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, n2777}), .clk ( clk ), .rnd ({Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214], Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210]}), .outt ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, new_AGEMA_signal_1479, n2650}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2775 ( .ina ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .inb ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}), .clk ( clk ), .rnd ({Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226], Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220]}), .outt ({new_AGEMA_signal_1184, new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2683}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2789 ( .ina ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .inb ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .rnd ({Fresh[2239], Fresh[2238], Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232], Fresh[2231], Fresh[2230]}), .outt ({new_AGEMA_signal_2000, new_AGEMA_signal_1999, new_AGEMA_signal_1998, n2711}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2790 ( .ina ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, new_AGEMA_signal_1320, n2709}), .inb ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .clk ( clk ), .rnd ({Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244], Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240]}), .outt ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, new_AGEMA_signal_2001, n2710}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2792 ( .ina ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .inb ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, n2712}), .clk ( clk ), .rnd ({Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256], Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250]}), .outt ({new_AGEMA_signal_1484, new_AGEMA_signal_1483, new_AGEMA_signal_1482, n2714}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2797 ( .ina ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .inb ({new_AGEMA_signal_1151, new_AGEMA_signal_1150, new_AGEMA_signal_1149, n2721}), .clk ( clk ), .rnd ({Fresh[2269], Fresh[2268], Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262], Fresh[2261], Fresh[2260]}), .outt ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, new_AGEMA_signal_1485, n2722}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2799 ( .ina ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .inb ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}), .clk ( clk ), .rnd ({Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274], Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270]}), .outt ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, new_AGEMA_signal_2007, n2726}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2806 ( .ina ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}), .inb ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}), .clk ( clk ), .rnd ({Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286], Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280]}), .outt ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, new_AGEMA_signal_2010, n2738}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2822 ( .ina ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .inb ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .clk ( clk ), .rnd ({Fresh[2299], Fresh[2298], Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292], Fresh[2291], Fresh[2290]}), .outt ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, new_AGEMA_signal_2019, n2768}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2828 ( .ina ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .inb ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, n2777}), .clk ( clk ), .rnd ({Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304], Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300]}), .outt ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, new_AGEMA_signal_1488, n2782}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2829 ( .ina ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .inb ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, new_AGEMA_signal_1017, n2779}), .clk ( clk ), .rnd ({Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316], Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310]}), .outt ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, new_AGEMA_signal_1491, n2781}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2832 ( .ina ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .inb ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, n2785}), .clk ( clk ), .rnd ({Fresh[2329], Fresh[2328], Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322], Fresh[2321], Fresh[2320]}), .outt ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, new_AGEMA_signal_2025, n2787}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2834 ( .ina ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .inb ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .clk ( clk ), .rnd ({Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334], Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330]}), .outt ({new_AGEMA_signal_2030, new_AGEMA_signal_2029, new_AGEMA_signal_2028, n2794}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2835 ( .ina ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .inb ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .rnd ({Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346], Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340]}), .outt ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, new_AGEMA_signal_2031, n2793}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2844 ( .ina ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .inb ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, n2809}), .clk ( clk ), .rnd ({Fresh[2359], Fresh[2358], Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352], Fresh[2351], Fresh[2350]}), .outt ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, new_AGEMA_signal_2034, n2812}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2847 ( .ina ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .inb ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .clk ( clk ), .rnd ({Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364], Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360]}), .outt ({new_AGEMA_signal_1496, new_AGEMA_signal_1495, new_AGEMA_signal_1494, n2820}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2851 ( .ina ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}), .inb ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}), .clk ( clk ), .rnd ({Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376], Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370]}), .outt ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, new_AGEMA_signal_2040, n2825}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1960 ( .ina ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, new_AGEMA_signal_1497, n2575}), .inb ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, new_AGEMA_signal_1500, n1962}), .clk ( clk ), .rnd ({Fresh[2389], Fresh[2388], Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382], Fresh[2381], Fresh[2380]}), .outt ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, new_AGEMA_signal_2043, n1924}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1967 ( .ina ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, new_AGEMA_signal_1503, n1922}), .inb ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .clk ( clk ), .rnd ({Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394], Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390]}), .outt ({new_AGEMA_signal_2048, new_AGEMA_signal_2047, new_AGEMA_signal_2046, n1923}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1981 ( .ina ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, new_AGEMA_signal_1506, n1926}), .inb ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, new_AGEMA_signal_1509, n1925}), .clk ( clk ), .rnd ({Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406], Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400]}), .outt ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, new_AGEMA_signal_2049, n1927}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1993 ( .ina ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, n2734}), .inb ({new_AGEMA_signal_1520, new_AGEMA_signal_1519, new_AGEMA_signal_1518, n2763}), .clk ( clk ), .rnd ({Fresh[2419], Fresh[2418], Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412], Fresh[2411], Fresh[2410]}), .outt ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, new_AGEMA_signal_2052, n1929}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2007 ( .ina ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .clk ( clk ), .rnd ({Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424], Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420]}), .outt ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, new_AGEMA_signal_2055, n2665}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2011 ( .ina ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .inb ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, new_AGEMA_signal_1524, n1937}), .clk ( clk ), .rnd ({Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436], Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430]}), .outt ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, new_AGEMA_signal_2058, n1938}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2019 ( .ina ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, n2174}), .inb ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .clk ( clk ), .rnd ({Fresh[2449], Fresh[2448], Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442], Fresh[2441], Fresh[2440]}), .outt ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, new_AGEMA_signal_2061, n2235}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2023 ( .ina ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .inb ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, new_AGEMA_signal_1242, n1942}), .clk ( clk ), .rnd ({Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454], Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450]}), .outt ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, new_AGEMA_signal_1527, n1943}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2027 ( .ina ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, new_AGEMA_signal_1245, n2676}), .inb ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466], Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460]}), .outt ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, new_AGEMA_signal_1530, n1946}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2031 ( .ina ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2570}), .inb ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, new_AGEMA_signal_1533, n1944}), .clk ( clk ), .rnd ({Fresh[2479], Fresh[2478], Fresh[2477], Fresh[2476], Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472], Fresh[2471], Fresh[2470]}), .outt ({new_AGEMA_signal_2066, new_AGEMA_signal_2065, new_AGEMA_signal_2064, n1945}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2034 ( .ina ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .inb ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, n2734}), .clk ( clk ), .rnd ({Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484], Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480]}), .outt ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, new_AGEMA_signal_2067, n1956}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2040 ( .ina ({new_AGEMA_signal_1538, new_AGEMA_signal_1537, new_AGEMA_signal_1536, n1950}), .inb ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, new_AGEMA_signal_1254, n1949}), .clk ( clk ), .rnd ({Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496], Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490]}), .outt ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, new_AGEMA_signal_2070, n1951}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2048 ( .ina ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1539, n2662}), .inb ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .clk ( clk ), .rnd ({Fresh[2509], Fresh[2508], Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504], Fresh[2503], Fresh[2502], Fresh[2501], Fresh[2500]}), .outt ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, new_AGEMA_signal_2073, n1952}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2057 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, new_AGEMA_signal_1542, n2088}), .clk ( clk ), .rnd ({Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514], Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510]}), .outt ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, n2687}) ) ;
    or_HPC1 #(.security_order(3), .pipeline(0)) U2061 ( .ina ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, new_AGEMA_signal_1500, n1962}), .inb ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, n2587}), .clk ( clk ), .rnd ({Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526], Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520]}), .outt ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, new_AGEMA_signal_2079, n1966}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2064 ( .ina ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, n2736}), .inb ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .clk ( clk ), .rnd ({Fresh[2539], Fresh[2538], Fresh[2537], Fresh[2536], Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532], Fresh[2531], Fresh[2530]}), .outt ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, new_AGEMA_signal_1545, n1963}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2077 ( .ina ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, n2720}), .inb ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .clk ( clk ), .rnd ({Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544], Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540]}), .outt ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, new_AGEMA_signal_2556, n1968}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2082 ( .ina ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2505}), .inb ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .rnd ({Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556], Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550]}), .outt ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, new_AGEMA_signal_2091, n2684}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2088 ( .ina ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .inb ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2625}), .clk ( clk ), .rnd ({Fresh[2569], Fresh[2568], Fresh[2567], Fresh[2566], Fresh[2565], Fresh[2564], Fresh[2563], Fresh[2562], Fresh[2561], Fresh[2560]}), .outt ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, new_AGEMA_signal_2094, n1972}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2092 ( .ina ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .inb ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, n2190}), .clk ( clk ), .rnd ({Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576], Fresh[2575], Fresh[2574], Fresh[2573], Fresh[2572], Fresh[2571], Fresh[2570]}), .outt ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, new_AGEMA_signal_1563, n1971}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2099 ( .ina ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .inb ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, new_AGEMA_signal_1566, n2535}), .clk ( clk ), .rnd ({Fresh[2589], Fresh[2588], Fresh[2587], Fresh[2586], Fresh[2585], Fresh[2584], Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580]}), .outt ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, new_AGEMA_signal_2097, n1974}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2106 ( .ina ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .inb ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .clk ( clk ), .rnd ({Fresh[2599], Fresh[2598], Fresh[2597], Fresh[2596], Fresh[2595], Fresh[2594], Fresh[2593], Fresh[2592], Fresh[2591], Fresh[2590]}), .outt ({new_AGEMA_signal_2102, new_AGEMA_signal_2101, new_AGEMA_signal_2100, n1979}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2112 ( .ina ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .inb ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .rnd ({Fresh[2609], Fresh[2608], Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604], Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600]}), .outt ({new_AGEMA_signal_1574, new_AGEMA_signal_1573, new_AGEMA_signal_1572, n1985}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2121 ( .ina ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, new_AGEMA_signal_1578, n1992}), .inb ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, new_AGEMA_signal_1581, n1991}), .clk ( clk ), .rnd ({Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616], Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612], Fresh[2611], Fresh[2610]}), .outt ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, new_AGEMA_signal_2106, n1994}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2126 ( .ina ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2400}), .inb ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, new_AGEMA_signal_1584, n1995}), .clk ( clk ), .rnd ({Fresh[2629], Fresh[2628], Fresh[2627], Fresh[2626], Fresh[2625], Fresh[2624], Fresh[2623], Fresh[2622], Fresh[2621], Fresh[2620]}), .outt ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, new_AGEMA_signal_2109, n1996}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2136 ( .ina ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .inb ({new_AGEMA_signal_1592, new_AGEMA_signal_1591, new_AGEMA_signal_1590, n2003}), .clk ( clk ), .rnd ({Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636], Fresh[2635], Fresh[2634], Fresh[2633], Fresh[2632], Fresh[2631], Fresh[2630]}), .outt ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, new_AGEMA_signal_2112, n2137}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2142 ( .ina ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .inb ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, n2572}), .clk ( clk ), .rnd ({Fresh[2649], Fresh[2648], Fresh[2647], Fresh[2646], Fresh[2645], Fresh[2644], Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640]}), .outt ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, new_AGEMA_signal_2115, n2006}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2144 ( .ina ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .inb ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, new_AGEMA_signal_1599, n2004}), .clk ( clk ), .rnd ({Fresh[2659], Fresh[2658], Fresh[2657], Fresh[2656], Fresh[2655], Fresh[2654], Fresh[2653], Fresh[2652], Fresh[2651], Fresh[2650]}), .outt ({new_AGEMA_signal_2120, new_AGEMA_signal_2119, new_AGEMA_signal_2118, n2005}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2152 ( .ina ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, new_AGEMA_signal_1320, n2709}), .inb ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .clk ( clk ), .rnd ({Fresh[2669], Fresh[2668], Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664], Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660]}), .outt ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, new_AGEMA_signal_2121, n2013}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2160 ( .ina ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}), .inb ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2227}), .clk ( clk ), .rnd ({Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676], Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672], Fresh[2671], Fresh[2670]}), .outt ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, new_AGEMA_signal_1611, n2020}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2164 ( .ina ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .inb ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2401}), .clk ( clk ), .rnd ({Fresh[2689], Fresh[2688], Fresh[2687], Fresh[2686], Fresh[2685], Fresh[2684], Fresh[2683], Fresh[2682], Fresh[2681], Fresh[2680]}), .outt ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, new_AGEMA_signal_1614, n2023}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2168 ( .ina ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, new_AGEMA_signal_1143, n2027}), .inb ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .clk ( clk ), .rnd ({Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696], Fresh[2695], Fresh[2694], Fresh[2693], Fresh[2692], Fresh[2691], Fresh[2690]}), .outt ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, new_AGEMA_signal_1329, n2028}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2172 ( .ina ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, new_AGEMA_signal_1617, n2214}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[2709], Fresh[2708], Fresh[2707], Fresh[2706], Fresh[2705], Fresh[2704], Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700]}), .outt ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, new_AGEMA_signal_2127, n2033}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2175 ( .ina ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}), .inb ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}), .clk ( clk ), .rnd ({Fresh[2719], Fresh[2718], Fresh[2717], Fresh[2716], Fresh[2715], Fresh[2714], Fresh[2713], Fresh[2712], Fresh[2711], Fresh[2710]}), .outt ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, new_AGEMA_signal_2130, n2031}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2184 ( .ina ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .inb ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, new_AGEMA_signal_1626, n2039}), .clk ( clk ), .rnd ({Fresh[2729], Fresh[2728], Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724], Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720]}), .outt ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, new_AGEMA_signal_2133, n2040}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2187 ( .ina ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .inb ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .rnd ({Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736], Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732], Fresh[2731], Fresh[2730]}), .outt ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, new_AGEMA_signal_1629, n2050}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2193 ( .ina ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}), .inb ({new_AGEMA_signal_1640, new_AGEMA_signal_1639, new_AGEMA_signal_1638, n2044}), .clk ( clk ), .rnd ({Fresh[2749], Fresh[2748], Fresh[2747], Fresh[2746], Fresh[2745], Fresh[2744], Fresh[2743], Fresh[2742], Fresh[2741], Fresh[2740]}), .outt ({new_AGEMA_signal_2138, new_AGEMA_signal_2137, new_AGEMA_signal_2136, n2045}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2199 ( .ina ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, n2654}), .inb ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .clk ( clk ), .rnd ({Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756], Fresh[2755], Fresh[2754], Fresh[2753], Fresh[2752], Fresh[2751], Fresh[2750]}), .outt ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, new_AGEMA_signal_2139, n2051}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2203 ( .ina ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .inb ({new_AGEMA_signal_1646, new_AGEMA_signal_1645, new_AGEMA_signal_1644, n2055}), .clk ( clk ), .rnd ({Fresh[2769], Fresh[2768], Fresh[2767], Fresh[2766], Fresh[2765], Fresh[2764], Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760]}), .outt ({new_AGEMA_signal_2144, new_AGEMA_signal_2143, new_AGEMA_signal_2142, n2056}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2209 ( .ina ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, new_AGEMA_signal_1650, n2407}), .inb ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}), .clk ( clk ), .rnd ({Fresh[2779], Fresh[2778], Fresh[2777], Fresh[2776], Fresh[2775], Fresh[2774], Fresh[2773], Fresh[2772], Fresh[2771], Fresh[2770]}), .outt ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, new_AGEMA_signal_2145, n2060}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2215 ( .ina ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .inb ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, n2654}), .clk ( clk ), .rnd ({Fresh[2789], Fresh[2788], Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784], Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780]}), .outt ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, new_AGEMA_signal_2148, n2066}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2217 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, new_AGEMA_signal_1656, n2731}), .clk ( clk ), .rnd ({Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796], Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792], Fresh[2791], Fresh[2790]}), .outt ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, new_AGEMA_signal_2151, n2065}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2221 ( .ina ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, new_AGEMA_signal_1659, n2068}), .inb ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .rnd ({Fresh[2809], Fresh[2808], Fresh[2807], Fresh[2806], Fresh[2805], Fresh[2804], Fresh[2803], Fresh[2802], Fresh[2801], Fresh[2800]}), .outt ({new_AGEMA_signal_2156, new_AGEMA_signal_2155, new_AGEMA_signal_2154, n2069}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2226 ( .ina ({new_AGEMA_signal_1055, new_AGEMA_signal_1054, new_AGEMA_signal_1053, n2073}), .inb ({new_AGEMA_signal_1664, new_AGEMA_signal_1663, new_AGEMA_signal_1662, n2252}), .clk ( clk ), .rnd ({Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816], Fresh[2815], Fresh[2814], Fresh[2813], Fresh[2812], Fresh[2811], Fresh[2810]}), .outt ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, new_AGEMA_signal_2157, n2074}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2235 ( .ina ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, new_AGEMA_signal_1344, n2081}), .inb ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, new_AGEMA_signal_1665, n2080}), .clk ( clk ), .rnd ({Fresh[2829], Fresh[2828], Fresh[2827], Fresh[2826], Fresh[2825], Fresh[2824], Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820]}), .outt ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, new_AGEMA_signal_2160, n2082}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2240 ( .ina ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .inb ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, new_AGEMA_signal_1671, n2083}), .clk ( clk ), .rnd ({Fresh[2839], Fresh[2838], Fresh[2837], Fresh[2836], Fresh[2835], Fresh[2834], Fresh[2833], Fresh[2832], Fresh[2831], Fresh[2830]}), .outt ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, new_AGEMA_signal_2163, n2084}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2242 ( .ina ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .inb ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[2849], Fresh[2848], Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844], Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840]}), .outt ({new_AGEMA_signal_2168, new_AGEMA_signal_2167, new_AGEMA_signal_2166, n2085}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2245 ( .ina ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .inb ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, new_AGEMA_signal_1674, n2562}), .clk ( clk ), .rnd ({Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856], Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852], Fresh[2851], Fresh[2850]}), .outt ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, new_AGEMA_signal_2169, n2131}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2248 ( .ina ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, new_AGEMA_signal_1542, n2088}), .inb ({new_AGEMA_signal_1352, new_AGEMA_signal_1351, new_AGEMA_signal_1350, n2087}), .clk ( clk ), .rnd ({Fresh[2869], Fresh[2868], Fresh[2867], Fresh[2866], Fresh[2865], Fresh[2864], Fresh[2863], Fresh[2862], Fresh[2861], Fresh[2860]}), .outt ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, new_AGEMA_signal_2172, n2089}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2252 ( .ina ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .inb ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, new_AGEMA_signal_1677, n2156}), .clk ( clk ), .rnd ({Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876], Fresh[2875], Fresh[2874], Fresh[2873], Fresh[2872], Fresh[2871], Fresh[2870]}), .outt ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, new_AGEMA_signal_2175, n2330}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2254 ( .ina ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}), .inb ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, new_AGEMA_signal_1512, n2151}), .clk ( clk ), .rnd ({Fresh[2889], Fresh[2888], Fresh[2887], Fresh[2886], Fresh[2885], Fresh[2884], Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880]}), .outt ({new_AGEMA_signal_2180, new_AGEMA_signal_2179, new_AGEMA_signal_2178, n2092}) ) ;
    or_HPC1 #(.security_order(3), .pipeline(0)) U2256 ( .ina ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}), .inb ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, new_AGEMA_signal_1557, n2359}), .clk ( clk ), .rnd ({Fresh[2899], Fresh[2898], Fresh[2897], Fresh[2896], Fresh[2895], Fresh[2894], Fresh[2893], Fresh[2892], Fresh[2891], Fresh[2890]}), .outt ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, new_AGEMA_signal_2181, n2094}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2261 ( .ina ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, n2101}), .inb ({new_AGEMA_signal_1682, new_AGEMA_signal_1681, new_AGEMA_signal_1680, n2100}), .clk ( clk ), .rnd ({Fresh[2909], Fresh[2908], Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904], Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900]}), .outt ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, new_AGEMA_signal_2184, n2160}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2265 ( .ina ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916], Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912], Fresh[2911], Fresh[2910]}), .outt ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, n2504}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2271 ( .ina ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .inb ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .rnd ({Fresh[2929], Fresh[2928], Fresh[2927], Fresh[2926], Fresh[2925], Fresh[2924], Fresh[2923], Fresh[2922], Fresh[2921], Fresh[2920]}), .outt ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, new_AGEMA_signal_2628, n2114}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2273 ( .ina ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, n2677}), .inb ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .clk ( clk ), .rnd ({Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936], Fresh[2935], Fresh[2934], Fresh[2933], Fresh[2932], Fresh[2931], Fresh[2930]}), .outt ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, new_AGEMA_signal_1686, n2115}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2280 ( .ina ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .inb ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, new_AGEMA_signal_1656, n2731}), .clk ( clk ), .rnd ({Fresh[2949], Fresh[2948], Fresh[2947], Fresh[2946], Fresh[2945], Fresh[2944], Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940]}), .outt ({new_AGEMA_signal_2192, new_AGEMA_signal_2191, new_AGEMA_signal_2190, n2291}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2281 ( .ina ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .clk ( clk ), .rnd ({Fresh[2959], Fresh[2958], Fresh[2957], Fresh[2956], Fresh[2955], Fresh[2954], Fresh[2953], Fresh[2952], Fresh[2951], Fresh[2950]}), .outt ({new_AGEMA_signal_1694, new_AGEMA_signal_1693, new_AGEMA_signal_1692, n2119}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2291 ( .ina ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .inb ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .clk ( clk ), .rnd ({Fresh[2969], Fresh[2968], Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964], Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960]}), .outt ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, new_AGEMA_signal_1701, n2130}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2292 ( .ina ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .inb ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2631}), .clk ( clk ), .rnd ({Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976], Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972], Fresh[2971], Fresh[2970]}), .outt ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, new_AGEMA_signal_1704, n2129}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2295 ( .ina ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, n2647}), .inb ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .rnd ({Fresh[2989], Fresh[2988], Fresh[2987], Fresh[2986], Fresh[2985], Fresh[2984], Fresh[2983], Fresh[2982], Fresh[2981], Fresh[2980]}), .outt ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, new_AGEMA_signal_1707, n2150}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2298 ( .ina ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}), .inb ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, new_AGEMA_signal_1362, n2132}), .clk ( clk ), .rnd ({Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996], Fresh[2995], Fresh[2994], Fresh[2993], Fresh[2992], Fresh[2991], Fresh[2990]}), .outt ({new_AGEMA_signal_1712, new_AGEMA_signal_1711, new_AGEMA_signal_1710, n2133}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2302 ( .ina ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .inb ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .clk ( clk ), .rnd ({Fresh[3009], Fresh[3008], Fresh[3007], Fresh[3006], Fresh[3005], Fresh[3004], Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000]}), .outt ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, new_AGEMA_signal_2199, n2136}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2306 ( .ina ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, n2572}), .inb ({new_AGEMA_signal_1718, new_AGEMA_signal_1717, new_AGEMA_signal_1716, n2138}), .clk ( clk ), .rnd ({Fresh[3019], Fresh[3018], Fresh[3017], Fresh[3016], Fresh[3015], Fresh[3014], Fresh[3013], Fresh[3012], Fresh[3011], Fresh[3010]}), .outt ({new_AGEMA_signal_2204, new_AGEMA_signal_2203, new_AGEMA_signal_2202, n2139}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2313 ( .ina ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}), .inb ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, new_AGEMA_signal_1719, n2555}), .clk ( clk ), .rnd ({Fresh[3029], Fresh[3028], Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024], Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020]}), .outt ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, new_AGEMA_signal_2205, n2144}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2318 ( .ina ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, new_AGEMA_signal_1512, n2151}), .inb ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .clk ( clk ), .rnd ({Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036], Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032], Fresh[3031], Fresh[3030]}), .outt ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, new_AGEMA_signal_2208, n2152}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2321 ( .ina ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .inb ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, new_AGEMA_signal_1677, n2156}), .clk ( clk ), .rnd ({Fresh[3049], Fresh[3048], Fresh[3047], Fresh[3046], Fresh[3045], Fresh[3044], Fresh[3043], Fresh[3042], Fresh[3041], Fresh[3040]}), .outt ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, new_AGEMA_signal_2211, n2170}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2323 ( .ina ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, n2429}), .inb ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .clk ( clk ), .rnd ({Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056], Fresh[3055], Fresh[3054], Fresh[3053], Fresh[3052], Fresh[3051], Fresh[3050]}), .outt ({new_AGEMA_signal_2216, new_AGEMA_signal_2215, new_AGEMA_signal_2214, n2157}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2329 ( .ina ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}), .inb ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, n2162}), .clk ( clk ), .rnd ({Fresh[3069], Fresh[3068], Fresh[3067], Fresh[3066], Fresh[3065], Fresh[3064], Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060]}), .outt ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, new_AGEMA_signal_1725, n2163}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2335 ( .ina ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335, n2171}), .inb ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}), .clk ( clk ), .rnd ({Fresh[3079], Fresh[3078], Fresh[3077], Fresh[3076], Fresh[3075], Fresh[3074], Fresh[3073], Fresh[3072], Fresh[3071], Fresh[3070]}), .outt ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, new_AGEMA_signal_2220, n2172}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2338 ( .ina ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2545}), .clk ( clk ), .rnd ({Fresh[3089], Fresh[3088], Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084], Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080]}), .outt ({new_AGEMA_signal_1370, new_AGEMA_signal_1369, new_AGEMA_signal_1368, n2186}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2339 ( .ina ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .inb ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, new_AGEMA_signal_1620, n2290}), .clk ( clk ), .rnd ({Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096], Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092], Fresh[3091], Fresh[3090]}), .outt ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, new_AGEMA_signal_2223, n2181}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2344 ( .ina ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, new_AGEMA_signal_1728, n2176}), .inb ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, new_AGEMA_signal_1731, n2175}), .clk ( clk ), .rnd ({Fresh[3109], Fresh[3108], Fresh[3107], Fresh[3106], Fresh[3105], Fresh[3104], Fresh[3103], Fresh[3102], Fresh[3101], Fresh[3100]}), .outt ({new_AGEMA_signal_2228, new_AGEMA_signal_2227, new_AGEMA_signal_2226, n2177}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2349 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_1166, new_AGEMA_signal_1165, new_AGEMA_signal_1164, n2182}), .clk ( clk ), .rnd ({Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116], Fresh[3115], Fresh[3114], Fresh[3113], Fresh[3112], Fresh[3111], Fresh[3110]}), .outt ({new_AGEMA_signal_1376, new_AGEMA_signal_1375, new_AGEMA_signal_1374, n2183}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2354 ( .ina ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .inb ({new_AGEMA_signal_1736, new_AGEMA_signal_1735, new_AGEMA_signal_1734, n2188}), .clk ( clk ), .rnd ({Fresh[3129], Fresh[3128], Fresh[3127], Fresh[3126], Fresh[3125], Fresh[3124], Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120]}), .outt ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, new_AGEMA_signal_2229, n2195}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2356 ( .ina ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, n2190}), .inb ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, new_AGEMA_signal_1737, n2189}), .clk ( clk ), .rnd ({Fresh[3139], Fresh[3138], Fresh[3137], Fresh[3136], Fresh[3135], Fresh[3134], Fresh[3133], Fresh[3132], Fresh[3131], Fresh[3130]}), .outt ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, new_AGEMA_signal_2232, n2193}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2358 ( .ina ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .inb ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, new_AGEMA_signal_1740, n2446}), .clk ( clk ), .rnd ({Fresh[3149], Fresh[3148], Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144], Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140]}), .outt ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, new_AGEMA_signal_2235, n2191}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2364 ( .ina ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, n2576}), .inb ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, new_AGEMA_signal_1380, n2748}), .clk ( clk ), .rnd ({Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156], Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152], Fresh[3151], Fresh[3150]}), .outt ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, new_AGEMA_signal_1743, n2196}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2367 ( .ina ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2505}), .clk ( clk ), .rnd ({Fresh[3169], Fresh[3168], Fresh[3167], Fresh[3166], Fresh[3165], Fresh[3164], Fresh[3163], Fresh[3162], Fresh[3161], Fresh[3160]}), .outt ({new_AGEMA_signal_2240, new_AGEMA_signal_2239, new_AGEMA_signal_2238, n2201}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2369 ( .ina ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, n2674}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176], Fresh[3175], Fresh[3174], Fresh[3173], Fresh[3172], Fresh[3171], Fresh[3170]}), .outt ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, new_AGEMA_signal_2661, n2200}) ) ;
    mux2_HPC1 #(.security_order(3), .pipeline(0)) U2371 ( .ins ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .inb ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, n2734}), .ina ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .clk ( clk ), .rnd ({Fresh[3189], Fresh[3188], Fresh[3187], Fresh[3186], Fresh[3185], Fresh[3184], Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180]}), .outt ({new_AGEMA_signal_2666, new_AGEMA_signal_2665, new_AGEMA_signal_2664, n2202}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2379 ( .ina ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, new_AGEMA_signal_1617, n2214}), .inb ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, n2213}), .clk ( clk ), .rnd ({Fresh[3199], Fresh[3198], Fresh[3197], Fresh[3196], Fresh[3195], Fresh[3194], Fresh[3193], Fresh[3192], Fresh[3191], Fresh[3190]}), .outt ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, new_AGEMA_signal_2244, n2217}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2381 ( .ina ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2640}), .inb ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, new_AGEMA_signal_1386, n2215}), .clk ( clk ), .rnd ({Fresh[3209], Fresh[3208], Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204], Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200]}), .outt ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, new_AGEMA_signal_1746, n2216}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2385 ( .ina ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, new_AGEMA_signal_1749, n2218}), .inb ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .clk ( clk ), .rnd ({Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216], Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212], Fresh[3211], Fresh[3210]}), .outt ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, new_AGEMA_signal_2247, n2222}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2387 ( .ina ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, new_AGEMA_signal_1713, n2220}), .inb ({new_AGEMA_signal_1754, new_AGEMA_signal_1753, new_AGEMA_signal_1752, n2219}), .clk ( clk ), .rnd ({Fresh[3229], Fresh[3228], Fresh[3227], Fresh[3226], Fresh[3225], Fresh[3224], Fresh[3223], Fresh[3222], Fresh[3221], Fresh[3220]}), .outt ({new_AGEMA_signal_2252, new_AGEMA_signal_2251, new_AGEMA_signal_2250, n2221}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2391 ( .ina ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .inb ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .rnd ({Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236], Fresh[3235], Fresh[3234], Fresh[3233], Fresh[3232], Fresh[3231], Fresh[3230]}), .outt ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, new_AGEMA_signal_1755, n2226}) ) ;
    mux2_HPC1 #(.security_order(3), .pipeline(0)) U2393 ( .ins ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .inb ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .ina ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2227}), .clk ( clk ), .rnd ({Fresh[3249], Fresh[3248], Fresh[3247], Fresh[3246], Fresh[3245], Fresh[3244], Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240]}), .outt ({new_AGEMA_signal_1760, new_AGEMA_signal_1759, new_AGEMA_signal_1758, n2228}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2397 ( .ina ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}), .inb ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .rnd ({Fresh[3259], Fresh[3258], Fresh[3257], Fresh[3256], Fresh[3255], Fresh[3254], Fresh[3253], Fresh[3252], Fresh[3251], Fresh[3250]}), .outt ({new_AGEMA_signal_1763, new_AGEMA_signal_1762, new_AGEMA_signal_1761, n2237}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2398 ( .ina ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .inb ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .rnd ({Fresh[3269], Fresh[3268], Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264], Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260]}), .outt ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, new_AGEMA_signal_2676, n2233}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2403 ( .ina ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, n2777}), .inb ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2631}), .clk ( clk ), .rnd ({Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276], Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272], Fresh[3271], Fresh[3270]}), .outt ({new_AGEMA_signal_1766, new_AGEMA_signal_1765, new_AGEMA_signal_1764, n2238}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2406 ( .ina ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, new_AGEMA_signal_1587, n2241}), .inb ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, new_AGEMA_signal_1767, n2240}), .clk ( clk ), .rnd ({Fresh[3289], Fresh[3288], Fresh[3287], Fresh[3286], Fresh[3285], Fresh[3284], Fresh[3283], Fresh[3282], Fresh[3281], Fresh[3280]}), .outt ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, new_AGEMA_signal_2256, n2248}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2409 ( .ina ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, new_AGEMA_signal_1770, n2561}), .inb ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, new_AGEMA_signal_1773, n2243}), .clk ( clk ), .rnd ({Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296], Fresh[3295], Fresh[3294], Fresh[3293], Fresh[3292], Fresh[3291], Fresh[3290]}), .outt ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, new_AGEMA_signal_2259, n2244}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2414 ( .ina ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}), .inb ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .clk ( clk ), .rnd ({Fresh[3309], Fresh[3308], Fresh[3307], Fresh[3306], Fresh[3305], Fresh[3304], Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300]}), .outt ({new_AGEMA_signal_2264, new_AGEMA_signal_2263, new_AGEMA_signal_2262, n2249}) ) ;
    mux2_HPC1 #(.security_order(3), .pipeline(0)) U2417 ( .ins ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .inb ({new_AGEMA_signal_1664, new_AGEMA_signal_1663, new_AGEMA_signal_1662, n2252}), .ina ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .rnd ({Fresh[3319], Fresh[3318], Fresh[3317], Fresh[3316], Fresh[3315], Fresh[3314], Fresh[3313], Fresh[3312], Fresh[3311], Fresh[3310]}), .outt ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, new_AGEMA_signal_2265, n2253}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2424 ( .ina ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .inb ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, new_AGEMA_signal_1782, n2259}), .clk ( clk ), .rnd ({Fresh[3329], Fresh[3328], Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324], Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320]}), .outt ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, new_AGEMA_signal_2268, n2260}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2429 ( .ina ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .inb ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .clk ( clk ), .rnd ({Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336], Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332], Fresh[3331], Fresh[3330]}), .outt ({new_AGEMA_signal_2690, new_AGEMA_signal_2689, new_AGEMA_signal_2688, n2273}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2430 ( .ina ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}), .inb ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, n2720}), .clk ( clk ), .rnd ({Fresh[3349], Fresh[3348], Fresh[3347], Fresh[3346], Fresh[3345], Fresh[3344], Fresh[3343], Fresh[3342], Fresh[3341], Fresh[3340]}), .outt ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, new_AGEMA_signal_2691, n2752}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2433 ( .ina ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, n2645}), .inb ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .rnd ({Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356], Fresh[3355], Fresh[3354], Fresh[3353], Fresh[3352], Fresh[3351], Fresh[3350]}), .outt ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, new_AGEMA_signal_1785, n2265}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2437 ( .ina ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}), .inb ({new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2268}), .clk ( clk ), .rnd ({Fresh[3369], Fresh[3368], Fresh[3367], Fresh[3366], Fresh[3365], Fresh[3364], Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360]}), .outt ({new_AGEMA_signal_1790, new_AGEMA_signal_1789, new_AGEMA_signal_1788, n2269}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2444 ( .ina ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .inb ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .rnd ({Fresh[3379], Fresh[3378], Fresh[3377], Fresh[3376], Fresh[3375], Fresh[3374], Fresh[3373], Fresh[3372], Fresh[3371], Fresh[3370]}), .outt ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, new_AGEMA_signal_1794, n2277}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2449 ( .ina ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .inb ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, n2383}), .clk ( clk ), .rnd ({Fresh[3389], Fresh[3388], Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384], Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380]}), .outt ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, new_AGEMA_signal_1797, n2282}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2452 ( .ina ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, n2736}), .inb ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .clk ( clk ), .rnd ({Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396], Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392], Fresh[3391], Fresh[3390]}), .outt ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, new_AGEMA_signal_2283, n2284}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2456 ( .ina ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, new_AGEMA_signal_1800, n2774}), .inb ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .clk ( clk ), .rnd ({Fresh[3409], Fresh[3408], Fresh[3407], Fresh[3406], Fresh[3405], Fresh[3404], Fresh[3403], Fresh[3402], Fresh[3401], Fresh[3400]}), .outt ({new_AGEMA_signal_2288, new_AGEMA_signal_2287, new_AGEMA_signal_2286, n2459}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2459 ( .ina ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .inb ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, new_AGEMA_signal_1803, n2287}), .clk ( clk ), .rnd ({Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416], Fresh[3415], Fresh[3414], Fresh[3413], Fresh[3412], Fresh[3411], Fresh[3410]}), .outt ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, new_AGEMA_signal_2289, n2288}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2462 ( .ina ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}), .clk ( clk ), .rnd ({Fresh[3429], Fresh[3428], Fresh[3427], Fresh[3426], Fresh[3425], Fresh[3424], Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420]}), .outt ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, new_AGEMA_signal_2292, n2458}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2464 ( .ina ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}), .inb ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, new_AGEMA_signal_1620, n2290}), .clk ( clk ), .rnd ({Fresh[3439], Fresh[3438], Fresh[3437], Fresh[3436], Fresh[3435], Fresh[3434], Fresh[3433], Fresh[3432], Fresh[3431], Fresh[3430]}), .outt ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, new_AGEMA_signal_2295, n2293}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2467 ( .ina ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}), .inb ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, new_AGEMA_signal_1338, n2642}), .clk ( clk ), .rnd ({Fresh[3449], Fresh[3448], Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444], Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440]}), .outt ({new_AGEMA_signal_1808, new_AGEMA_signal_1807, new_AGEMA_signal_1806, n2294}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2472 ( .ina ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, new_AGEMA_signal_1809, n2438}), .inb ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, new_AGEMA_signal_1404, n2299}), .clk ( clk ), .rnd ({Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456], Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452], Fresh[3451], Fresh[3450]}), .outt ({new_AGEMA_signal_2300, new_AGEMA_signal_2299, new_AGEMA_signal_2298, n2300}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2480 ( .ina ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, n2734}), .inb ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .clk ( clk ), .rnd ({Fresh[3469], Fresh[3468], Fresh[3467], Fresh[3466], Fresh[3465], Fresh[3464], Fresh[3463], Fresh[3462], Fresh[3461], Fresh[3460]}), .outt ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, new_AGEMA_signal_2301, n2323}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(0)) U2482 ( .ina ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, n2571}), .inb ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, new_AGEMA_signal_1812, n2371}), .clk ( clk ), .rnd ({Fresh[3479], Fresh[3478], Fresh[3477], Fresh[3476], Fresh[3475], Fresh[3474], Fresh[3473], Fresh[3472], Fresh[3471], Fresh[3470]}), .outt ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, new_AGEMA_signal_2304, n2314}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2485 ( .ina ({new_AGEMA_signal_1172, new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2316}), .inb ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}), .clk ( clk ), .rnd ({Fresh[3489], Fresh[3488], Fresh[3487], Fresh[3486], Fresh[3485], Fresh[3484], Fresh[3483], Fresh[3482], Fresh[3481], Fresh[3480]}), .outt ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, n2319}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2491 ( .ina ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, new_AGEMA_signal_1338, n2642}), .inb ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .clk ( clk ), .rnd ({Fresh[3499], Fresh[3498], Fresh[3497], Fresh[3496], Fresh[3495], Fresh[3494], Fresh[3493], Fresh[3492], Fresh[3491], Fresh[3490]}), .outt ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, new_AGEMA_signal_1818, n2326}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2496 ( .ina ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, new_AGEMA_signal_1824, n2328}), .inb ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, new_AGEMA_signal_1413, n2327}), .clk ( clk ), .rnd ({Fresh[3509], Fresh[3508], Fresh[3507], Fresh[3506], Fresh[3505], Fresh[3504], Fresh[3503], Fresh[3502], Fresh[3501], Fresh[3500]}), .outt ({new_AGEMA_signal_2312, new_AGEMA_signal_2311, new_AGEMA_signal_2310, n2329}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2501 ( .ina ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .inb ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, n2674}), .clk ( clk ), .rnd ({Fresh[3519], Fresh[3518], Fresh[3517], Fresh[3516], Fresh[3515], Fresh[3514], Fresh[3513], Fresh[3512], Fresh[3511], Fresh[3510]}), .outt ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, new_AGEMA_signal_2727, n2335}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2506 ( .ina ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, new_AGEMA_signal_1320, n2709}), .inb ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}), .clk ( clk ), .rnd ({Fresh[3529], Fresh[3528], Fresh[3527], Fresh[3526], Fresh[3525], Fresh[3524], Fresh[3523], Fresh[3522], Fresh[3521], Fresh[3520]}), .outt ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, new_AGEMA_signal_2313, n2341}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2507 ( .ina ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .inb ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, n2736}), .clk ( clk ), .rnd ({Fresh[3539], Fresh[3538], Fresh[3537], Fresh[3536], Fresh[3535], Fresh[3534], Fresh[3533], Fresh[3532], Fresh[3531], Fresh[3530]}), .outt ({new_AGEMA_signal_1832, new_AGEMA_signal_1831, new_AGEMA_signal_1830, n2340}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2514 ( .ina ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, new_AGEMA_signal_1416, n2348}), .inb ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, n2347}), .clk ( clk ), .rnd ({Fresh[3549], Fresh[3548], Fresh[3547], Fresh[3546], Fresh[3545], Fresh[3544], Fresh[3543], Fresh[3542], Fresh[3541], Fresh[3540]}), .outt ({new_AGEMA_signal_1838, new_AGEMA_signal_1837, new_AGEMA_signal_1836, n2349}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2517 ( .ina ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, new_AGEMA_signal_1125, n2624}), .inb ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, n2690}), .clk ( clk ), .rnd ({Fresh[3559], Fresh[3558], Fresh[3557], Fresh[3556], Fresh[3555], Fresh[3554], Fresh[3553], Fresh[3552], Fresh[3551], Fresh[3550]}), .outt ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, new_AGEMA_signal_1839, n2375}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2518 ( .ina ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}), .inb ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, n2736}), .clk ( clk ), .rnd ({Fresh[3569], Fresh[3568], Fresh[3567], Fresh[3566], Fresh[3565], Fresh[3564], Fresh[3563], Fresh[3562], Fresh[3561], Fresh[3560]}), .outt ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, new_AGEMA_signal_1842, n2352}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2522 ( .ina ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, new_AGEMA_signal_1845, n2353}), .inb ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .clk ( clk ), .rnd ({Fresh[3579], Fresh[3578], Fresh[3577], Fresh[3576], Fresh[3575], Fresh[3574], Fresh[3573], Fresh[3572], Fresh[3571], Fresh[3570]}), .outt ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319, n2354}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2525 ( .ina ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2356}), .inb ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, new_AGEMA_signal_1848, n2355}), .clk ( clk ), .rnd ({Fresh[3589], Fresh[3588], Fresh[3587], Fresh[3586], Fresh[3585], Fresh[3584], Fresh[3583], Fresh[3582], Fresh[3581], Fresh[3580]}), .outt ({new_AGEMA_signal_2324, new_AGEMA_signal_2323, new_AGEMA_signal_2322, n2357}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2527 ( .ina ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, new_AGEMA_signal_1557, n2359}), .inb ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .clk ( clk ), .rnd ({Fresh[3599], Fresh[3598], Fresh[3597], Fresh[3596], Fresh[3595], Fresh[3594], Fresh[3593], Fresh[3592], Fresh[3591], Fresh[3590]}), .outt ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, new_AGEMA_signal_2325, n2360}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2534 ( .ina ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, n2674}), .clk ( clk ), .rnd ({Fresh[3609], Fresh[3608], Fresh[3607], Fresh[3606], Fresh[3605], Fresh[3604], Fresh[3603], Fresh[3602], Fresh[3601], Fresh[3600]}), .outt ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, new_AGEMA_signal_2736, n2369}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2536 ( .ina ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, new_AGEMA_signal_1812, n2371}), .inb ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .rnd ({Fresh[3619], Fresh[3618], Fresh[3617], Fresh[3616], Fresh[3615], Fresh[3614], Fresh[3613], Fresh[3612], Fresh[3611], Fresh[3610]}), .outt ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, new_AGEMA_signal_2328, n2372}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2539 ( .ina ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, n2576}), .inb ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}), .clk ( clk ), .rnd ({Fresh[3629], Fresh[3628], Fresh[3627], Fresh[3626], Fresh[3625], Fresh[3624], Fresh[3623], Fresh[3622], Fresh[3621], Fresh[3620]}), .outt ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, new_AGEMA_signal_2331, n2377}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2544 ( .ina ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .inb ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, new_AGEMA_signal_1425, n2415}), .clk ( clk ), .rnd ({Fresh[3639], Fresh[3638], Fresh[3637], Fresh[3636], Fresh[3635], Fresh[3634], Fresh[3633], Fresh[3632], Fresh[3631], Fresh[3630]}), .outt ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, new_AGEMA_signal_1854, n2467}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2545 ( .ina ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .inb ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, n2383}), .clk ( clk ), .rnd ({Fresh[3649], Fresh[3648], Fresh[3647], Fresh[3646], Fresh[3645], Fresh[3644], Fresh[3643], Fresh[3642], Fresh[3641], Fresh[3640]}), .outt ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, new_AGEMA_signal_1857, n2385}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2546 ( .ina ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[3659], Fresh[3658], Fresh[3657], Fresh[3656], Fresh[3655], Fresh[3654], Fresh[3653], Fresh[3652], Fresh[3651], Fresh[3650]}), .outt ({new_AGEMA_signal_1862, new_AGEMA_signal_1861, new_AGEMA_signal_1860, n2384}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2548 ( .ina ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .inb ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, n2429}), .clk ( clk ), .rnd ({Fresh[3669], Fresh[3668], Fresh[3667], Fresh[3666], Fresh[3665], Fresh[3664], Fresh[3663], Fresh[3662], Fresh[3661], Fresh[3660]}), .outt ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, new_AGEMA_signal_2337, n2386}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2552 ( .ina ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .inb ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, n2647}), .clk ( clk ), .rnd ({Fresh[3679], Fresh[3678], Fresh[3677], Fresh[3676], Fresh[3675], Fresh[3674], Fresh[3673], Fresh[3672], Fresh[3671], Fresh[3670]}), .outt ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, new_AGEMA_signal_1863, n2394}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2553 ( .ina ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .inb ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .clk ( clk ), .rnd ({Fresh[3689], Fresh[3688], Fresh[3687], Fresh[3686], Fresh[3685], Fresh[3684], Fresh[3683], Fresh[3682], Fresh[3681], Fresh[3680]}), .outt ({new_AGEMA_signal_1868, new_AGEMA_signal_1867, new_AGEMA_signal_1866, n2391}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2554 ( .ina ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2505}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[3699], Fresh[3698], Fresh[3697], Fresh[3696], Fresh[3695], Fresh[3694], Fresh[3693], Fresh[3692], Fresh[3691], Fresh[3690]}), .outt ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, new_AGEMA_signal_2340, n2390}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2559 ( .ina ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}), .inb ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, new_AGEMA_signal_1428, n2700}), .clk ( clk ), .rnd ({Fresh[3709], Fresh[3708], Fresh[3707], Fresh[3706], Fresh[3705], Fresh[3704], Fresh[3703], Fresh[3702], Fresh[3701], Fresh[3700]}), .outt ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, new_AGEMA_signal_1869, n2396}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2562 ( .ina ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .inb ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, new_AGEMA_signal_1809, n2438}), .clk ( clk ), .rnd ({Fresh[3719], Fresh[3718], Fresh[3717], Fresh[3716], Fresh[3715], Fresh[3714], Fresh[3713], Fresh[3712], Fresh[3711], Fresh[3710]}), .outt ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, new_AGEMA_signal_2343, n2406}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2565 ( .ina ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, n2594}), .inb ({new_AGEMA_signal_1436, new_AGEMA_signal_1435, new_AGEMA_signal_1434, n2402}), .clk ( clk ), .rnd ({Fresh[3729], Fresh[3728], Fresh[3727], Fresh[3726], Fresh[3725], Fresh[3724], Fresh[3723], Fresh[3722], Fresh[3721], Fresh[3720]}), .outt ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, new_AGEMA_signal_1872, n2403}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2569 ( .ina ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, new_AGEMA_signal_1650, n2407}), .inb ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .clk ( clk ), .rnd ({Fresh[3739], Fresh[3738], Fresh[3737], Fresh[3736], Fresh[3735], Fresh[3734], Fresh[3733], Fresh[3732], Fresh[3731], Fresh[3730]}), .outt ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, new_AGEMA_signal_2349, n2408}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2573 ( .ina ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, new_AGEMA_signal_1551, n2412}), .inb ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, n2777}), .clk ( clk ), .rnd ({Fresh[3749], Fresh[3748], Fresh[3747], Fresh[3746], Fresh[3745], Fresh[3744], Fresh[3743], Fresh[3742], Fresh[3741], Fresh[3740]}), .outt ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, new_AGEMA_signal_2352, n2574}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2574 ( .ina ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .inb ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}), .clk ( clk ), .rnd ({Fresh[3759], Fresh[3758], Fresh[3757], Fresh[3756], Fresh[3755], Fresh[3754], Fresh[3753], Fresh[3752], Fresh[3751], Fresh[3750]}), .outt ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, new_AGEMA_signal_1875, n2413}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2577 ( .ina ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, new_AGEMA_signal_1425, n2415}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[3769], Fresh[3768], Fresh[3767], Fresh[3766], Fresh[3765], Fresh[3764], Fresh[3763], Fresh[3762], Fresh[3761], Fresh[3760]}), .outt ({new_AGEMA_signal_1880, new_AGEMA_signal_1879, new_AGEMA_signal_1878, n2416}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2586 ( .ina ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, new_AGEMA_signal_1881, n2428}), .inb ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .clk ( clk ), .rnd ({Fresh[3779], Fresh[3778], Fresh[3777], Fresh[3776], Fresh[3775], Fresh[3774], Fresh[3773], Fresh[3772], Fresh[3771], Fresh[3770]}), .outt ({new_AGEMA_signal_2360, new_AGEMA_signal_2359, new_AGEMA_signal_2358, n2433}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2587 ( .ina ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, n2429}), .clk ( clk ), .rnd ({Fresh[3789], Fresh[3788], Fresh[3787], Fresh[3786], Fresh[3785], Fresh[3784], Fresh[3783], Fresh[3782], Fresh[3781], Fresh[3780]}), .outt ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, new_AGEMA_signal_2361, n2689}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2591 ( .ina ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, n2647}), .inb ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}), .clk ( clk ), .rnd ({Fresh[3799], Fresh[3798], Fresh[3797], Fresh[3796], Fresh[3795], Fresh[3794], Fresh[3793], Fresh[3792], Fresh[3791], Fresh[3790]}), .outt ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, new_AGEMA_signal_1887, n2434}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2595 ( .ina ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, new_AGEMA_signal_1809, n2438}), .inb ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, n2483}), .clk ( clk ), .rnd ({Fresh[3809], Fresh[3808], Fresh[3807], Fresh[3806], Fresh[3805], Fresh[3804], Fresh[3803], Fresh[3802], Fresh[3801], Fresh[3800]}), .outt ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, new_AGEMA_signal_2367, n2439}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2598 ( .ina ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .inb ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, new_AGEMA_signal_1779, n2540}), .clk ( clk ), .rnd ({Fresh[3819], Fresh[3818], Fresh[3817], Fresh[3816], Fresh[3815], Fresh[3814], Fresh[3813], Fresh[3812], Fresh[3811], Fresh[3810]}), .outt ({new_AGEMA_signal_2372, new_AGEMA_signal_2371, new_AGEMA_signal_2370, n2445}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2600 ( .ina ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, n2690}), .inb ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, new_AGEMA_signal_1890, n2443}), .clk ( clk ), .rnd ({Fresh[3829], Fresh[3828], Fresh[3827], Fresh[3826], Fresh[3825], Fresh[3824], Fresh[3823], Fresh[3822], Fresh[3821], Fresh[3820]}), .outt ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2373, n2444}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2602 ( .ina ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .inb ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, new_AGEMA_signal_1740, n2446}), .clk ( clk ), .rnd ({Fresh[3839], Fresh[3838], Fresh[3837], Fresh[3836], Fresh[3835], Fresh[3834], Fresh[3833], Fresh[3832], Fresh[3831], Fresh[3830]}), .outt ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, new_AGEMA_signal_2376, n2447}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2607 ( .ina ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}), .inb ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, new_AGEMA_signal_1893, n2693}), .clk ( clk ), .rnd ({Fresh[3849], Fresh[3848], Fresh[3847], Fresh[3846], Fresh[3845], Fresh[3844], Fresh[3843], Fresh[3842], Fresh[3841], Fresh[3840]}), .outt ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, new_AGEMA_signal_2379, n2454}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2617 ( .ina ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .inb ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443, n2464}), .clk ( clk ), .rnd ({Fresh[3859], Fresh[3858], Fresh[3857], Fresh[3856], Fresh[3855], Fresh[3854], Fresh[3853], Fresh[3852], Fresh[3851], Fresh[3850]}), .outt ({new_AGEMA_signal_1898, new_AGEMA_signal_1897, new_AGEMA_signal_1896, n2465}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2622 ( .ina ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .inb ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, n2576}), .clk ( clk ), .rnd ({Fresh[3869], Fresh[3868], Fresh[3867], Fresh[3866], Fresh[3865], Fresh[3864], Fresh[3863], Fresh[3862], Fresh[3861], Fresh[3860]}), .outt ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, new_AGEMA_signal_1899, n2470}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2626 ( .ina ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, new_AGEMA_signal_1449, n2473}), .inb ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, new_AGEMA_signal_1452, n2472}), .clk ( clk ), .rnd ({Fresh[3879], Fresh[3878], Fresh[3877], Fresh[3876], Fresh[3875], Fresh[3874], Fresh[3873], Fresh[3872], Fresh[3871], Fresh[3870]}), .outt ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, new_AGEMA_signal_1902, n2476}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2633 ( .ina ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .inb ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, new_AGEMA_signal_1905, n2480}), .clk ( clk ), .rnd ({Fresh[3889], Fresh[3888], Fresh[3887], Fresh[3886], Fresh[3885], Fresh[3884], Fresh[3883], Fresh[3882], Fresh[3881], Fresh[3880]}), .outt ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, new_AGEMA_signal_2388, n2481}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2639 ( .ina ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .inb ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .rnd ({Fresh[3899], Fresh[3898], Fresh[3897], Fresh[3896], Fresh[3895], Fresh[3894], Fresh[3893], Fresh[3892], Fresh[3891], Fresh[3890]}), .outt ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, new_AGEMA_signal_1911, n2486}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2642 ( .ina ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}), .inb ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, new_AGEMA_signal_1458, n2488}), .clk ( clk ), .rnd ({Fresh[3909], Fresh[3908], Fresh[3907], Fresh[3906], Fresh[3905], Fresh[3904], Fresh[3903], Fresh[3902], Fresh[3901], Fresh[3900]}), .outt ({new_AGEMA_signal_1916, new_AGEMA_signal_1915, new_AGEMA_signal_1914, n2489}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2645 ( .ina ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2493}), .inb ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}), .clk ( clk ), .rnd ({Fresh[3919], Fresh[3918], Fresh[3917], Fresh[3916], Fresh[3915], Fresh[3914], Fresh[3913], Fresh[3912], Fresh[3911], Fresh[3910]}), .outt ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, new_AGEMA_signal_1917, n2497}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2646 ( .ina ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, n2577}), .inb ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, new_AGEMA_signal_1428, n2700}), .clk ( clk ), .rnd ({Fresh[3929], Fresh[3928], Fresh[3927], Fresh[3926], Fresh[3925], Fresh[3924], Fresh[3923], Fresh[3922], Fresh[3921], Fresh[3920]}), .outt ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, new_AGEMA_signal_1920, n2495}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2647 ( .ina ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .inb ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2625}), .clk ( clk ), .rnd ({Fresh[3939], Fresh[3938], Fresh[3937], Fresh[3936], Fresh[3935], Fresh[3934], Fresh[3933], Fresh[3932], Fresh[3931], Fresh[3930]}), .outt ({new_AGEMA_signal_2396, new_AGEMA_signal_2395, new_AGEMA_signal_2394, n2494}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2650 ( .ina ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .inb ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[3949], Fresh[3948], Fresh[3947], Fresh[3946], Fresh[3945], Fresh[3944], Fresh[3943], Fresh[3942], Fresh[3941], Fresh[3940]}), .outt ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, new_AGEMA_signal_1923, n2499}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2653 ( .ina ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, n2674}), .clk ( clk ), .rnd ({Fresh[3959], Fresh[3958], Fresh[3957], Fresh[3956], Fresh[3955], Fresh[3954], Fresh[3953], Fresh[3952], Fresh[3951], Fresh[3950]}), .outt ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, new_AGEMA_signal_2787, n2503}) ) ;
    mux2_HPC1 #(.security_order(3), .pipeline(0)) U2655 ( .ins ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .inb ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2505}), .ina ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .rnd ({Fresh[3969], Fresh[3968], Fresh[3967], Fresh[3966], Fresh[3965], Fresh[3964], Fresh[3963], Fresh[3962], Fresh[3961], Fresh[3960]}), .outt ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, new_AGEMA_signal_2397, n2506}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2662 ( .ina ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1539, n2662}), .inb ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .rnd ({Fresh[3979], Fresh[3978], Fresh[3977], Fresh[3976], Fresh[3975], Fresh[3974], Fresh[3973], Fresh[3972], Fresh[3971], Fresh[3970]}), .outt ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, new_AGEMA_signal_2400, n2518}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2663 ( .ina ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, n2720}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[3989], Fresh[3988], Fresh[3987], Fresh[3986], Fresh[3985], Fresh[3984], Fresh[3983], Fresh[3982], Fresh[3981], Fresh[3980]}), .outt ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, new_AGEMA_signal_2790, n2517}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2666 ( .ina ({new_AGEMA_signal_1928, new_AGEMA_signal_1927, new_AGEMA_signal_1926, n2520}), .inb ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .clk ( clk ), .rnd ({Fresh[3999], Fresh[3998], Fresh[3997], Fresh[3996], Fresh[3995], Fresh[3994], Fresh[3993], Fresh[3992], Fresh[3991], Fresh[3990]}), .outt ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, new_AGEMA_signal_2403, n2523}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2668 ( .ina ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, new_AGEMA_signal_1800, n2774}), .inb ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, new_AGEMA_signal_1461, n2521}), .clk ( clk ), .rnd ({Fresh[4009], Fresh[4008], Fresh[4007], Fresh[4006], Fresh[4005], Fresh[4004], Fresh[4003], Fresh[4002], Fresh[4001], Fresh[4000]}), .outt ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, new_AGEMA_signal_2406, n2522}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2675 ( .ina ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .inb ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, new_AGEMA_signal_1929, n2531}), .clk ( clk ), .rnd ({Fresh[4019], Fresh[4018], Fresh[4017], Fresh[4016], Fresh[4015], Fresh[4014], Fresh[4013], Fresh[4012], Fresh[4011], Fresh[4010]}), .outt ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2409, n2532}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2677 ( .ina ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .inb ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .clk ( clk ), .rnd ({Fresh[4029], Fresh[4028], Fresh[4027], Fresh[4026], Fresh[4025], Fresh[4024], Fresh[4023], Fresh[4022], Fresh[4021], Fresh[4020]}), .outt ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, new_AGEMA_signal_2412, n2534}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2681 ( .ina ({new_AGEMA_signal_1214, new_AGEMA_signal_1213, new_AGEMA_signal_1212, n2541}), .inb ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, new_AGEMA_signal_1779, n2540}), .clk ( clk ), .rnd ({Fresh[4039], Fresh[4038], Fresh[4037], Fresh[4036], Fresh[4035], Fresh[4034], Fresh[4033], Fresh[4032], Fresh[4031], Fresh[4030]}), .outt ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, new_AGEMA_signal_2415, n2542}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2683 ( .ina ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2545}), .inb ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, new_AGEMA_signal_1353, n2544}), .clk ( clk ), .rnd ({Fresh[4049], Fresh[4048], Fresh[4047], Fresh[4046], Fresh[4045], Fresh[4044], Fresh[4043], Fresh[4042], Fresh[4041], Fresh[4040]}), .outt ({new_AGEMA_signal_1934, new_AGEMA_signal_1933, new_AGEMA_signal_1932, n2546}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2687 ( .ina ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, new_AGEMA_signal_1272, n2673}), .inb ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .clk ( clk ), .rnd ({Fresh[4059], Fresh[4058], Fresh[4057], Fresh[4056], Fresh[4055], Fresh[4054], Fresh[4053], Fresh[4052], Fresh[4051], Fresh[4050]}), .outt ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, new_AGEMA_signal_2421, n2551}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2690 ( .ina ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, new_AGEMA_signal_1935, n2553}), .inb ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2679}), .clk ( clk ), .rnd ({Fresh[4069], Fresh[4068], Fresh[4067], Fresh[4066], Fresh[4065], Fresh[4064], Fresh[4063], Fresh[4062], Fresh[4061], Fresh[4060]}), .outt ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, new_AGEMA_signal_2424, n2558}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2692 ( .ina ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, new_AGEMA_signal_1719, n2555}), .inb ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, new_AGEMA_signal_1938, n2554}), .clk ( clk ), .rnd ({Fresh[4079], Fresh[4078], Fresh[4077], Fresh[4076], Fresh[4075], Fresh[4074], Fresh[4073], Fresh[4072], Fresh[4071], Fresh[4070]}), .outt ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, n2556}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2696 ( .ina ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, new_AGEMA_signal_1770, n2561}), .inb ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, new_AGEMA_signal_1464, n2560}), .clk ( clk ), .rnd ({Fresh[4089], Fresh[4088], Fresh[4087], Fresh[4086], Fresh[4085], Fresh[4084], Fresh[4083], Fresh[4082], Fresh[4081], Fresh[4080]}), .outt ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, new_AGEMA_signal_2430, n2566}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2697 ( .ina ({new_AGEMA_signal_1040, new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2699}), .inb ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, new_AGEMA_signal_1674, n2562}), .clk ( clk ), .rnd ({Fresh[4099], Fresh[4098], Fresh[4097], Fresh[4096], Fresh[4095], Fresh[4094], Fresh[4093], Fresh[4092], Fresh[4091], Fresh[4090]}), .outt ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2433, n2715}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2703 ( .ina ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, n2572}), .inb ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, n2571}), .clk ( clk ), .rnd ({Fresh[4109], Fresh[4108], Fresh[4107], Fresh[4106], Fresh[4105], Fresh[4104], Fresh[4103], Fresh[4102], Fresh[4101], Fresh[4100]}), .outt ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, new_AGEMA_signal_2436, n2573}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2705 ( .ina ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .inb ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, new_AGEMA_signal_1635, n2754}), .clk ( clk ), .rnd ({Fresh[4119], Fresh[4118], Fresh[4117], Fresh[4116], Fresh[4115], Fresh[4114], Fresh[4113], Fresh[4112], Fresh[4111], Fresh[4110]}), .outt ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, new_AGEMA_signal_2439, n2585}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2706 ( .ina ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .inb ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .clk ( clk ), .rnd ({Fresh[4129], Fresh[4128], Fresh[4127], Fresh[4126], Fresh[4125], Fresh[4124], Fresh[4123], Fresh[4122], Fresh[4121], Fresh[4120]}), .outt ({new_AGEMA_signal_1946, new_AGEMA_signal_1945, new_AGEMA_signal_1944, n2581}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2707 ( .ina ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, new_AGEMA_signal_1497, n2575}), .inb ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .rnd ({Fresh[4139], Fresh[4138], Fresh[4137], Fresh[4136], Fresh[4135], Fresh[4134], Fresh[4133], Fresh[4132], Fresh[4131], Fresh[4130]}), .outt ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, new_AGEMA_signal_2442, n2579}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2708 ( .ina ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, n2577}), .inb ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, n2576}), .clk ( clk ), .rnd ({Fresh[4149], Fresh[4148], Fresh[4147], Fresh[4146], Fresh[4145], Fresh[4144], Fresh[4143], Fresh[4142], Fresh[4141], Fresh[4140]}), .outt ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, new_AGEMA_signal_1947, n2578}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2711 ( .ina ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2625}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[4159], Fresh[4158], Fresh[4157], Fresh[4156], Fresh[4155], Fresh[4154], Fresh[4153], Fresh[4152], Fresh[4151], Fresh[4150]}), .outt ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, new_AGEMA_signal_2445, n2582}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2715 ( .ina ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, n2587}), .inb ({new_AGEMA_signal_1952, new_AGEMA_signal_1951, new_AGEMA_signal_1950, n2586}), .clk ( clk ), .rnd ({Fresh[4169], Fresh[4168], Fresh[4167], Fresh[4166], Fresh[4165], Fresh[4164], Fresh[4163], Fresh[4162], Fresh[4161], Fresh[4160]}), .outt ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, new_AGEMA_signal_2448, n2588}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2719 ( .ina ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, n2594}), .inb ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .clk ( clk ), .rnd ({Fresh[4179], Fresh[4178], Fresh[4177], Fresh[4176], Fresh[4175], Fresh[4174], Fresh[4173], Fresh[4172], Fresh[4171], Fresh[4170]}), .outt ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, new_AGEMA_signal_1953, n2607}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2722 ( .ina ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, new_AGEMA_signal_1467, n2597}), .inb ({new_AGEMA_signal_1958, new_AGEMA_signal_1957, new_AGEMA_signal_1956, n2596}), .clk ( clk ), .rnd ({Fresh[4189], Fresh[4188], Fresh[4187], Fresh[4186], Fresh[4185], Fresh[4184], Fresh[4183], Fresh[4182], Fresh[4181], Fresh[4180]}), .outt ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, new_AGEMA_signal_2451, n2605}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2724 ( .ina ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, new_AGEMA_signal_1959, n2598}), .inb ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .clk ( clk ), .rnd ({Fresh[4199], Fresh[4198], Fresh[4197], Fresh[4196], Fresh[4195], Fresh[4194], Fresh[4193], Fresh[4192], Fresh[4191], Fresh[4190]}), .outt ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, n2603}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2726 ( .ina ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, n2599}), .inb ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, n2777}), .clk ( clk ), .rnd ({Fresh[4209], Fresh[4208], Fresh[4207], Fresh[4206], Fresh[4205], Fresh[4204], Fresh[4203], Fresh[4202], Fresh[4201], Fresh[4200]}), .outt ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, new_AGEMA_signal_1470, n2601}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2733 ( .ina ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, new_AGEMA_signal_1965, n2610}), .inb ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .clk ( clk ), .rnd ({Fresh[4219], Fresh[4218], Fresh[4217], Fresh[4216], Fresh[4215], Fresh[4214], Fresh[4213], Fresh[4212], Fresh[4211], Fresh[4210]}), .outt ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, new_AGEMA_signal_2457, n2620}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2736 ( .ina ({new_AGEMA_signal_1970, new_AGEMA_signal_1969, new_AGEMA_signal_1968, n2614}), .inb ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, new_AGEMA_signal_1971, n2613}), .clk ( clk ), .rnd ({Fresh[4229], Fresh[4228], Fresh[4227], Fresh[4226], Fresh[4225], Fresh[4224], Fresh[4223], Fresh[4222], Fresh[4221], Fresh[4220]}), .outt ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, new_AGEMA_signal_2460, n2618}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2743 ( .ina ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .inb ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2625}), .clk ( clk ), .rnd ({Fresh[4239], Fresh[4238], Fresh[4237], Fresh[4236], Fresh[4235], Fresh[4234], Fresh[4233], Fresh[4232], Fresh[4231], Fresh[4230]}), .outt ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, new_AGEMA_signal_2463, n2626}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2746 ( .ina ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2631}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[4249], Fresh[4248], Fresh[4247], Fresh[4246], Fresh[4245], Fresh[4244], Fresh[4243], Fresh[4242], Fresh[4241], Fresh[4240]}), .outt ({new_AGEMA_signal_1976, new_AGEMA_signal_1975, new_AGEMA_signal_1974, n2632}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2752 ( .ina ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, new_AGEMA_signal_1977, n2784}), .inb ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, new_AGEMA_signal_1338, n2642}), .clk ( clk ), .rnd ({Fresh[4259], Fresh[4258], Fresh[4257], Fresh[4256], Fresh[4255], Fresh[4254], Fresh[4253], Fresh[4252], Fresh[4251], Fresh[4250]}), .outt ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, new_AGEMA_signal_2466, n2644}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2754 ( .ina ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .inb ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, n2645}), .clk ( clk ), .rnd ({Fresh[4269], Fresh[4268], Fresh[4267], Fresh[4266], Fresh[4265], Fresh[4264], Fresh[4263], Fresh[4262], Fresh[4261], Fresh[4260]}), .outt ({new_AGEMA_signal_1982, new_AGEMA_signal_1981, new_AGEMA_signal_1980, n2646}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2758 ( .ina ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .inb ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, new_AGEMA_signal_1479, n2650}), .clk ( clk ), .rnd ({Fresh[4279], Fresh[4278], Fresh[4277], Fresh[4276], Fresh[4275], Fresh[4274], Fresh[4273], Fresh[4272], Fresh[4271], Fresh[4270]}), .outt ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, new_AGEMA_signal_1983, n2653}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2760 ( .ina ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, n2777}), .inb ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, n2654}), .clk ( clk ), .rnd ({Fresh[4289], Fresh[4288], Fresh[4287], Fresh[4286], Fresh[4285], Fresh[4284], Fresh[4283], Fresh[4282], Fresh[4281], Fresh[4280]}), .outt ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, new_AGEMA_signal_2472, n2655}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2764 ( .ina ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1539, n2662}), .inb ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}), .clk ( clk ), .rnd ({Fresh[4299], Fresh[4298], Fresh[4297], Fresh[4296], Fresh[4295], Fresh[4294], Fresh[4293], Fresh[4292], Fresh[4291], Fresh[4290]}), .outt ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, new_AGEMA_signal_2475, n2663}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2770 ( .ina ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, new_AGEMA_signal_1272, n2673}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[4309], Fresh[4308], Fresh[4307], Fresh[4306], Fresh[4305], Fresh[4304], Fresh[4303], Fresh[4302], Fresh[4301], Fresh[4300]}), .outt ({new_AGEMA_signal_1988, new_AGEMA_signal_1987, new_AGEMA_signal_1986, n2675}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2772 ( .ina ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, n2677}), .inb ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, new_AGEMA_signal_1245, n2676}), .clk ( clk ), .rnd ({Fresh[4319], Fresh[4318], Fresh[4317], Fresh[4316], Fresh[4315], Fresh[4314], Fresh[4313], Fresh[4312], Fresh[4311], Fresh[4310]}), .outt ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, new_AGEMA_signal_1989, n2678}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2780 ( .ina ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, n2690}), .inb ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .clk ( clk ), .rnd ({Fresh[4329], Fresh[4328], Fresh[4327], Fresh[4326], Fresh[4325], Fresh[4324], Fresh[4323], Fresh[4322], Fresh[4321], Fresh[4320]}), .outt ({new_AGEMA_signal_1994, new_AGEMA_signal_1993, new_AGEMA_signal_1992, n2691}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2782 ( .ina ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .inb ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, new_AGEMA_signal_1893, n2693}), .clk ( clk ), .rnd ({Fresh[4339], Fresh[4338], Fresh[4337], Fresh[4336], Fresh[4335], Fresh[4334], Fresh[4333], Fresh[4332], Fresh[4331], Fresh[4330]}), .outt ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, new_AGEMA_signal_2481, n2695}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2785 ( .ina ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, new_AGEMA_signal_1428, n2700}), .inb ({new_AGEMA_signal_1040, new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2699}), .clk ( clk ), .rnd ({Fresh[4349], Fresh[4348], Fresh[4347], Fresh[4346], Fresh[4345], Fresh[4344], Fresh[4343], Fresh[4342], Fresh[4341], Fresh[4340]}), .outt ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, new_AGEMA_signal_1995, n2701}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2791 ( .ina ({new_AGEMA_signal_2000, new_AGEMA_signal_1999, new_AGEMA_signal_1998, n2711}), .inb ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, new_AGEMA_signal_2001, n2710}), .clk ( clk ), .rnd ({Fresh[4359], Fresh[4358], Fresh[4357], Fresh[4356], Fresh[4355], Fresh[4354], Fresh[4353], Fresh[4352], Fresh[4351], Fresh[4350]}), .outt ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, new_AGEMA_signal_2484, n2717}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2796 ( .ina ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, n2720}), .inb ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .rnd ({Fresh[4369], Fresh[4368], Fresh[4367], Fresh[4366], Fresh[4365], Fresh[4364], Fresh[4363], Fresh[4362], Fresh[4361], Fresh[4360]}), .outt ({new_AGEMA_signal_2846, new_AGEMA_signal_2845, new_AGEMA_signal_2844, n2729}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2798 ( .ina ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .inb ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, new_AGEMA_signal_1485, n2722}), .clk ( clk ), .rnd ({Fresh[4379], Fresh[4378], Fresh[4377], Fresh[4376], Fresh[4375], Fresh[4374], Fresh[4373], Fresh[4372], Fresh[4371], Fresh[4370]}), .outt ({new_AGEMA_signal_2006, new_AGEMA_signal_2005, new_AGEMA_signal_2004, n2727}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2803 ( .ina ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .inb ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, new_AGEMA_signal_1656, n2731}), .clk ( clk ), .rnd ({Fresh[4389], Fresh[4388], Fresh[4387], Fresh[4386], Fresh[4385], Fresh[4384], Fresh[4383], Fresh[4382], Fresh[4381], Fresh[4380]}), .outt ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, new_AGEMA_signal_2490, n2733}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2807 ( .ina ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, new_AGEMA_signal_1101, n2739}), .inb ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, new_AGEMA_signal_2010, n2738}), .clk ( clk ), .rnd ({Fresh[4399], Fresh[4398], Fresh[4397], Fresh[4396], Fresh[4395], Fresh[4394], Fresh[4393], Fresh[4392], Fresh[4391], Fresh[4390]}), .outt ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, new_AGEMA_signal_2493, n2740}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2812 ( .ina ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, new_AGEMA_signal_1380, n2748}), .inb ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .clk ( clk ), .rnd ({Fresh[4409], Fresh[4408], Fresh[4407], Fresh[4406], Fresh[4405], Fresh[4404], Fresh[4403], Fresh[4402], Fresh[4401], Fresh[4400]}), .outt ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, new_AGEMA_signal_2013, n2749}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2815 ( .ina ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, new_AGEMA_signal_1635, n2754}), .inb ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}), .clk ( clk ), .rnd ({Fresh[4419], Fresh[4418], Fresh[4417], Fresh[4416], Fresh[4415], Fresh[4414], Fresh[4413], Fresh[4412], Fresh[4411], Fresh[4410]}), .outt ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, new_AGEMA_signal_2499, n2757}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2816 ( .ina ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, new_AGEMA_signal_1206, n2755}), .inb ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2772}), .clk ( clk ), .rnd ({Fresh[4429], Fresh[4428], Fresh[4427], Fresh[4426], Fresh[4425], Fresh[4424], Fresh[4423], Fresh[4422], Fresh[4421], Fresh[4420]}), .outt ({new_AGEMA_signal_2018, new_AGEMA_signal_2017, new_AGEMA_signal_2016, n2756}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2819 ( .ina ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}), .inb ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .clk ( clk ), .rnd ({Fresh[4439], Fresh[4438], Fresh[4437], Fresh[4436], Fresh[4435], Fresh[4434], Fresh[4433], Fresh[4432], Fresh[4431], Fresh[4430]}), .outt ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, new_AGEMA_signal_2502, n2762}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2823 ( .ina ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .inb ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, new_AGEMA_signal_2019, n2768}), .clk ( clk ), .rnd ({Fresh[4449], Fresh[4448], Fresh[4447], Fresh[4446], Fresh[4445], Fresh[4444], Fresh[4443], Fresh[4442], Fresh[4441], Fresh[4440]}), .outt ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, new_AGEMA_signal_2505, n2770}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2825 ( .ina ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, new_AGEMA_signal_1668, n2773}), .inb ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2772}), .clk ( clk ), .rnd ({Fresh[4459], Fresh[4458], Fresh[4457], Fresh[4456], Fresh[4455], Fresh[4454], Fresh[4453], Fresh[4452], Fresh[4451], Fresh[4450]}), .outt ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, new_AGEMA_signal_2508, n2776}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2826 ( .ina ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, new_AGEMA_signal_1800, n2774}), .inb ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .rnd ({Fresh[4469], Fresh[4468], Fresh[4467], Fresh[4466], Fresh[4465], Fresh[4464], Fresh[4463], Fresh[4462], Fresh[4461], Fresh[4460]}), .outt ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, new_AGEMA_signal_2511, n2775}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2830 ( .ina ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, new_AGEMA_signal_1488, n2782}), .inb ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, new_AGEMA_signal_1491, n2781}), .clk ( clk ), .rnd ({Fresh[4479], Fresh[4478], Fresh[4477], Fresh[4476], Fresh[4475], Fresh[4474], Fresh[4473], Fresh[4472], Fresh[4471], Fresh[4470]}), .outt ({new_AGEMA_signal_2024, new_AGEMA_signal_2023, new_AGEMA_signal_2022, n2783}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2836 ( .ina ({new_AGEMA_signal_2030, new_AGEMA_signal_2029, new_AGEMA_signal_2028, n2794}), .inb ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, new_AGEMA_signal_2031, n2793}), .clk ( clk ), .rnd ({Fresh[4489], Fresh[4488], Fresh[4487], Fresh[4486], Fresh[4485], Fresh[4484], Fresh[4483], Fresh[4482], Fresh[4481], Fresh[4480]}), .outt ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, new_AGEMA_signal_2517, n2795}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2845 ( .ina ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, new_AGEMA_signal_2034, n2812}), .inb ({new_AGEMA_signal_1700, new_AGEMA_signal_1699, new_AGEMA_signal_1698, n2811}), .clk ( clk ), .rnd ({Fresh[4499], Fresh[4498], Fresh[4497], Fresh[4496], Fresh[4495], Fresh[4494], Fresh[4493], Fresh[4492], Fresh[4491], Fresh[4490]}), .outt ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, new_AGEMA_signal_2520, n2814}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2848 ( .ina ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .inb ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .rnd ({Fresh[4509], Fresh[4508], Fresh[4507], Fresh[4506], Fresh[4505], Fresh[4504], Fresh[4503], Fresh[4502], Fresh[4501], Fresh[4500]}), .outt ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, new_AGEMA_signal_2037, n2819}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1968 ( .ina ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, new_AGEMA_signal_2043, n1924}), .inb ({new_AGEMA_signal_2048, new_AGEMA_signal_2047, new_AGEMA_signal_2046, n1923}), .clk ( clk ), .rnd ({Fresh[4519], Fresh[4518], Fresh[4517], Fresh[4516], Fresh[4515], Fresh[4514], Fresh[4513], Fresh[4512], Fresh[4511], Fresh[4510]}), .outt ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, new_AGEMA_signal_2526, n1936}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1982 ( .ina ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, new_AGEMA_signal_1206, n2755}), .inb ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, new_AGEMA_signal_2049, n1927}), .clk ( clk ), .rnd ({Fresh[4529], Fresh[4528], Fresh[4527], Fresh[4526], Fresh[4525], Fresh[4524], Fresh[4523], Fresh[4522], Fresh[4521], Fresh[4520]}), .outt ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, new_AGEMA_signal_2529, n1928}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U1994 ( .ina ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, new_AGEMA_signal_1512, n2151}), .inb ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, new_AGEMA_signal_2052, n1929}), .clk ( clk ), .rnd ({Fresh[4539], Fresh[4538], Fresh[4537], Fresh[4536], Fresh[4535], Fresh[4534], Fresh[4533], Fresh[4532], Fresh[4531], Fresh[4530]}), .outt ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, new_AGEMA_signal_2532, n1931}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2012 ( .ina ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, new_AGEMA_signal_2055, n2665}), .inb ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, new_AGEMA_signal_2058, n1938}), .clk ( clk ), .rnd ({Fresh[4549], Fresh[4548], Fresh[4547], Fresh[4546], Fresh[4545], Fresh[4544], Fresh[4543], Fresh[4542], Fresh[4541], Fresh[4540]}), .outt ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, new_AGEMA_signal_2535, n1939}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2024 ( .ina ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, new_AGEMA_signal_2061, n2235}), .inb ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, new_AGEMA_signal_1527, n1943}), .clk ( clk ), .rnd ({Fresh[4559], Fresh[4558], Fresh[4557], Fresh[4556], Fresh[4555], Fresh[4554], Fresh[4553], Fresh[4552], Fresh[4551], Fresh[4550]}), .outt ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, new_AGEMA_signal_2538, n1948}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2032 ( .ina ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, new_AGEMA_signal_1530, n1946}), .inb ({new_AGEMA_signal_2066, new_AGEMA_signal_2065, new_AGEMA_signal_2064, n1945}), .clk ( clk ), .rnd ({Fresh[4569], Fresh[4568], Fresh[4567], Fresh[4566], Fresh[4565], Fresh[4564], Fresh[4563], Fresh[4562], Fresh[4561], Fresh[4560]}), .outt ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, new_AGEMA_signal_2541, n1947}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2041 ( .ina ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .inb ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, new_AGEMA_signal_2070, n1951}), .clk ( clk ), .rnd ({Fresh[4579], Fresh[4578], Fresh[4577], Fresh[4576], Fresh[4575], Fresh[4574], Fresh[4573], Fresh[4572], Fresh[4571], Fresh[4570]}), .outt ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, new_AGEMA_signal_2544, n1954}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2049 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, new_AGEMA_signal_2073, n1952}), .clk ( clk ), .rnd ({Fresh[4589], Fresh[4588], Fresh[4587], Fresh[4586], Fresh[4585], Fresh[4584], Fresh[4583], Fresh[4582], Fresh[4581], Fresh[4580]}), .outt ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, new_AGEMA_signal_2547, n1953}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2058 ( .ina ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, n2687}), .clk ( clk ), .rnd ({Fresh[4599], Fresh[4598], Fresh[4597], Fresh[4596], Fresh[4595], Fresh[4594], Fresh[4593], Fresh[4592], Fresh[4591], Fresh[4590]}), .outt ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, new_AGEMA_signal_2550, n2658}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2065 ( .ina ({new_AGEMA_signal_1115, new_AGEMA_signal_1114, new_AGEMA_signal_1113, n1964}), .inb ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, new_AGEMA_signal_1545, n1963}), .clk ( clk ), .rnd ({Fresh[4609], Fresh[4608], Fresh[4607], Fresh[4606], Fresh[4605], Fresh[4604], Fresh[4603], Fresh[4602], Fresh[4601], Fresh[4600]}), .outt ({new_AGEMA_signal_2084, new_AGEMA_signal_2083, new_AGEMA_signal_2082, n1965}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2078 ( .ina ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, new_AGEMA_signal_1272, n2673}), .inb ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, new_AGEMA_signal_2556, n1968}), .clk ( clk ), .rnd ({Fresh[4619], Fresh[4618], Fresh[4617], Fresh[4616], Fresh[4615], Fresh[4614], Fresh[4613], Fresh[4612], Fresh[4611], Fresh[4610]}), .outt ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, new_AGEMA_signal_2889, n1970}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2084 ( .ina ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, new_AGEMA_signal_2091, n2684}), .inb ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, new_AGEMA_signal_1557, n2359}), .clk ( clk ), .rnd ({Fresh[4629], Fresh[4628], Fresh[4627], Fresh[4626], Fresh[4625], Fresh[4624], Fresh[4623], Fresh[4622], Fresh[4621], Fresh[4620]}), .outt ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, new_AGEMA_signal_2559, n1969}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2093 ( .ina ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, new_AGEMA_signal_2094, n1972}), .inb ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, new_AGEMA_signal_1563, n1971}), .clk ( clk ), .rnd ({Fresh[4639], Fresh[4638], Fresh[4637], Fresh[4636], Fresh[4635], Fresh[4634], Fresh[4633], Fresh[4632], Fresh[4631], Fresh[4630]}), .outt ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, new_AGEMA_signal_2562, n1978}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2102 ( .ina ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, new_AGEMA_signal_2097, n1974}), .inb ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, new_AGEMA_signal_1569, n1973}), .clk ( clk ), .rnd ({Fresh[4649], Fresh[4648], Fresh[4647], Fresh[4646], Fresh[4645], Fresh[4644], Fresh[4643], Fresh[4642], Fresh[4641], Fresh[4640]}), .outt ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, new_AGEMA_signal_2565, n1975}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2107 ( .ina ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, n2690}), .inb ({new_AGEMA_signal_2102, new_AGEMA_signal_2101, new_AGEMA_signal_2100, n1979}), .clk ( clk ), .rnd ({Fresh[4659], Fresh[4658], Fresh[4657], Fresh[4656], Fresh[4655], Fresh[4654], Fresh[4653], Fresh[4652], Fresh[4651], Fresh[4650]}), .outt ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, new_AGEMA_signal_2568, n1980}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2114 ( .ina ({new_AGEMA_signal_1574, new_AGEMA_signal_1573, new_AGEMA_signal_1572, n1985}), .inb ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, new_AGEMA_signal_1575, n2741}), .clk ( clk ), .rnd ({Fresh[4669], Fresh[4668], Fresh[4667], Fresh[4666], Fresh[4665], Fresh[4664], Fresh[4663], Fresh[4662], Fresh[4661], Fresh[4660]}), .outt ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, new_AGEMA_signal_2103, n1986}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2124 ( .ina ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, new_AGEMA_signal_2106, n1994}), .inb ({new_AGEMA_signal_1310, new_AGEMA_signal_1309, new_AGEMA_signal_1308, n1993}), .clk ( clk ), .rnd ({Fresh[4679], Fresh[4678], Fresh[4677], Fresh[4676], Fresh[4675], Fresh[4674], Fresh[4673], Fresh[4672], Fresh[4671], Fresh[4670]}), .outt ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, new_AGEMA_signal_2574, n1997}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2137 ( .ina ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, new_AGEMA_signal_1587, n2241}), .inb ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, new_AGEMA_signal_2112, n2137}), .clk ( clk ), .rnd ({Fresh[4689], Fresh[4688], Fresh[4687], Fresh[4686], Fresh[4685], Fresh[4684], Fresh[4683], Fresh[4682], Fresh[4681], Fresh[4680]}), .outt ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, new_AGEMA_signal_2577, n2012}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2145 ( .ina ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, new_AGEMA_signal_2115, n2006}), .inb ({new_AGEMA_signal_2120, new_AGEMA_signal_2119, new_AGEMA_signal_2118, n2005}), .clk ( clk ), .rnd ({Fresh[4699], Fresh[4698], Fresh[4697], Fresh[4696], Fresh[4695], Fresh[4694], Fresh[4693], Fresh[4692], Fresh[4691], Fresh[4690]}), .outt ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, new_AGEMA_signal_2580, n2007}) ) ;
    mux2_HPC1 #(.security_order(3), .pipeline(0)) U2161 ( .ins ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .inb ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, new_AGEMA_signal_1611, n2020}), .ina ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, new_AGEMA_signal_1017, n2779}), .clk ( clk ), .rnd ({Fresh[4709], Fresh[4708], Fresh[4707], Fresh[4706], Fresh[4705], Fresh[4704], Fresh[4703], Fresh[4702], Fresh[4701], Fresh[4700]}), .outt ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, new_AGEMA_signal_2124, n2021}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2176 ( .ina ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, new_AGEMA_signal_1620, n2290}), .inb ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, new_AGEMA_signal_2130, n2031}), .clk ( clk ), .rnd ({Fresh[4719], Fresh[4718], Fresh[4717], Fresh[4716], Fresh[4715], Fresh[4714], Fresh[4713], Fresh[4712], Fresh[4711], Fresh[4710]}), .outt ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, new_AGEMA_signal_2586, n2032}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2185 ( .ina ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335, n2171}), .inb ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, new_AGEMA_signal_2133, n2040}), .clk ( clk ), .rnd ({Fresh[4729], Fresh[4728], Fresh[4727], Fresh[4726], Fresh[4725], Fresh[4724], Fresh[4723], Fresh[4722], Fresh[4721], Fresh[4720]}), .outt ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, new_AGEMA_signal_2589, n2041}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2189 ( .ina ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, new_AGEMA_signal_2055, n2665}), .inb ({new_AGEMA_signal_1634, new_AGEMA_signal_1633, new_AGEMA_signal_1632, n2042}), .clk ( clk ), .rnd ({Fresh[4739], Fresh[4738], Fresh[4737], Fresh[4736], Fresh[4735], Fresh[4734], Fresh[4733], Fresh[4732], Fresh[4731], Fresh[4730]}), .outt ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, new_AGEMA_signal_2592, n2043}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2194 ( .ina ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, new_AGEMA_signal_1635, n2754}), .inb ({new_AGEMA_signal_2138, new_AGEMA_signal_2137, new_AGEMA_signal_2136, n2045}), .clk ( clk ), .rnd ({Fresh[4749], Fresh[4748], Fresh[4747], Fresh[4746], Fresh[4745], Fresh[4744], Fresh[4743], Fresh[4742], Fresh[4741], Fresh[4740]}), .outt ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, new_AGEMA_signal_2595, n2046}) ) ;
    mux2_HPC1 #(.security_order(3), .pipeline(0)) U2204 ( .ins ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .inb ({new_AGEMA_signal_2144, new_AGEMA_signal_2143, new_AGEMA_signal_2142, n2056}), .ina ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .clk ( clk ), .rnd ({Fresh[4759], Fresh[4758], Fresh[4757], Fresh[4756], Fresh[4755], Fresh[4754], Fresh[4753], Fresh[4752], Fresh[4751], Fresh[4750]}), .outt ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, new_AGEMA_signal_2598, n2058}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2210 ( .ina ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, new_AGEMA_signal_1566, n2535}), .inb ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, new_AGEMA_signal_2145, n2060}), .clk ( clk ), .rnd ({Fresh[4769], Fresh[4768], Fresh[4767], Fresh[4766], Fresh[4765], Fresh[4764], Fresh[4763], Fresh[4762], Fresh[4761], Fresh[4760]}), .outt ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, new_AGEMA_signal_2601, n2063}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2218 ( .ina ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, new_AGEMA_signal_2148, n2066}), .inb ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, new_AGEMA_signal_2151, n2065}), .clk ( clk ), .rnd ({Fresh[4779], Fresh[4778], Fresh[4777], Fresh[4776], Fresh[4775], Fresh[4774], Fresh[4773], Fresh[4772], Fresh[4771], Fresh[4770]}), .outt ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, new_AGEMA_signal_2604, n2652}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2227 ( .ina ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, new_AGEMA_signal_1338, n2642}), .inb ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, new_AGEMA_signal_2157, n2074}), .clk ( clk ), .rnd ({Fresh[4789], Fresh[4788], Fresh[4787], Fresh[4786], Fresh[4785], Fresh[4784], Fresh[4783], Fresh[4782], Fresh[4781], Fresh[4780]}), .outt ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, new_AGEMA_signal_2607, n2076}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2236 ( .ina ({new_AGEMA_signal_1151, new_AGEMA_signal_1150, new_AGEMA_signal_1149, n2721}), .inb ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, new_AGEMA_signal_2160, n2082}), .clk ( clk ), .rnd ({Fresh[4799], Fresh[4798], Fresh[4797], Fresh[4796], Fresh[4795], Fresh[4794], Fresh[4793], Fresh[4792], Fresh[4791], Fresh[4790]}), .outt ({new_AGEMA_signal_2612, new_AGEMA_signal_2611, new_AGEMA_signal_2610, n2105}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2241 ( .ina ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, new_AGEMA_signal_1668, n2773}), .inb ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, new_AGEMA_signal_2163, n2084}), .clk ( clk ), .rnd ({Fresh[4809], Fresh[4808], Fresh[4807], Fresh[4806], Fresh[4805], Fresh[4804], Fresh[4803], Fresh[4802], Fresh[4801], Fresh[4800]}), .outt ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, new_AGEMA_signal_2613, n2099}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2243 ( .ina ({new_AGEMA_signal_2168, new_AGEMA_signal_2167, new_AGEMA_signal_2166, n2085}), .inb ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .clk ( clk ), .rnd ({Fresh[4819], Fresh[4818], Fresh[4817], Fresh[4816], Fresh[4815], Fresh[4814], Fresh[4813], Fresh[4812], Fresh[4811], Fresh[4810]}), .outt ({new_AGEMA_signal_2618, new_AGEMA_signal_2617, new_AGEMA_signal_2616, n2091}) ) ;
    and_HPC1 #(.security_order(3), .pipeline(0)) U2246 ( .ina ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}), .inb ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, new_AGEMA_signal_2169, n2131}), .clk ( clk ), .rnd ({Fresh[4829], Fresh[4828], Fresh[4827], Fresh[4826], Fresh[4825], Fresh[4824], Fresh[4823], Fresh[4822], Fresh[4821], Fresh[4820]}), .outt ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, new_AGEMA_signal_2619, n2090}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2253 ( .ina ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2631}), .inb ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, new_AGEMA_signal_2175, n2330}), .clk ( clk ), .rnd ({Fresh[4839], Fresh[4838], Fresh[4837], Fresh[4836], Fresh[4835], Fresh[4834], Fresh[4833], Fresh[4832], Fresh[4831], Fresh[4830]}), .outt ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, new_AGEMA_signal_2622, n2093}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2262 ( .ina ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}), .inb ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, new_AGEMA_signal_2184, n2160}), .clk ( clk ), .rnd ({Fresh[4849], Fresh[4848], Fresh[4847], Fresh[4846], Fresh[4845], Fresh[4844], Fresh[4843], Fresh[4842], Fresh[4841], Fresh[4840]}), .outt ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, new_AGEMA_signal_2625, n2102}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2266 ( .ina ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, n2504}), .inb ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}), .clk ( clk ), .rnd ({Fresh[4859], Fresh[4858], Fresh[4857], Fresh[4856], Fresh[4855], Fresh[4854], Fresh[4853], Fresh[4852], Fresh[4851], Fresh[4850]}), .outt ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, new_AGEMA_signal_2187, n2106}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2272 ( .ina ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .inb ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, new_AGEMA_signal_2628, n2114}), .clk ( clk ), .rnd ({Fresh[4869], Fresh[4868], Fresh[4867], Fresh[4866], Fresh[4865], Fresh[4864], Fresh[4863], Fresh[4862], Fresh[4861], Fresh[4860]}), .outt ({new_AGEMA_signal_2936, new_AGEMA_signal_2935, new_AGEMA_signal_2934, n2116}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2282 ( .ina ({new_AGEMA_signal_2192, new_AGEMA_signal_2191, new_AGEMA_signal_2190, n2291}), .inb ({new_AGEMA_signal_1694, new_AGEMA_signal_1693, new_AGEMA_signal_1692, n2119}), .clk ( clk ), .rnd ({Fresh[4879], Fresh[4878], Fresh[4877], Fresh[4876], Fresh[4875], Fresh[4874], Fresh[4873], Fresh[4872], Fresh[4871], Fresh[4870]}), .outt ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, new_AGEMA_signal_2631, n2120}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2293 ( .ina ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, new_AGEMA_signal_1701, n2130}), .inb ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, new_AGEMA_signal_1704, n2129}), .clk ( clk ), .rnd ({Fresh[4889], Fresh[4888], Fresh[4887], Fresh[4886], Fresh[4885], Fresh[4884], Fresh[4883], Fresh[4882], Fresh[4881], Fresh[4880]}), .outt ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, new_AGEMA_signal_2193, n2155}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2296 ( .ina ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .inb ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, new_AGEMA_signal_2169, n2131}), .clk ( clk ), .rnd ({Fresh[4899], Fresh[4898], Fresh[4897], Fresh[4896], Fresh[4895], Fresh[4894], Fresh[4893], Fresh[4892], Fresh[4891], Fresh[4890]}), .outt ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, new_AGEMA_signal_2634, n2543}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2299 ( .ina ({new_AGEMA_signal_1712, new_AGEMA_signal_1711, new_AGEMA_signal_1710, n2133}), .inb ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .clk ( clk ), .rnd ({Fresh[4909], Fresh[4908], Fresh[4907], Fresh[4906], Fresh[4905], Fresh[4904], Fresh[4903], Fresh[4902], Fresh[4901], Fresh[4900]}), .outt ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, new_AGEMA_signal_2196, n2134}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2303 ( .ina ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, new_AGEMA_signal_2112, n2137}), .inb ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, new_AGEMA_signal_2199, n2136}), .clk ( clk ), .rnd ({Fresh[4919], Fresh[4918], Fresh[4917], Fresh[4916], Fresh[4915], Fresh[4914], Fresh[4913], Fresh[4912], Fresh[4911], Fresh[4910]}), .outt ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, new_AGEMA_signal_2640, n2143}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2308 ( .ina ({new_AGEMA_signal_2204, new_AGEMA_signal_2203, new_AGEMA_signal_2202, n2139}), .inb ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, new_AGEMA_signal_1155, n2346}), .clk ( clk ), .rnd ({Fresh[4929], Fresh[4928], Fresh[4927], Fresh[4926], Fresh[4925], Fresh[4924], Fresh[4923], Fresh[4922], Fresh[4921], Fresh[4920]}), .outt ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, new_AGEMA_signal_2643, n2140}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2324 ( .ina ({new_AGEMA_signal_2216, new_AGEMA_signal_2215, new_AGEMA_signal_2214, n2157}), .inb ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2679}), .clk ( clk ), .rnd ({Fresh[4939], Fresh[4938], Fresh[4937], Fresh[4936], Fresh[4935], Fresh[4934], Fresh[4933], Fresh[4932], Fresh[4931], Fresh[4930]}), .outt ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, new_AGEMA_signal_2646, n2159}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2326 ( .ina ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, new_AGEMA_signal_2184, n2160}), .inb ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .clk ( clk ), .rnd ({Fresh[4949], Fresh[4948], Fresh[4947], Fresh[4946], Fresh[4945], Fresh[4944], Fresh[4943], Fresh[4942], Fresh[4941], Fresh[4940]}), .outt ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, new_AGEMA_signal_2649, n2161}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2330 ( .ina ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .inb ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, new_AGEMA_signal_1725, n2163}), .clk ( clk ), .rnd ({Fresh[4959], Fresh[4958], Fresh[4957], Fresh[4956], Fresh[4955], Fresh[4954], Fresh[4953], Fresh[4952], Fresh[4951], Fresh[4950]}), .outt ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, new_AGEMA_signal_2217, n2164}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2345 ( .ina ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, new_AGEMA_signal_1371, n2178}), .inb ({new_AGEMA_signal_2228, new_AGEMA_signal_2227, new_AGEMA_signal_2226, n2177}), .clk ( clk ), .rnd ({Fresh[4969], Fresh[4968], Fresh[4967], Fresh[4966], Fresh[4965], Fresh[4964], Fresh[4963], Fresh[4962], Fresh[4961], Fresh[4960]}), .outt ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, new_AGEMA_signal_2655, n2179}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2359 ( .ina ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .inb ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, new_AGEMA_signal_2235, n2191}), .clk ( clk ), .rnd ({Fresh[4979], Fresh[4978], Fresh[4977], Fresh[4976], Fresh[4975], Fresh[4974], Fresh[4973], Fresh[4972], Fresh[4971], Fresh[4970]}), .outt ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, new_AGEMA_signal_2658, n2192}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2370 ( .ina ({new_AGEMA_signal_2240, new_AGEMA_signal_2239, new_AGEMA_signal_2238, n2201}), .inb ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, new_AGEMA_signal_2661, n2200}), .clk ( clk ), .rnd ({Fresh[4989], Fresh[4988], Fresh[4987], Fresh[4986], Fresh[4985], Fresh[4984], Fresh[4983], Fresh[4982], Fresh[4981], Fresh[4980]}), .outt ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, new_AGEMA_signal_2955, n2203}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2382 ( .ina ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, new_AGEMA_signal_2244, n2217}), .inb ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, new_AGEMA_signal_1746, n2216}), .clk ( clk ), .rnd ({Fresh[4999], Fresh[4998], Fresh[4997], Fresh[4996], Fresh[4995], Fresh[4994], Fresh[4993], Fresh[4992], Fresh[4991], Fresh[4990]}), .outt ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, new_AGEMA_signal_2667, n2224}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2388 ( .ina ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, new_AGEMA_signal_2247, n2222}), .inb ({new_AGEMA_signal_2252, new_AGEMA_signal_2251, new_AGEMA_signal_2250, n2221}), .clk ( clk ), .rnd ({Fresh[5009], Fresh[5008], Fresh[5007], Fresh[5006], Fresh[5005], Fresh[5004], Fresh[5003], Fresh[5002], Fresh[5001], Fresh[5000]}), .outt ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, new_AGEMA_signal_2670, n2223}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2392 ( .ina ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, n2504}), .inb ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, new_AGEMA_signal_1755, n2226}), .clk ( clk ), .rnd ({Fresh[5019], Fresh[5018], Fresh[5017], Fresh[5016], Fresh[5015], Fresh[5014], Fresh[5013], Fresh[5012], Fresh[5011], Fresh[5010]}), .outt ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, new_AGEMA_signal_2253, n2229}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2399 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, new_AGEMA_signal_2676, n2233}), .clk ( clk ), .rnd ({Fresh[5029], Fresh[5028], Fresh[5027], Fresh[5026], Fresh[5025], Fresh[5024], Fresh[5023], Fresh[5022], Fresh[5021], Fresh[5020]}), .outt ({new_AGEMA_signal_2966, new_AGEMA_signal_2965, new_AGEMA_signal_2964, n2234}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2410 ( .ina ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, new_AGEMA_signal_2259, n2244}), .clk ( clk ), .rnd ({Fresh[5039], Fresh[5038], Fresh[5037], Fresh[5036], Fresh[5035], Fresh[5034], Fresh[5033], Fresh[5032], Fresh[5031], Fresh[5030]}), .outt ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, new_AGEMA_signal_2679, n2246}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2418 ( .ina ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2505}), .inb ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, new_AGEMA_signal_2265, n2253}), .clk ( clk ), .rnd ({Fresh[5049], Fresh[5048], Fresh[5047], Fresh[5046], Fresh[5045], Fresh[5044], Fresh[5043], Fresh[5042], Fresh[5041], Fresh[5040]}), .outt ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, new_AGEMA_signal_2682, n2254}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2425 ( .ina ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, new_AGEMA_signal_1779, n2540}), .inb ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, new_AGEMA_signal_2268, n2260}), .clk ( clk ), .rnd ({Fresh[5059], Fresh[5058], Fresh[5057], Fresh[5056], Fresh[5055], Fresh[5054], Fresh[5053], Fresh[5052], Fresh[5051], Fresh[5050]}), .outt ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, new_AGEMA_signal_2685, n2263}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2434 ( .ina ({new_AGEMA_signal_1394, new_AGEMA_signal_1393, new_AGEMA_signal_1392, n2266}), .inb ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, new_AGEMA_signal_1785, n2265}), .clk ( clk ), .rnd ({Fresh[5069], Fresh[5068], Fresh[5067], Fresh[5066], Fresh[5065], Fresh[5064], Fresh[5063], Fresh[5062], Fresh[5061], Fresh[5060]}), .outt ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, new_AGEMA_signal_2271, n2267}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2438 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_1790, new_AGEMA_signal_1789, new_AGEMA_signal_1788, n2269}), .clk ( clk ), .rnd ({Fresh[5079], Fresh[5078], Fresh[5077], Fresh[5076], Fresh[5075], Fresh[5074], Fresh[5073], Fresh[5072], Fresh[5071], Fresh[5070]}), .outt ({new_AGEMA_signal_2276, new_AGEMA_signal_2275, new_AGEMA_signal_2274, n2270}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2445 ( .ina ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, new_AGEMA_signal_1791, n2278}), .inb ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, new_AGEMA_signal_1794, n2277}), .clk ( clk ), .rnd ({Fresh[5089], Fresh[5088], Fresh[5087], Fresh[5086], Fresh[5085], Fresh[5084], Fresh[5083], Fresh[5082], Fresh[5081], Fresh[5080]}), .outt ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, new_AGEMA_signal_2277, n2279}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2450 ( .ina ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, new_AGEMA_signal_1017, n2779}), .inb ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, new_AGEMA_signal_1797, n2282}), .clk ( clk ), .rnd ({Fresh[5099], Fresh[5098], Fresh[5097], Fresh[5096], Fresh[5095], Fresh[5094], Fresh[5093], Fresh[5092], Fresh[5091], Fresh[5090]}), .outt ({new_AGEMA_signal_2282, new_AGEMA_signal_2281, new_AGEMA_signal_2280, n2283}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2453 ( .ina ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, new_AGEMA_signal_1668, n2773}), .inb ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, new_AGEMA_signal_2283, n2284}), .clk ( clk ), .rnd ({Fresh[5109], Fresh[5108], Fresh[5107], Fresh[5106], Fresh[5105], Fresh[5104], Fresh[5103], Fresh[5102], Fresh[5101], Fresh[5100]}), .outt ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, new_AGEMA_signal_2700, n2285}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2457 ( .ina ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .inb ({new_AGEMA_signal_2288, new_AGEMA_signal_2287, new_AGEMA_signal_2286, n2459}), .clk ( clk ), .rnd ({Fresh[5119], Fresh[5118], Fresh[5117], Fresh[5116], Fresh[5115], Fresh[5114], Fresh[5113], Fresh[5112], Fresh[5111], Fresh[5110]}), .outt ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, new_AGEMA_signal_2703, n2686}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2460 ( .ina ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, new_AGEMA_signal_2289, n2288}), .clk ( clk ), .rnd ({Fresh[5129], Fresh[5128], Fresh[5127], Fresh[5126], Fresh[5125], Fresh[5124], Fresh[5123], Fresh[5122], Fresh[5121], Fresh[5120]}), .outt ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, new_AGEMA_signal_2706, n2289}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2463 ( .ina ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, new_AGEMA_signal_2292, n2458}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[5139], Fresh[5138], Fresh[5137], Fresh[5136], Fresh[5135], Fresh[5134], Fresh[5133], Fresh[5132], Fresh[5131], Fresh[5130]}), .outt ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, new_AGEMA_signal_2709, n2297}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2465 ( .ina ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, new_AGEMA_signal_1125, n2624}), .inb ({new_AGEMA_signal_2192, new_AGEMA_signal_2191, new_AGEMA_signal_2190, n2291}), .clk ( clk ), .rnd ({Fresh[5149], Fresh[5148], Fresh[5147], Fresh[5146], Fresh[5145], Fresh[5144], Fresh[5143], Fresh[5142], Fresh[5141], Fresh[5140]}), .outt ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, new_AGEMA_signal_2712, n2292}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2473 ( .ina ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .inb ({new_AGEMA_signal_2300, new_AGEMA_signal_2299, new_AGEMA_signal_2298, n2300}), .clk ( clk ), .rnd ({Fresh[5159], Fresh[5158], Fresh[5157], Fresh[5156], Fresh[5155], Fresh[5154], Fresh[5153], Fresh[5152], Fresh[5151], Fresh[5150]}), .outt ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, new_AGEMA_signal_2715, n2301}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2483 ( .ina ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .inb ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, new_AGEMA_signal_2304, n2314}), .clk ( clk ), .rnd ({Fresh[5169], Fresh[5168], Fresh[5167], Fresh[5166], Fresh[5165], Fresh[5164], Fresh[5163], Fresh[5162], Fresh[5161], Fresh[5160]}), .outt ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, new_AGEMA_signal_2718, n2321}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2487 ( .ina ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, n2319}), .inb ({new_AGEMA_signal_1412, new_AGEMA_signal_1411, new_AGEMA_signal_1410, n2318}), .clk ( clk ), .rnd ({Fresh[5179], Fresh[5178], Fresh[5177], Fresh[5176], Fresh[5175], Fresh[5174], Fresh[5173], Fresh[5172], Fresh[5171], Fresh[5170]}), .outt ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, new_AGEMA_signal_1815, n2320}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2493 ( .ina ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, new_AGEMA_signal_1818, n2326}), .inb ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, new_AGEMA_signal_1821, n2325}), .clk ( clk ), .rnd ({Fresh[5189], Fresh[5188], Fresh[5187], Fresh[5186], Fresh[5185], Fresh[5184], Fresh[5183], Fresh[5182], Fresh[5181], Fresh[5180]}), .outt ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, new_AGEMA_signal_2307, n2334}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2497 ( .ina ({new_AGEMA_signal_2312, new_AGEMA_signal_2311, new_AGEMA_signal_2310, n2329}), .inb ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, new_AGEMA_signal_1017, n2779}), .clk ( clk ), .rnd ({Fresh[5199], Fresh[5198], Fresh[5197], Fresh[5196], Fresh[5195], Fresh[5194], Fresh[5193], Fresh[5192], Fresh[5191], Fresh[5190]}), .outt ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, new_AGEMA_signal_2721, n2332}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2498 ( .ina ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, n2677}), .inb ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, new_AGEMA_signal_2175, n2330}), .clk ( clk ), .rnd ({Fresh[5209], Fresh[5208], Fresh[5207], Fresh[5206], Fresh[5205], Fresh[5204], Fresh[5203], Fresh[5202], Fresh[5201], Fresh[5200]}), .outt ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, new_AGEMA_signal_2724, n2331}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2502 ( .ina ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, n2577}), .inb ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, new_AGEMA_signal_2727, n2335}), .clk ( clk ), .rnd ({Fresh[5219], Fresh[5218], Fresh[5217], Fresh[5216], Fresh[5215], Fresh[5214], Fresh[5213], Fresh[5212], Fresh[5211], Fresh[5210]}), .outt ({new_AGEMA_signal_2996, new_AGEMA_signal_2995, new_AGEMA_signal_2994, n2336}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2508 ( .ina ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, new_AGEMA_signal_2313, n2341}), .inb ({new_AGEMA_signal_1832, new_AGEMA_signal_1831, new_AGEMA_signal_1830, n2340}), .clk ( clk ), .rnd ({Fresh[5229], Fresh[5228], Fresh[5227], Fresh[5226], Fresh[5225], Fresh[5224], Fresh[5223], Fresh[5222], Fresh[5221], Fresh[5220]}), .outt ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, new_AGEMA_signal_2730, n2342}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2519 ( .ina ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, new_AGEMA_signal_1842, n2352}), .inb ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .clk ( clk ), .rnd ({Fresh[5239], Fresh[5238], Fresh[5237], Fresh[5236], Fresh[5235], Fresh[5234], Fresh[5233], Fresh[5232], Fresh[5231], Fresh[5230]}), .outt ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, new_AGEMA_signal_2316, n2367}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2523 ( .ina ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319, n2354}), .inb ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .clk ( clk ), .rnd ({Fresh[5249], Fresh[5248], Fresh[5247], Fresh[5246], Fresh[5245], Fresh[5244], Fresh[5243], Fresh[5242], Fresh[5241], Fresh[5240]}), .outt ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, new_AGEMA_signal_2733, n2358}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2547 ( .ina ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, new_AGEMA_signal_1857, n2385}), .inb ({new_AGEMA_signal_1862, new_AGEMA_signal_1861, new_AGEMA_signal_1860, n2384}), .clk ( clk ), .rnd ({Fresh[5259], Fresh[5258], Fresh[5257], Fresh[5256], Fresh[5255], Fresh[5254], Fresh[5253], Fresh[5252], Fresh[5251], Fresh[5250]}), .outt ({new_AGEMA_signal_2336, new_AGEMA_signal_2335, new_AGEMA_signal_2334, n2387}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2555 ( .ina ({new_AGEMA_signal_1868, new_AGEMA_signal_1867, new_AGEMA_signal_1866, n2391}), .inb ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, new_AGEMA_signal_2340, n2390}), .clk ( clk ), .rnd ({Fresh[5269], Fresh[5268], Fresh[5267], Fresh[5266], Fresh[5265], Fresh[5264], Fresh[5263], Fresh[5262], Fresh[5261], Fresh[5260]}), .outt ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, new_AGEMA_signal_2742, n2392}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2566 ( .ina ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, new_AGEMA_signal_1872, n2403}), .inb ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .clk ( clk ), .rnd ({Fresh[5279], Fresh[5278], Fresh[5277], Fresh[5276], Fresh[5275], Fresh[5274], Fresh[5273], Fresh[5272], Fresh[5271], Fresh[5270]}), .outt ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346, n2404}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2570 ( .ina ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, new_AGEMA_signal_1566, n2535}), .inb ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, new_AGEMA_signal_2349, n2408}), .clk ( clk ), .rnd ({Fresh[5289], Fresh[5288], Fresh[5287], Fresh[5286], Fresh[5285], Fresh[5284], Fresh[5283], Fresh[5282], Fresh[5281], Fresh[5280]}), .outt ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, new_AGEMA_signal_2748, n2409}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2575 ( .ina ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, new_AGEMA_signal_2352, n2574}), .inb ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, new_AGEMA_signal_1875, n2413}), .clk ( clk ), .rnd ({Fresh[5299], Fresh[5298], Fresh[5297], Fresh[5296], Fresh[5295], Fresh[5294], Fresh[5293], Fresh[5292], Fresh[5291], Fresh[5290]}), .outt ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, new_AGEMA_signal_2751, n2414}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2578 ( .ina ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2625}), .inb ({new_AGEMA_signal_1880, new_AGEMA_signal_1879, new_AGEMA_signal_1878, n2416}), .clk ( clk ), .rnd ({Fresh[5309], Fresh[5308], Fresh[5307], Fresh[5306], Fresh[5305], Fresh[5304], Fresh[5303], Fresh[5302], Fresh[5301], Fresh[5300]}), .outt ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, n2418}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2589 ( .ina ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, new_AGEMA_signal_2361, n2689}), .inb ({new_AGEMA_signal_1886, new_AGEMA_signal_1885, new_AGEMA_signal_1884, n2431}), .clk ( clk ), .rnd ({Fresh[5319], Fresh[5318], Fresh[5317], Fresh[5316], Fresh[5315], Fresh[5314], Fresh[5313], Fresh[5312], Fresh[5311], Fresh[5310]}), .outt ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, new_AGEMA_signal_2757, n2432}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2592 ( .ina ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, new_AGEMA_signal_1887, n2434}), .clk ( clk ), .rnd ({Fresh[5329], Fresh[5328], Fresh[5327], Fresh[5326], Fresh[5325], Fresh[5324], Fresh[5323], Fresh[5322], Fresh[5321], Fresh[5320]}), .outt ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, new_AGEMA_signal_2364, n2435}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2601 ( .ina ({new_AGEMA_signal_2372, new_AGEMA_signal_2371, new_AGEMA_signal_2370, n2445}), .inb ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2373, n2444}), .clk ( clk ), .rnd ({Fresh[5339], Fresh[5338], Fresh[5337], Fresh[5336], Fresh[5335], Fresh[5334], Fresh[5333], Fresh[5332], Fresh[5331], Fresh[5330]}), .outt ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, new_AGEMA_signal_2760, n2449}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2603 ( .ina ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .inb ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, new_AGEMA_signal_2376, n2447}), .clk ( clk ), .rnd ({Fresh[5349], Fresh[5348], Fresh[5347], Fresh[5346], Fresh[5345], Fresh[5344], Fresh[5343], Fresh[5342], Fresh[5341], Fresh[5340]}), .outt ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, new_AGEMA_signal_2763, n2448}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2609 ( .ina ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, new_AGEMA_signal_2379, n2454}), .inb ({new_AGEMA_signal_1442, new_AGEMA_signal_1441, new_AGEMA_signal_1440, n2453}), .clk ( clk ), .rnd ({Fresh[5359], Fresh[5358], Fresh[5357], Fresh[5356], Fresh[5355], Fresh[5354], Fresh[5353], Fresh[5352], Fresh[5351], Fresh[5350]}), .outt ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, new_AGEMA_signal_2766, n2455}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2612 ( .ina ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, n2687}), .inb ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, new_AGEMA_signal_2292, n2458}), .clk ( clk ), .rnd ({Fresh[5369], Fresh[5368], Fresh[5367], Fresh[5366], Fresh[5365], Fresh[5364], Fresh[5363], Fresh[5362], Fresh[5361], Fresh[5360]}), .outt ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, new_AGEMA_signal_2769, n2460}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2618 ( .ina ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, new_AGEMA_signal_1125, n2624}), .inb ({new_AGEMA_signal_1898, new_AGEMA_signal_1897, new_AGEMA_signal_1896, n2465}), .clk ( clk ), .rnd ({Fresh[5379], Fresh[5378], Fresh[5377], Fresh[5376], Fresh[5375], Fresh[5374], Fresh[5373], Fresh[5372], Fresh[5371], Fresh[5370]}), .outt ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, n2466}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2629 ( .ina ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, new_AGEMA_signal_1902, n2476}), .inb ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, new_AGEMA_signal_1455, n2475}), .clk ( clk ), .rnd ({Fresh[5389], Fresh[5388], Fresh[5387], Fresh[5386], Fresh[5385], Fresh[5384], Fresh[5383], Fresh[5382], Fresh[5381], Fresh[5380]}), .outt ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, new_AGEMA_signal_2385, n2477}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2634 ( .ina ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .inb ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, new_AGEMA_signal_2388, n2481}), .clk ( clk ), .rnd ({Fresh[5399], Fresh[5398], Fresh[5397], Fresh[5396], Fresh[5395], Fresh[5394], Fresh[5393], Fresh[5392], Fresh[5391], Fresh[5390]}), .outt ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, new_AGEMA_signal_2778, n2482}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2640 ( .ina ({new_AGEMA_signal_1910, new_AGEMA_signal_1909, new_AGEMA_signal_1908, n2487}), .inb ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, new_AGEMA_signal_1911, n2486}), .clk ( clk ), .rnd ({Fresh[5409], Fresh[5408], Fresh[5407], Fresh[5406], Fresh[5405], Fresh[5404], Fresh[5403], Fresh[5402], Fresh[5401], Fresh[5400]}), .outt ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, n2490}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2648 ( .ina ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, new_AGEMA_signal_1920, n2495}), .inb ({new_AGEMA_signal_2396, new_AGEMA_signal_2395, new_AGEMA_signal_2394, n2494}), .clk ( clk ), .rnd ({Fresh[5419], Fresh[5418], Fresh[5417], Fresh[5416], Fresh[5415], Fresh[5414], Fresh[5413], Fresh[5412], Fresh[5411], Fresh[5410]}), .outt ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, new_AGEMA_signal_2784, n2496}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2654 ( .ina ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, n2504}), .inb ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, new_AGEMA_signal_2787, n2503}), .clk ( clk ), .rnd ({Fresh[5429], Fresh[5428], Fresh[5427], Fresh[5426], Fresh[5425], Fresh[5424], Fresh[5423], Fresh[5422], Fresh[5421], Fresh[5420]}), .outt ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, new_AGEMA_signal_3045, n2507}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2664 ( .ina ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, new_AGEMA_signal_2400, n2518}), .inb ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, new_AGEMA_signal_2790, n2517}), .clk ( clk ), .rnd ({Fresh[5439], Fresh[5438], Fresh[5437], Fresh[5436], Fresh[5435], Fresh[5434], Fresh[5433], Fresh[5432], Fresh[5431], Fresh[5430]}), .outt ({new_AGEMA_signal_3050, new_AGEMA_signal_3049, new_AGEMA_signal_3048, n2525}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2669 ( .ina ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, new_AGEMA_signal_2403, n2523}), .inb ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, new_AGEMA_signal_2406, n2522}), .clk ( clk ), .rnd ({Fresh[5449], Fresh[5448], Fresh[5447], Fresh[5446], Fresh[5445], Fresh[5444], Fresh[5443], Fresh[5442], Fresh[5441], Fresh[5440]}), .outt ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, new_AGEMA_signal_2793, n2524}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2676 ( .ina ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2409, n2532}), .inb ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .clk ( clk ), .rnd ({Fresh[5459], Fresh[5458], Fresh[5457], Fresh[5456], Fresh[5455], Fresh[5454], Fresh[5453], Fresh[5452], Fresh[5451], Fresh[5450]}), .outt ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, new_AGEMA_signal_2796, n2537}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2678 ( .ina ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, new_AGEMA_signal_1566, n2535}), .inb ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, new_AGEMA_signal_2412, n2534}), .clk ( clk ), .rnd ({Fresh[5469], Fresh[5468], Fresh[5467], Fresh[5466], Fresh[5465], Fresh[5464], Fresh[5463], Fresh[5462], Fresh[5461], Fresh[5460]}), .outt ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, new_AGEMA_signal_2799, n2536}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2684 ( .ina ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}), .inb ({new_AGEMA_signal_1934, new_AGEMA_signal_1933, new_AGEMA_signal_1932, n2546}), .clk ( clk ), .rnd ({Fresh[5479], Fresh[5478], Fresh[5477], Fresh[5476], Fresh[5475], Fresh[5474], Fresh[5473], Fresh[5472], Fresh[5471], Fresh[5470]}), .outt ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, new_AGEMA_signal_2418, n2547}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2693 ( .ina ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .inb ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, n2556}), .clk ( clk ), .rnd ({Fresh[5489], Fresh[5488], Fresh[5487], Fresh[5486], Fresh[5485], Fresh[5484], Fresh[5483], Fresh[5482], Fresh[5481], Fresh[5480]}), .outt ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, new_AGEMA_signal_2802, n2557}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2699 ( .ina ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2433, n2715}), .inb ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, new_AGEMA_signal_1941, n2564}), .clk ( clk ), .rnd ({Fresh[5499], Fresh[5498], Fresh[5497], Fresh[5496], Fresh[5495], Fresh[5494], Fresh[5493], Fresh[5492], Fresh[5491], Fresh[5490]}), .outt ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, new_AGEMA_signal_2805, n2565}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2704 ( .ina ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, new_AGEMA_signal_2352, n2574}), .inb ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, new_AGEMA_signal_2436, n2573}), .clk ( clk ), .rnd ({Fresh[5509], Fresh[5508], Fresh[5507], Fresh[5506], Fresh[5505], Fresh[5504], Fresh[5503], Fresh[5502], Fresh[5501], Fresh[5500]}), .outt ({new_AGEMA_signal_2810, new_AGEMA_signal_2809, new_AGEMA_signal_2808, n2591}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2709 ( .ina ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, new_AGEMA_signal_2442, n2579}), .inb ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, new_AGEMA_signal_1947, n2578}), .clk ( clk ), .rnd ({Fresh[5519], Fresh[5518], Fresh[5517], Fresh[5516], Fresh[5515], Fresh[5514], Fresh[5513], Fresh[5512], Fresh[5511], Fresh[5510]}), .outt ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, new_AGEMA_signal_2811, n2580}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2727 ( .ina ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, new_AGEMA_signal_1470, n2601}), .inb ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2600}), .clk ( clk ), .rnd ({Fresh[5529], Fresh[5528], Fresh[5527], Fresh[5526], Fresh[5525], Fresh[5524], Fresh[5523], Fresh[5522], Fresh[5521], Fresh[5520]}), .outt ({new_AGEMA_signal_1964, new_AGEMA_signal_1963, new_AGEMA_signal_1962, n2602}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2738 ( .ina ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, new_AGEMA_signal_2460, n2618}), .inb ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, new_AGEMA_signal_1473, n2617}), .clk ( clk ), .rnd ({Fresh[5539], Fresh[5538], Fresh[5537], Fresh[5536], Fresh[5535], Fresh[5534], Fresh[5533], Fresh[5532], Fresh[5531], Fresh[5530]}), .outt ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, new_AGEMA_signal_2817, n2619}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2744 ( .ina ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .inb ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, new_AGEMA_signal_2463, n2626}), .clk ( clk ), .rnd ({Fresh[5549], Fresh[5548], Fresh[5547], Fresh[5546], Fresh[5545], Fresh[5544], Fresh[5543], Fresh[5542], Fresh[5541], Fresh[5540]}), .outt ({new_AGEMA_signal_2822, new_AGEMA_signal_2821, new_AGEMA_signal_2820, n2628}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2753 ( .ina ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, new_AGEMA_signal_2466, n2644}), .inb ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .clk ( clk ), .rnd ({Fresh[5559], Fresh[5558], Fresh[5557], Fresh[5556], Fresh[5555], Fresh[5554], Fresh[5553], Fresh[5552], Fresh[5551], Fresh[5550]}), .outt ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, new_AGEMA_signal_2823, n2649}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2755 ( .ina ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, n2647}), .inb ({new_AGEMA_signal_1982, new_AGEMA_signal_1981, new_AGEMA_signal_1980, n2646}), .clk ( clk ), .rnd ({Fresh[5569], Fresh[5568], Fresh[5567], Fresh[5566], Fresh[5565], Fresh[5564], Fresh[5563], Fresh[5562], Fresh[5561], Fresh[5560]}), .outt ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, new_AGEMA_signal_2469, n2648}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2765 ( .ina ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, new_AGEMA_signal_2475, n2663}), .clk ( clk ), .rnd ({Fresh[5579], Fresh[5578], Fresh[5577], Fresh[5576], Fresh[5575], Fresh[5574], Fresh[5573], Fresh[5572], Fresh[5571], Fresh[5570]}), .outt ({new_AGEMA_signal_2828, new_AGEMA_signal_2827, new_AGEMA_signal_2826, n2664}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2771 ( .ina ({new_AGEMA_signal_1988, new_AGEMA_signal_1987, new_AGEMA_signal_1986, n2675}), .inb ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, n2674}), .clk ( clk ), .rnd ({Fresh[5589], Fresh[5588], Fresh[5587], Fresh[5586], Fresh[5585], Fresh[5584], Fresh[5583], Fresh[5582], Fresh[5581], Fresh[5580]}), .outt ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, new_AGEMA_signal_2829, n2681}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2773 ( .ina ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2679}), .inb ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, new_AGEMA_signal_1989, n2678}), .clk ( clk ), .rnd ({Fresh[5599], Fresh[5598], Fresh[5597], Fresh[5596], Fresh[5595], Fresh[5594], Fresh[5593], Fresh[5592], Fresh[5591], Fresh[5590]}), .outt ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, new_AGEMA_signal_2478, n2680}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2776 ( .ina ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, new_AGEMA_signal_2091, n2684}), .inb ({new_AGEMA_signal_1184, new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2683}), .clk ( clk ), .rnd ({Fresh[5609], Fresh[5608], Fresh[5607], Fresh[5606], Fresh[5605], Fresh[5604], Fresh[5603], Fresh[5602], Fresh[5601], Fresh[5600]}), .outt ({new_AGEMA_signal_2834, new_AGEMA_signal_2833, new_AGEMA_signal_2832, n2685}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2778 ( .ina ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, n2687}), .inb ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}), .clk ( clk ), .rnd ({Fresh[5619], Fresh[5618], Fresh[5617], Fresh[5616], Fresh[5615], Fresh[5614], Fresh[5613], Fresh[5612], Fresh[5611], Fresh[5610]}), .outt ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, new_AGEMA_signal_2835, n2698}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2779 ( .ina ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, new_AGEMA_signal_2361, n2689}), .inb ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .clk ( clk ), .rnd ({Fresh[5629], Fresh[5628], Fresh[5627], Fresh[5626], Fresh[5625], Fresh[5624], Fresh[5623], Fresh[5622], Fresh[5621], Fresh[5620]}), .outt ({new_AGEMA_signal_2840, new_AGEMA_signal_2839, new_AGEMA_signal_2838, n2692}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2793 ( .ina ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2433, n2715}), .inb ({new_AGEMA_signal_1484, new_AGEMA_signal_1483, new_AGEMA_signal_1482, n2714}), .clk ( clk ), .rnd ({Fresh[5639], Fresh[5638], Fresh[5637], Fresh[5636], Fresh[5635], Fresh[5634], Fresh[5633], Fresh[5632], Fresh[5631], Fresh[5630]}), .outt ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, new_AGEMA_signal_2841, n2716}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2800 ( .ina ({new_AGEMA_signal_2006, new_AGEMA_signal_2005, new_AGEMA_signal_2004, n2727}), .inb ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, new_AGEMA_signal_2007, n2726}), .clk ( clk ), .rnd ({Fresh[5649], Fresh[5648], Fresh[5647], Fresh[5646], Fresh[5645], Fresh[5644], Fresh[5643], Fresh[5642], Fresh[5641], Fresh[5640]}), .outt ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, new_AGEMA_signal_2487, n2728}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2804 ( .ina ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, n2734}), .inb ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, new_AGEMA_signal_2490, n2733}), .clk ( clk ), .rnd ({Fresh[5659], Fresh[5658], Fresh[5657], Fresh[5656], Fresh[5655], Fresh[5654], Fresh[5653], Fresh[5652], Fresh[5651], Fresh[5650]}), .outt ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, new_AGEMA_signal_2847, n2735}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2808 ( .ina ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, new_AGEMA_signal_1575, n2741}), .inb ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, new_AGEMA_signal_2493, n2740}), .clk ( clk ), .rnd ({Fresh[5669], Fresh[5668], Fresh[5667], Fresh[5666], Fresh[5665], Fresh[5664], Fresh[5663], Fresh[5662], Fresh[5661], Fresh[5660]}), .outt ({new_AGEMA_signal_2852, new_AGEMA_signal_2851, new_AGEMA_signal_2850, n2743}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2813 ( .ina ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .inb ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, new_AGEMA_signal_2013, n2749}), .clk ( clk ), .rnd ({Fresh[5679], Fresh[5678], Fresh[5677], Fresh[5676], Fresh[5675], Fresh[5674], Fresh[5673], Fresh[5672], Fresh[5671], Fresh[5670]}), .outt ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, new_AGEMA_signal_2496, n2751}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2817 ( .ina ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, new_AGEMA_signal_2499, n2757}), .inb ({new_AGEMA_signal_2018, new_AGEMA_signal_2017, new_AGEMA_signal_2016, n2756}), .clk ( clk ), .rnd ({Fresh[5689], Fresh[5688], Fresh[5687], Fresh[5686], Fresh[5685], Fresh[5684], Fresh[5683], Fresh[5682], Fresh[5681], Fresh[5680]}), .outt ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, new_AGEMA_signal_2853, n2758}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2820 ( .ina ({new_AGEMA_signal_1520, new_AGEMA_signal_1519, new_AGEMA_signal_1518, n2763}), .inb ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, new_AGEMA_signal_2502, n2762}), .clk ( clk ), .rnd ({Fresh[5699], Fresh[5698], Fresh[5697], Fresh[5696], Fresh[5695], Fresh[5694], Fresh[5693], Fresh[5692], Fresh[5691], Fresh[5690]}), .outt ({new_AGEMA_signal_2858, new_AGEMA_signal_2857, new_AGEMA_signal_2856, n2764}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2827 ( .ina ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, new_AGEMA_signal_2508, n2776}), .inb ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, new_AGEMA_signal_2511, n2775}), .clk ( clk ), .rnd ({Fresh[5709], Fresh[5708], Fresh[5707], Fresh[5706], Fresh[5705], Fresh[5704], Fresh[5703], Fresh[5702], Fresh[5701], Fresh[5700]}), .outt ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, new_AGEMA_signal_2859, n2800}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2831 ( .ina ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, new_AGEMA_signal_1977, n2784}), .inb ({new_AGEMA_signal_2024, new_AGEMA_signal_2023, new_AGEMA_signal_2022, n2783}), .clk ( clk ), .rnd ({Fresh[5719], Fresh[5718], Fresh[5717], Fresh[5716], Fresh[5715], Fresh[5714], Fresh[5713], Fresh[5712], Fresh[5711], Fresh[5710]}), .outt ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, new_AGEMA_signal_2514, n2788}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2837 ( .ina ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .inb ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, new_AGEMA_signal_2517, n2795}), .clk ( clk ), .rnd ({Fresh[5729], Fresh[5728], Fresh[5727], Fresh[5726], Fresh[5725], Fresh[5724], Fresh[5723], Fresh[5722], Fresh[5721], Fresh[5720]}), .outt ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, new_AGEMA_signal_2865, n2797}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2846 ( .ina ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, new_AGEMA_signal_2520, n2814}), .inb ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .rnd ({Fresh[5739], Fresh[5738], Fresh[5737], Fresh[5736], Fresh[5735], Fresh[5734], Fresh[5733], Fresh[5732], Fresh[5731], Fresh[5730]}), .outt ({new_AGEMA_signal_2870, new_AGEMA_signal_2869, new_AGEMA_signal_2868, n2822}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2849 ( .ina ({new_AGEMA_signal_1496, new_AGEMA_signal_1495, new_AGEMA_signal_1494, n2820}), .inb ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, new_AGEMA_signal_2037, n2819}), .clk ( clk ), .rnd ({Fresh[5749], Fresh[5748], Fresh[5747], Fresh[5746], Fresh[5745], Fresh[5744], Fresh[5743], Fresh[5742], Fresh[5741], Fresh[5740]}), .outt ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, new_AGEMA_signal_2523, n2821}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1983 ( .ina ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .inb ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, new_AGEMA_signal_2529, n1928}), .clk ( clk ), .rnd ({Fresh[5759], Fresh[5758], Fresh[5757], Fresh[5756], Fresh[5755], Fresh[5754], Fresh[5753], Fresh[5752], Fresh[5751], Fresh[5750]}), .outt ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, new_AGEMA_signal_2871, n1934}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U1998 ( .ina ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, new_AGEMA_signal_2532, n1931}), .inb ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, new_AGEMA_signal_1224, n1930}), .clk ( clk ), .rnd ({Fresh[5769], Fresh[5768], Fresh[5767], Fresh[5766], Fresh[5765], Fresh[5764], Fresh[5763], Fresh[5762], Fresh[5761], Fresh[5760]}), .outt ({new_AGEMA_signal_2876, new_AGEMA_signal_2875, new_AGEMA_signal_2874, n1932}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2015 ( .ina ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, new_AGEMA_signal_2535, n1939}), .inb ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}), .clk ( clk ), .rnd ({Fresh[5779], Fresh[5778], Fresh[5777], Fresh[5776], Fresh[5775], Fresh[5774], Fresh[5773], Fresh[5772], Fresh[5771], Fresh[5770]}), .outt ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, new_AGEMA_signal_2877, n1940}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2033 ( .ina ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, new_AGEMA_signal_2538, n1948}), .inb ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, new_AGEMA_signal_2541, n1947}), .clk ( clk ), .rnd ({Fresh[5789], Fresh[5788], Fresh[5787], Fresh[5786], Fresh[5785], Fresh[5784], Fresh[5783], Fresh[5782], Fresh[5781], Fresh[5780]}), .outt ({new_AGEMA_signal_2882, new_AGEMA_signal_2881, new_AGEMA_signal_2880, n1961}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2050 ( .ina ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, new_AGEMA_signal_2544, n1954}), .inb ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, new_AGEMA_signal_2547, n1953}), .clk ( clk ), .rnd ({Fresh[5799], Fresh[5798], Fresh[5797], Fresh[5796], Fresh[5795], Fresh[5794], Fresh[5793], Fresh[5792], Fresh[5791], Fresh[5790]}), .outt ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, new_AGEMA_signal_2883, n1955}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2066 ( .ina ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, new_AGEMA_signal_2079, n1966}), .inb ({new_AGEMA_signal_2084, new_AGEMA_signal_2083, new_AGEMA_signal_2082, n1965}), .clk ( clk ), .rnd ({Fresh[5809], Fresh[5808], Fresh[5807], Fresh[5806], Fresh[5805], Fresh[5804], Fresh[5803], Fresh[5802], Fresh[5801], Fresh[5800]}), .outt ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, new_AGEMA_signal_2553, n1967}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2085 ( .ina ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, new_AGEMA_signal_2889, n1970}), .inb ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, new_AGEMA_signal_2559, n1969}), .clk ( clk ), .rnd ({Fresh[5819], Fresh[5818], Fresh[5817], Fresh[5816], Fresh[5815], Fresh[5814], Fresh[5813], Fresh[5812], Fresh[5811], Fresh[5810]}), .outt ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, new_AGEMA_signal_3123, n1984}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2103 ( .ina ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, new_AGEMA_signal_1296, n1976}), .inb ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, new_AGEMA_signal_2565, n1975}), .clk ( clk ), .rnd ({Fresh[5829], Fresh[5828], Fresh[5827], Fresh[5826], Fresh[5825], Fresh[5824], Fresh[5823], Fresh[5822], Fresh[5821], Fresh[5820]}), .outt ({new_AGEMA_signal_2894, new_AGEMA_signal_2893, new_AGEMA_signal_2892, n1977}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2108 ( .ina ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .inb ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, new_AGEMA_signal_2568, n1980}), .clk ( clk ), .rnd ({Fresh[5839], Fresh[5838], Fresh[5837], Fresh[5836], Fresh[5835], Fresh[5834], Fresh[5833], Fresh[5832], Fresh[5831], Fresh[5830]}), .outt ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, new_AGEMA_signal_2895, n1981}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2115 ( .ina ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .inb ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, new_AGEMA_signal_2103, n1986}), .clk ( clk ), .rnd ({Fresh[5849], Fresh[5848], Fresh[5847], Fresh[5846], Fresh[5845], Fresh[5844], Fresh[5843], Fresh[5842], Fresh[5841], Fresh[5840]}), .outt ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, new_AGEMA_signal_2571, n1987}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2127 ( .ina ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, new_AGEMA_signal_2574, n1997}), .inb ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, new_AGEMA_signal_2109, n1996}), .clk ( clk ), .rnd ({Fresh[5859], Fresh[5858], Fresh[5857], Fresh[5856], Fresh[5855], Fresh[5854], Fresh[5853], Fresh[5852], Fresh[5851], Fresh[5850]}), .outt ({new_AGEMA_signal_2900, new_AGEMA_signal_2899, new_AGEMA_signal_2898, n1998}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2146 ( .ina ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, new_AGEMA_signal_1593, n2008}), .inb ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, new_AGEMA_signal_2580, n2007}), .clk ( clk ), .rnd ({Fresh[5869], Fresh[5868], Fresh[5867], Fresh[5866], Fresh[5865], Fresh[5864], Fresh[5863], Fresh[5862], Fresh[5861], Fresh[5860]}), .outt ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, new_AGEMA_signal_2901, n2010}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2162 ( .ina ({new_AGEMA_signal_1610, new_AGEMA_signal_1609, new_AGEMA_signal_1608, n2022}), .inb ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, new_AGEMA_signal_2124, n2021}), .clk ( clk ), .rnd ({Fresh[5879], Fresh[5878], Fresh[5877], Fresh[5876], Fresh[5875], Fresh[5874], Fresh[5873], Fresh[5872], Fresh[5871], Fresh[5870]}), .outt ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, new_AGEMA_signal_2583, n2024}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2177 ( .ina ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, new_AGEMA_signal_2127, n2033}), .inb ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, new_AGEMA_signal_2586, n2032}), .clk ( clk ), .rnd ({Fresh[5889], Fresh[5888], Fresh[5887], Fresh[5886], Fresh[5885], Fresh[5884], Fresh[5883], Fresh[5882], Fresh[5881], Fresh[5880]}), .outt ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, new_AGEMA_signal_2907, n2035}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2186 ( .ina ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, new_AGEMA_signal_2589, n2041}), .inb ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}), .clk ( clk ), .rnd ({Fresh[5899], Fresh[5898], Fresh[5897], Fresh[5896], Fresh[5895], Fresh[5894], Fresh[5893], Fresh[5892], Fresh[5891], Fresh[5890]}), .outt ({new_AGEMA_signal_2912, new_AGEMA_signal_2911, new_AGEMA_signal_2910, n2054}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2190 ( .ina ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .inb ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, new_AGEMA_signal_2592, n2043}), .clk ( clk ), .rnd ({Fresh[5909], Fresh[5908], Fresh[5907], Fresh[5906], Fresh[5905], Fresh[5904], Fresh[5903], Fresh[5902], Fresh[5901], Fresh[5900]}), .outt ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, new_AGEMA_signal_2913, n2048}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2195 ( .ina ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, new_AGEMA_signal_2595, n2046}), .inb ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .rnd ({Fresh[5919], Fresh[5918], Fresh[5917], Fresh[5916], Fresh[5915], Fresh[5914], Fresh[5913], Fresh[5912], Fresh[5911], Fresh[5910]}), .outt ({new_AGEMA_signal_2918, new_AGEMA_signal_2917, new_AGEMA_signal_2916, n2047}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2206 ( .ina ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, new_AGEMA_signal_2598, n2058}), .inb ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, new_AGEMA_signal_1647, n2057}), .clk ( clk ), .rnd ({Fresh[5929], Fresh[5928], Fresh[5927], Fresh[5926], Fresh[5925], Fresh[5924], Fresh[5923], Fresh[5922], Fresh[5921], Fresh[5920]}), .outt ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, new_AGEMA_signal_2919, n2059}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2213 ( .ina ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, new_AGEMA_signal_2601, n2063}), .inb ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, new_AGEMA_signal_1653, n2062}), .clk ( clk ), .rnd ({Fresh[5939], Fresh[5938], Fresh[5937], Fresh[5936], Fresh[5935], Fresh[5934], Fresh[5933], Fresh[5932], Fresh[5931], Fresh[5930]}), .outt ({new_AGEMA_signal_2924, new_AGEMA_signal_2923, new_AGEMA_signal_2922, n2064}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2229 ( .ina ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, new_AGEMA_signal_2607, n2076}), .inb ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, new_AGEMA_signal_1341, n2075}), .clk ( clk ), .rnd ({Fresh[5949], Fresh[5948], Fresh[5947], Fresh[5946], Fresh[5945], Fresh[5944], Fresh[5943], Fresh[5942], Fresh[5941], Fresh[5940]}), .outt ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, new_AGEMA_signal_2925, n2077}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2249 ( .ina ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, new_AGEMA_signal_2619, n2090}), .inb ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, new_AGEMA_signal_2172, n2089}), .clk ( clk ), .rnd ({Fresh[5959], Fresh[5958], Fresh[5957], Fresh[5956], Fresh[5955], Fresh[5954], Fresh[5953], Fresh[5952], Fresh[5951], Fresh[5950]}), .outt ({new_AGEMA_signal_2930, new_AGEMA_signal_2929, new_AGEMA_signal_2928, n2158}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2255 ( .ina ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, new_AGEMA_signal_2622, n2093}), .inb ({new_AGEMA_signal_2180, new_AGEMA_signal_2179, new_AGEMA_signal_2178, n2092}), .clk ( clk ), .rnd ({Fresh[5969], Fresh[5968], Fresh[5967], Fresh[5966], Fresh[5965], Fresh[5964], Fresh[5963], Fresh[5962], Fresh[5961], Fresh[5960]}), .outt ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, new_AGEMA_signal_2931, n2095}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2274 ( .ina ({new_AGEMA_signal_2936, new_AGEMA_signal_2935, new_AGEMA_signal_2934, n2116}), .inb ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, new_AGEMA_signal_1686, n2115}), .clk ( clk ), .rnd ({Fresh[5979], Fresh[5978], Fresh[5977], Fresh[5976], Fresh[5975], Fresh[5974], Fresh[5973], Fresh[5972], Fresh[5971], Fresh[5970]}), .outt ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, new_AGEMA_signal_3159, n2117}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2283 ( .ina ({new_AGEMA_signal_1691, new_AGEMA_signal_1690, new_AGEMA_signal_1689, n2121}), .inb ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, new_AGEMA_signal_2631, n2120}), .clk ( clk ), .rnd ({Fresh[5989], Fresh[5988], Fresh[5987], Fresh[5986], Fresh[5985], Fresh[5984], Fresh[5983], Fresh[5982], Fresh[5981], Fresh[5980]}), .outt ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, new_AGEMA_signal_2937, n2123}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2300 ( .ina ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, n2687}), .inb ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, new_AGEMA_signal_2196, n2134}), .clk ( clk ), .rnd ({Fresh[5999], Fresh[5998], Fresh[5997], Fresh[5996], Fresh[5995], Fresh[5994], Fresh[5993], Fresh[5992], Fresh[5991], Fresh[5990]}), .outt ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, new_AGEMA_signal_2637, n2135}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2309 ( .ina ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .inb ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, new_AGEMA_signal_2643, n2140}), .clk ( clk ), .rnd ({Fresh[6009], Fresh[6008], Fresh[6007], Fresh[6006], Fresh[6005], Fresh[6004], Fresh[6003], Fresh[6002], Fresh[6001], Fresh[6000]}), .outt ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, new_AGEMA_signal_2943, n2141}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2327 ( .ina ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}), .inb ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, new_AGEMA_signal_2649, n2161}), .clk ( clk ), .rnd ({Fresh[6019], Fresh[6018], Fresh[6017], Fresh[6016], Fresh[6015], Fresh[6014], Fresh[6013], Fresh[6012], Fresh[6011], Fresh[6010]}), .outt ({new_AGEMA_signal_2948, new_AGEMA_signal_2947, new_AGEMA_signal_2946, n2166}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2331 ( .ina ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .inb ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, new_AGEMA_signal_2217, n2164}), .clk ( clk ), .rnd ({Fresh[6029], Fresh[6028], Fresh[6027], Fresh[6026], Fresh[6025], Fresh[6024], Fresh[6023], Fresh[6022], Fresh[6021], Fresh[6020]}), .outt ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, new_AGEMA_signal_2652, n2165}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2346 ( .ina ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, new_AGEMA_signal_2655, n2179}), .inb ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .clk ( clk ), .rnd ({Fresh[6039], Fresh[6038], Fresh[6037], Fresh[6036], Fresh[6035], Fresh[6034], Fresh[6033], Fresh[6032], Fresh[6031], Fresh[6030]}), .outt ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, new_AGEMA_signal_2949, n2180}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2360 ( .ina ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, new_AGEMA_signal_2232, n2193}), .inb ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, new_AGEMA_signal_2658, n2192}), .clk ( clk ), .rnd ({Fresh[6049], Fresh[6048], Fresh[6047], Fresh[6046], Fresh[6045], Fresh[6044], Fresh[6043], Fresh[6042], Fresh[6041], Fresh[6040]}), .outt ({new_AGEMA_signal_2954, new_AGEMA_signal_2953, new_AGEMA_signal_2952, n2194}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2372 ( .ina ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, new_AGEMA_signal_2955, n2203}), .inb ({new_AGEMA_signal_2666, new_AGEMA_signal_2665, new_AGEMA_signal_2664, n2202}), .clk ( clk ), .rnd ({Fresh[6059], Fresh[6058], Fresh[6057], Fresh[6056], Fresh[6055], Fresh[6054], Fresh[6053], Fresh[6052], Fresh[6051], Fresh[6050]}), .outt ({new_AGEMA_signal_3182, new_AGEMA_signal_3181, new_AGEMA_signal_3180, n2204}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2389 ( .ina ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, new_AGEMA_signal_2667, n2224}), .inb ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, new_AGEMA_signal_2670, n2223}), .clk ( clk ), .rnd ({Fresh[6069], Fresh[6068], Fresh[6067], Fresh[6066], Fresh[6065], Fresh[6064], Fresh[6063], Fresh[6062], Fresh[6061], Fresh[6060]}), .outt ({new_AGEMA_signal_2960, new_AGEMA_signal_2959, new_AGEMA_signal_2958, n2225}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2394 ( .ina ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, new_AGEMA_signal_2253, n2229}), .inb ({new_AGEMA_signal_1760, new_AGEMA_signal_1759, new_AGEMA_signal_1758, n2228}), .clk ( clk ), .rnd ({Fresh[6079], Fresh[6078], Fresh[6077], Fresh[6076], Fresh[6075], Fresh[6074], Fresh[6073], Fresh[6072], Fresh[6071], Fresh[6070]}), .outt ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, new_AGEMA_signal_2673, n2230}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2400 ( .ina ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, new_AGEMA_signal_2061, n2235}), .inb ({new_AGEMA_signal_2966, new_AGEMA_signal_2965, new_AGEMA_signal_2964, n2234}), .clk ( clk ), .rnd ({Fresh[6089], Fresh[6088], Fresh[6087], Fresh[6086], Fresh[6085], Fresh[6084], Fresh[6083], Fresh[6082], Fresh[6081], Fresh[6080]}), .outt ({new_AGEMA_signal_3188, new_AGEMA_signal_3187, new_AGEMA_signal_3186, n2236}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2412 ( .ina ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, new_AGEMA_signal_2679, n2246}), .inb ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, new_AGEMA_signal_1776, n2245}), .clk ( clk ), .rnd ({Fresh[6099], Fresh[6098], Fresh[6097], Fresh[6096], Fresh[6095], Fresh[6094], Fresh[6093], Fresh[6092], Fresh[6091], Fresh[6090]}), .outt ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, new_AGEMA_signal_2967, n2247}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2419 ( .ina ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, new_AGEMA_signal_2682, n2254}), .inb ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, n2785}), .clk ( clk ), .rnd ({Fresh[6109], Fresh[6108], Fresh[6107], Fresh[6106], Fresh[6105], Fresh[6104], Fresh[6103], Fresh[6102], Fresh[6101], Fresh[6100]}), .outt ({new_AGEMA_signal_2972, new_AGEMA_signal_2971, new_AGEMA_signal_2970, n2255}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2427 ( .ina ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, new_AGEMA_signal_2685, n2263}), .inb ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, new_AGEMA_signal_1389, n2262}), .clk ( clk ), .rnd ({Fresh[6119], Fresh[6118], Fresh[6117], Fresh[6116], Fresh[6115], Fresh[6114], Fresh[6113], Fresh[6112], Fresh[6111], Fresh[6110]}), .outt ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, new_AGEMA_signal_2973, n2264}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2435 ( .ina ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, new_AGEMA_signal_2691, n2752}), .inb ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, new_AGEMA_signal_2271, n2267}), .clk ( clk ), .rnd ({Fresh[6129], Fresh[6128], Fresh[6127], Fresh[6126], Fresh[6125], Fresh[6124], Fresh[6123], Fresh[6122], Fresh[6121], Fresh[6120]}), .outt ({new_AGEMA_signal_2978, new_AGEMA_signal_2977, new_AGEMA_signal_2976, n2271}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2446 ( .ina ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .inb ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, new_AGEMA_signal_2277, n2279}), .clk ( clk ), .rnd ({Fresh[6139], Fresh[6138], Fresh[6137], Fresh[6136], Fresh[6135], Fresh[6134], Fresh[6133], Fresh[6132], Fresh[6131], Fresh[6130]}), .outt ({new_AGEMA_signal_2696, new_AGEMA_signal_2695, new_AGEMA_signal_2694, n2280}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2451 ( .ina ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({new_AGEMA_signal_2282, new_AGEMA_signal_2281, new_AGEMA_signal_2280, n2283}), .clk ( clk ), .rnd ({Fresh[6149], Fresh[6148], Fresh[6147], Fresh[6146], Fresh[6145], Fresh[6144], Fresh[6143], Fresh[6142], Fresh[6141], Fresh[6140]}), .outt ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, new_AGEMA_signal_2697, n2286}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2461 ( .ina ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, new_AGEMA_signal_2703, n2686}), .inb ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, new_AGEMA_signal_2706, n2289}), .clk ( clk ), .rnd ({Fresh[6159], Fresh[6158], Fresh[6157], Fresh[6156], Fresh[6155], Fresh[6154], Fresh[6153], Fresh[6152], Fresh[6151], Fresh[6150]}), .outt ({new_AGEMA_signal_2984, new_AGEMA_signal_2983, new_AGEMA_signal_2982, n2304}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2466 ( .ina ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, new_AGEMA_signal_2295, n2293}), .inb ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, new_AGEMA_signal_2712, n2292}), .clk ( clk ), .rnd ({Fresh[6169], Fresh[6168], Fresh[6167], Fresh[6166], Fresh[6165], Fresh[6164], Fresh[6163], Fresh[6162], Fresh[6161], Fresh[6160]}), .outt ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, new_AGEMA_signal_2985, n2295}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2488 ( .ina ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, new_AGEMA_signal_2718, n2321}), .inb ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, new_AGEMA_signal_1815, n2320}), .clk ( clk ), .rnd ({Fresh[6179], Fresh[6178], Fresh[6177], Fresh[6176], Fresh[6175], Fresh[6174], Fresh[6173], Fresh[6172], Fresh[6171], Fresh[6170]}), .outt ({new_AGEMA_signal_2990, new_AGEMA_signal_2989, new_AGEMA_signal_2988, n2322}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2499 ( .ina ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, new_AGEMA_signal_2721, n2332}), .inb ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, new_AGEMA_signal_2724, n2331}), .clk ( clk ), .rnd ({Fresh[6189], Fresh[6188], Fresh[6187], Fresh[6186], Fresh[6185], Fresh[6184], Fresh[6183], Fresh[6182], Fresh[6181], Fresh[6180]}), .outt ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, new_AGEMA_signal_2991, n2333}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2509 ( .ina ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, new_AGEMA_signal_1827, n2343}), .inb ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, new_AGEMA_signal_2730, n2342}), .clk ( clk ), .rnd ({Fresh[6199], Fresh[6198], Fresh[6197], Fresh[6196], Fresh[6195], Fresh[6194], Fresh[6193], Fresh[6192], Fresh[6191], Fresh[6190]}), .outt ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, new_AGEMA_signal_2997, n2345}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2526 ( .ina ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, new_AGEMA_signal_2733, n2358}), .inb ({new_AGEMA_signal_2324, new_AGEMA_signal_2323, new_AGEMA_signal_2322, n2357}), .clk ( clk ), .rnd ({Fresh[6209], Fresh[6208], Fresh[6207], Fresh[6206], Fresh[6205], Fresh[6204], Fresh[6203], Fresh[6202], Fresh[6201], Fresh[6200]}), .outt ({new_AGEMA_signal_3002, new_AGEMA_signal_3001, new_AGEMA_signal_3000, n2361}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2549 ( .ina ({new_AGEMA_signal_2336, new_AGEMA_signal_2335, new_AGEMA_signal_2334, n2387}), .inb ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, new_AGEMA_signal_2337, n2386}), .clk ( clk ), .rnd ({Fresh[6219], Fresh[6218], Fresh[6217], Fresh[6216], Fresh[6215], Fresh[6214], Fresh[6213], Fresh[6212], Fresh[6211], Fresh[6210]}), .outt ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, new_AGEMA_signal_2739, n2388}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2556 ( .ina ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .inb ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, new_AGEMA_signal_2742, n2392}), .clk ( clk ), .rnd ({Fresh[6229], Fresh[6228], Fresh[6227], Fresh[6226], Fresh[6225], Fresh[6224], Fresh[6223], Fresh[6222], Fresh[6221], Fresh[6220]}), .outt ({new_AGEMA_signal_3008, new_AGEMA_signal_3007, new_AGEMA_signal_3006, n2393}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2567 ( .ina ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .inb ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346, n2404}), .clk ( clk ), .rnd ({Fresh[6239], Fresh[6238], Fresh[6237], Fresh[6236], Fresh[6235], Fresh[6234], Fresh[6233], Fresh[6232], Fresh[6231], Fresh[6230]}), .outt ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, new_AGEMA_signal_2745, n2405}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2571 ( .ina ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, new_AGEMA_signal_2748, n2409}), .inb ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .clk ( clk ), .rnd ({Fresh[6249], Fresh[6248], Fresh[6247], Fresh[6246], Fresh[6245], Fresh[6244], Fresh[6243], Fresh[6242], Fresh[6241], Fresh[6240]}), .outt ({new_AGEMA_signal_3014, new_AGEMA_signal_3013, new_AGEMA_signal_3012, n2410}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2576 ( .ina ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .inb ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, new_AGEMA_signal_2751, n2414}), .clk ( clk ), .rnd ({Fresh[6259], Fresh[6258], Fresh[6257], Fresh[6256], Fresh[6255], Fresh[6254], Fresh[6253], Fresh[6252], Fresh[6251], Fresh[6250]}), .outt ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, new_AGEMA_signal_3015, n2421}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2579 ( .ina ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, n2418}), .inb ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .clk ( clk ), .rnd ({Fresh[6269], Fresh[6268], Fresh[6267], Fresh[6266], Fresh[6265], Fresh[6264], Fresh[6263], Fresh[6262], Fresh[6261], Fresh[6260]}), .outt ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, new_AGEMA_signal_2754, n2419}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2590 ( .ina ({new_AGEMA_signal_2360, new_AGEMA_signal_2359, new_AGEMA_signal_2358, n2433}), .inb ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, new_AGEMA_signal_2757, n2432}), .clk ( clk ), .rnd ({Fresh[6279], Fresh[6278], Fresh[6277], Fresh[6276], Fresh[6275], Fresh[6274], Fresh[6273], Fresh[6272], Fresh[6271], Fresh[6270]}), .outt ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, new_AGEMA_signal_3021, n2436}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2604 ( .ina ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, new_AGEMA_signal_2760, n2449}), .inb ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, new_AGEMA_signal_2763, n2448}), .clk ( clk ), .rnd ({Fresh[6289], Fresh[6288], Fresh[6287], Fresh[6286], Fresh[6285], Fresh[6284], Fresh[6283], Fresh[6282], Fresh[6281], Fresh[6280]}), .outt ({new_AGEMA_signal_3026, new_AGEMA_signal_3025, new_AGEMA_signal_3024, n2450}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2610 ( .ina ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}), .inb ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, new_AGEMA_signal_2766, n2455}), .clk ( clk ), .rnd ({Fresh[6299], Fresh[6298], Fresh[6297], Fresh[6296], Fresh[6295], Fresh[6294], Fresh[6293], Fresh[6292], Fresh[6291], Fresh[6290]}), .outt ({new_AGEMA_signal_3029, new_AGEMA_signal_3028, new_AGEMA_signal_3027, n2456}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2613 ( .ina ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, new_AGEMA_signal_2769, n2460}), .inb ({new_AGEMA_signal_2288, new_AGEMA_signal_2287, new_AGEMA_signal_2286, n2459}), .clk ( clk ), .rnd ({Fresh[6309], Fresh[6308], Fresh[6307], Fresh[6306], Fresh[6305], Fresh[6304], Fresh[6303], Fresh[6302], Fresh[6301], Fresh[6300]}), .outt ({new_AGEMA_signal_3032, new_AGEMA_signal_3031, new_AGEMA_signal_3030, n2461}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2619 ( .ina ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, new_AGEMA_signal_1854, n2467}), .inb ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, n2466}), .clk ( clk ), .rnd ({Fresh[6319], Fresh[6318], Fresh[6317], Fresh[6316], Fresh[6315], Fresh[6314], Fresh[6313], Fresh[6312], Fresh[6311], Fresh[6310]}), .outt ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, new_AGEMA_signal_2772, n2469}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2630 ( .ina ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .inb ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, new_AGEMA_signal_2385, n2477}), .clk ( clk ), .rnd ({Fresh[6329], Fresh[6328], Fresh[6327], Fresh[6326], Fresh[6325], Fresh[6324], Fresh[6323], Fresh[6322], Fresh[6321], Fresh[6320]}), .outt ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, new_AGEMA_signal_2775, n2478}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2635 ( .ina ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, n2483}), .inb ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, new_AGEMA_signal_2778, n2482}), .clk ( clk ), .rnd ({Fresh[6339], Fresh[6338], Fresh[6337], Fresh[6336], Fresh[6335], Fresh[6334], Fresh[6333], Fresh[6332], Fresh[6331], Fresh[6330]}), .outt ({new_AGEMA_signal_3038, new_AGEMA_signal_3037, new_AGEMA_signal_3036, n2484}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2643 ( .ina ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, n2490}), .inb ({new_AGEMA_signal_1916, new_AGEMA_signal_1915, new_AGEMA_signal_1914, n2489}), .clk ( clk ), .rnd ({Fresh[6349], Fresh[6348], Fresh[6347], Fresh[6346], Fresh[6345], Fresh[6344], Fresh[6343], Fresh[6342], Fresh[6341], Fresh[6340]}), .outt ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, new_AGEMA_signal_2781, n2491}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2649 ( .ina ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, new_AGEMA_signal_1917, n2497}), .inb ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, new_AGEMA_signal_2784, n2496}), .clk ( clk ), .rnd ({Fresh[6359], Fresh[6358], Fresh[6357], Fresh[6356], Fresh[6355], Fresh[6354], Fresh[6353], Fresh[6352], Fresh[6351], Fresh[6350]}), .outt ({new_AGEMA_signal_3044, new_AGEMA_signal_3043, new_AGEMA_signal_3042, n2500}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2656 ( .ina ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, new_AGEMA_signal_3045, n2507}), .inb ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, new_AGEMA_signal_2397, n2506}), .clk ( clk ), .rnd ({Fresh[6369], Fresh[6368], Fresh[6367], Fresh[6366], Fresh[6365], Fresh[6364], Fresh[6363], Fresh[6362], Fresh[6361], Fresh[6360]}), .outt ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, new_AGEMA_signal_3240, n2508}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2670 ( .ina ({new_AGEMA_signal_3050, new_AGEMA_signal_3049, new_AGEMA_signal_3048, n2525}), .inb ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, new_AGEMA_signal_2793, n2524}), .clk ( clk ), .rnd ({Fresh[6379], Fresh[6378], Fresh[6377], Fresh[6376], Fresh[6375], Fresh[6374], Fresh[6373], Fresh[6372], Fresh[6371], Fresh[6370]}), .outt ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, new_AGEMA_signal_3243, n2526}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2679 ( .ina ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, new_AGEMA_signal_2796, n2537}), .inb ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, new_AGEMA_signal_2799, n2536}), .clk ( clk ), .rnd ({Fresh[6389], Fresh[6388], Fresh[6387], Fresh[6386], Fresh[6385], Fresh[6384], Fresh[6383], Fresh[6382], Fresh[6381], Fresh[6380]}), .outt ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, new_AGEMA_signal_3051, n2539}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2682 ( .ina ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, new_AGEMA_signal_2634, n2543}), .inb ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, new_AGEMA_signal_2415, n2542}), .clk ( clk ), .rnd ({Fresh[6399], Fresh[6398], Fresh[6397], Fresh[6396], Fresh[6395], Fresh[6394], Fresh[6393], Fresh[6392], Fresh[6391], Fresh[6390]}), .outt ({new_AGEMA_signal_3056, new_AGEMA_signal_3055, new_AGEMA_signal_3054, n2548}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2694 ( .ina ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, new_AGEMA_signal_2424, n2558}), .inb ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, new_AGEMA_signal_2802, n2557}), .clk ( clk ), .rnd ({Fresh[6409], Fresh[6408], Fresh[6407], Fresh[6406], Fresh[6405], Fresh[6404], Fresh[6403], Fresh[6402], Fresh[6401], Fresh[6400]}), .outt ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, new_AGEMA_signal_3057, n2568}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2700 ( .ina ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, new_AGEMA_signal_2430, n2566}), .inb ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, new_AGEMA_signal_2805, n2565}), .clk ( clk ), .rnd ({Fresh[6419], Fresh[6418], Fresh[6417], Fresh[6416], Fresh[6415], Fresh[6414], Fresh[6413], Fresh[6412], Fresh[6411], Fresh[6410]}), .outt ({new_AGEMA_signal_3062, new_AGEMA_signal_3061, new_AGEMA_signal_3060, n2567}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2710 ( .ina ({new_AGEMA_signal_1946, new_AGEMA_signal_1945, new_AGEMA_signal_1944, n2581}), .inb ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, new_AGEMA_signal_2811, n2580}), .clk ( clk ), .rnd ({Fresh[6429], Fresh[6428], Fresh[6427], Fresh[6426], Fresh[6425], Fresh[6424], Fresh[6423], Fresh[6422], Fresh[6421], Fresh[6420]}), .outt ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, new_AGEMA_signal_3063, n2583}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2728 ( .ina ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, n2603}), .inb ({new_AGEMA_signal_1964, new_AGEMA_signal_1963, new_AGEMA_signal_1962, n2602}), .clk ( clk ), .rnd ({Fresh[6439], Fresh[6438], Fresh[6437], Fresh[6436], Fresh[6435], Fresh[6434], Fresh[6433], Fresh[6432], Fresh[6431], Fresh[6430]}), .outt ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, new_AGEMA_signal_2814, n2604}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2739 ( .ina ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, new_AGEMA_signal_2457, n2620}), .inb ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, new_AGEMA_signal_2817, n2619}), .clk ( clk ), .rnd ({Fresh[6449], Fresh[6448], Fresh[6447], Fresh[6446], Fresh[6445], Fresh[6444], Fresh[6443], Fresh[6442], Fresh[6441], Fresh[6440]}), .outt ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, new_AGEMA_signal_3069, n2621}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2745 ( .ina ({new_AGEMA_signal_1478, new_AGEMA_signal_1477, new_AGEMA_signal_1476, n2629}), .inb ({new_AGEMA_signal_2822, new_AGEMA_signal_2821, new_AGEMA_signal_2820, n2628}), .clk ( clk ), .rnd ({Fresh[6459], Fresh[6458], Fresh[6457], Fresh[6456], Fresh[6455], Fresh[6454], Fresh[6453], Fresh[6452], Fresh[6451], Fresh[6450]}), .outt ({new_AGEMA_signal_3074, new_AGEMA_signal_3073, new_AGEMA_signal_3072, n2633}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2756 ( .ina ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, new_AGEMA_signal_2823, n2649}), .inb ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, new_AGEMA_signal_2469, n2648}), .clk ( clk ), .rnd ({Fresh[6469], Fresh[6468], Fresh[6467], Fresh[6466], Fresh[6465], Fresh[6464], Fresh[6463], Fresh[6462], Fresh[6461], Fresh[6460]}), .outt ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, new_AGEMA_signal_3075, n2660}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2759 ( .ina ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, new_AGEMA_signal_1983, n2653}), .inb ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, new_AGEMA_signal_2604, n2652}), .clk ( clk ), .rnd ({Fresh[6479], Fresh[6478], Fresh[6477], Fresh[6476], Fresh[6475], Fresh[6474], Fresh[6473], Fresh[6472], Fresh[6471], Fresh[6470]}), .outt ({new_AGEMA_signal_3080, new_AGEMA_signal_3079, new_AGEMA_signal_3078, n2656}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2766 ( .ina ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, new_AGEMA_signal_2055, n2665}), .inb ({new_AGEMA_signal_2828, new_AGEMA_signal_2827, new_AGEMA_signal_2826, n2664}), .clk ( clk ), .rnd ({Fresh[6489], Fresh[6488], Fresh[6487], Fresh[6486], Fresh[6485], Fresh[6484], Fresh[6483], Fresh[6482], Fresh[6481], Fresh[6480]}), .outt ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, new_AGEMA_signal_3081, n2666}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2774 ( .ina ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, new_AGEMA_signal_2829, n2681}), .inb ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, new_AGEMA_signal_2478, n2680}), .clk ( clk ), .rnd ({Fresh[6499], Fresh[6498], Fresh[6497], Fresh[6496], Fresh[6495], Fresh[6494], Fresh[6493], Fresh[6492], Fresh[6491], Fresh[6490]}), .outt ({new_AGEMA_signal_3086, new_AGEMA_signal_3085, new_AGEMA_signal_3084, n2706}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2777 ( .ina ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, new_AGEMA_signal_2703, n2686}), .inb ({new_AGEMA_signal_2834, new_AGEMA_signal_2833, new_AGEMA_signal_2832, n2685}), .clk ( clk ), .rnd ({Fresh[6509], Fresh[6508], Fresh[6507], Fresh[6506], Fresh[6505], Fresh[6504], Fresh[6503], Fresh[6502], Fresh[6501], Fresh[6500]}), .outt ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, new_AGEMA_signal_3087, n2704}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2781 ( .ina ({new_AGEMA_signal_2840, new_AGEMA_signal_2839, new_AGEMA_signal_2838, n2692}), .inb ({new_AGEMA_signal_1994, new_AGEMA_signal_1993, new_AGEMA_signal_1992, n2691}), .clk ( clk ), .rnd ({Fresh[6519], Fresh[6518], Fresh[6517], Fresh[6516], Fresh[6515], Fresh[6514], Fresh[6513], Fresh[6512], Fresh[6511], Fresh[6510]}), .outt ({new_AGEMA_signal_3092, new_AGEMA_signal_3091, new_AGEMA_signal_3090, n2696}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2794 ( .ina ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, new_AGEMA_signal_2484, n2717}), .inb ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, new_AGEMA_signal_2841, n2716}), .clk ( clk ), .rnd ({Fresh[6529], Fresh[6528], Fresh[6527], Fresh[6526], Fresh[6525], Fresh[6524], Fresh[6523], Fresh[6522], Fresh[6521], Fresh[6520]}), .outt ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, new_AGEMA_signal_3093, n2718}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2801 ( .ina ({new_AGEMA_signal_2846, new_AGEMA_signal_2845, new_AGEMA_signal_2844, n2729}), .inb ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, new_AGEMA_signal_2487, n2728}), .clk ( clk ), .rnd ({Fresh[6539], Fresh[6538], Fresh[6537], Fresh[6536], Fresh[6535], Fresh[6534], Fresh[6533], Fresh[6532], Fresh[6531], Fresh[6530]}), .outt ({new_AGEMA_signal_3098, new_AGEMA_signal_3097, new_AGEMA_signal_3096, n2730}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2805 ( .ina ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, n2736}), .inb ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, new_AGEMA_signal_2847, n2735}), .clk ( clk ), .rnd ({Fresh[6549], Fresh[6548], Fresh[6547], Fresh[6546], Fresh[6545], Fresh[6544], Fresh[6543], Fresh[6542], Fresh[6541], Fresh[6540]}), .outt ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, new_AGEMA_signal_3099, n2745}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2809 ( .ina ({new_AGEMA_signal_2852, new_AGEMA_signal_2851, new_AGEMA_signal_2850, n2743}), .inb ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .clk ( clk ), .rnd ({Fresh[6559], Fresh[6558], Fresh[6557], Fresh[6556], Fresh[6555], Fresh[6554], Fresh[6553], Fresh[6552], Fresh[6551], Fresh[6550]}), .outt ({new_AGEMA_signal_3104, new_AGEMA_signal_3103, new_AGEMA_signal_3102, n2744}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2814 ( .ina ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, new_AGEMA_signal_2691, n2752}), .inb ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, new_AGEMA_signal_2496, n2751}), .clk ( clk ), .rnd ({Fresh[6569], Fresh[6568], Fresh[6567], Fresh[6566], Fresh[6565], Fresh[6564], Fresh[6563], Fresh[6562], Fresh[6561], Fresh[6560]}), .outt ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, new_AGEMA_signal_3105, n2759}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2821 ( .ina ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .inb ({new_AGEMA_signal_2858, new_AGEMA_signal_2857, new_AGEMA_signal_2856, n2764}), .clk ( clk ), .rnd ({Fresh[6579], Fresh[6578], Fresh[6577], Fresh[6576], Fresh[6575], Fresh[6574], Fresh[6573], Fresh[6572], Fresh[6571], Fresh[6570]}), .outt ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, new_AGEMA_signal_3108, n2771}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2833 ( .ina ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, new_AGEMA_signal_2514, n2788}), .inb ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, new_AGEMA_signal_2025, n2787}), .clk ( clk ), .rnd ({Fresh[6589], Fresh[6588], Fresh[6587], Fresh[6586], Fresh[6585], Fresh[6584], Fresh[6583], Fresh[6582], Fresh[6581], Fresh[6580]}), .outt ({new_AGEMA_signal_2864, new_AGEMA_signal_2863, new_AGEMA_signal_2862, n2798}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2850 ( .ina ({new_AGEMA_signal_2870, new_AGEMA_signal_2869, new_AGEMA_signal_2868, n2822}), .inb ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, new_AGEMA_signal_2523, n2821}), .clk ( clk ), .rnd ({Fresh[6599], Fresh[6598], Fresh[6597], Fresh[6596], Fresh[6595], Fresh[6594], Fresh[6593], Fresh[6592], Fresh[6591], Fresh[6590]}), .outt ({new_AGEMA_signal_3116, new_AGEMA_signal_3115, new_AGEMA_signal_3114, n2826}) ) ;

    /* cells in depth 11 */

    /* cells in depth 12 */
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2001 ( .ina ({new_AGEMA_signal_2876, new_AGEMA_signal_2875, new_AGEMA_signal_2874, n1932}), .inb ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, n2577}), .clk ( clk ), .rnd ({Fresh[6609], Fresh[6608], Fresh[6607], Fresh[6606], Fresh[6605], Fresh[6604], Fresh[6603], Fresh[6602], Fresh[6601], Fresh[6600]}), .outt ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, new_AGEMA_signal_3117, n1933}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2051 ( .ina ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, new_AGEMA_signal_2067, n1956}), .inb ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, new_AGEMA_signal_2883, n1955}), .clk ( clk ), .rnd ({Fresh[6619], Fresh[6618], Fresh[6617], Fresh[6616], Fresh[6615], Fresh[6614], Fresh[6613], Fresh[6612], Fresh[6611], Fresh[6610]}), .outt ({new_AGEMA_signal_3122, new_AGEMA_signal_3121, new_AGEMA_signal_3120, n1958}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2067 ( .ina ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, new_AGEMA_signal_2553, n1967}), .inb ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, new_AGEMA_signal_1005, n2595}), .clk ( clk ), .rnd ({Fresh[6629], Fresh[6628], Fresh[6627], Fresh[6626], Fresh[6625], Fresh[6624], Fresh[6623], Fresh[6622], Fresh[6621], Fresh[6620]}), .outt ({new_AGEMA_signal_2888, new_AGEMA_signal_2887, new_AGEMA_signal_2886, n1990}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2104 ( .ina ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, new_AGEMA_signal_2562, n1978}), .inb ({new_AGEMA_signal_2894, new_AGEMA_signal_2893, new_AGEMA_signal_2892, n1977}), .clk ( clk ), .rnd ({Fresh[6639], Fresh[6638], Fresh[6637], Fresh[6636], Fresh[6635], Fresh[6634], Fresh[6633], Fresh[6632], Fresh[6631], Fresh[6630]}), .outt ({new_AGEMA_signal_3128, new_AGEMA_signal_3127, new_AGEMA_signal_3126, n1982}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2128 ( .ina ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .inb ({new_AGEMA_signal_2900, new_AGEMA_signal_2899, new_AGEMA_signal_2898, n1998}), .clk ( clk ), .rnd ({Fresh[6649], Fresh[6648], Fresh[6647], Fresh[6646], Fresh[6645], Fresh[6644], Fresh[6643], Fresh[6642], Fresh[6641], Fresh[6640]}), .outt ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, new_AGEMA_signal_3129, n1999}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2148 ( .ina ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, new_AGEMA_signal_2901, n2010}), .inb ({new_AGEMA_signal_1604, new_AGEMA_signal_1603, new_AGEMA_signal_1602, n2009}), .clk ( clk ), .rnd ({Fresh[6659], Fresh[6658], Fresh[6657], Fresh[6656], Fresh[6655], Fresh[6654], Fresh[6653], Fresh[6652], Fresh[6651], Fresh[6650]}), .outt ({new_AGEMA_signal_3134, new_AGEMA_signal_3133, new_AGEMA_signal_3132, n2011}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2165 ( .ina ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, new_AGEMA_signal_2583, n2024}), .inb ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, new_AGEMA_signal_1614, n2023}), .clk ( clk ), .rnd ({Fresh[6669], Fresh[6668], Fresh[6667], Fresh[6666], Fresh[6665], Fresh[6664], Fresh[6663], Fresh[6662], Fresh[6661], Fresh[6660]}), .outt ({new_AGEMA_signal_2906, new_AGEMA_signal_2905, new_AGEMA_signal_2904, n2025}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2179 ( .ina ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, new_AGEMA_signal_2907, n2035}), .inb ({new_AGEMA_signal_1334, new_AGEMA_signal_1333, new_AGEMA_signal_1332, n2034}), .clk ( clk ), .rnd ({Fresh[6679], Fresh[6678], Fresh[6677], Fresh[6676], Fresh[6675], Fresh[6674], Fresh[6673], Fresh[6672], Fresh[6671], Fresh[6670]}), .outt ({new_AGEMA_signal_3140, new_AGEMA_signal_3139, new_AGEMA_signal_3138, n2036}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2196 ( .ina ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, new_AGEMA_signal_2913, n2048}), .inb ({new_AGEMA_signal_2918, new_AGEMA_signal_2917, new_AGEMA_signal_2916, n2047}), .clk ( clk ), .rnd ({Fresh[6689], Fresh[6688], Fresh[6687], Fresh[6686], Fresh[6685], Fresh[6684], Fresh[6683], Fresh[6682], Fresh[6681], Fresh[6680]}), .outt ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, new_AGEMA_signal_3141, n2049}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2207 ( .ina ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .inb ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, new_AGEMA_signal_2919, n2059}), .clk ( clk ), .rnd ({Fresh[6699], Fresh[6698], Fresh[6697], Fresh[6696], Fresh[6695], Fresh[6694], Fresh[6693], Fresh[6692], Fresh[6691], Fresh[6690]}), .outt ({new_AGEMA_signal_3146, new_AGEMA_signal_3145, new_AGEMA_signal_3144, n2072}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2214 ( .ina ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .inb ({new_AGEMA_signal_2924, new_AGEMA_signal_2923, new_AGEMA_signal_2922, n2064}), .clk ( clk ), .rnd ({Fresh[6709], Fresh[6708], Fresh[6707], Fresh[6706], Fresh[6705], Fresh[6704], Fresh[6703], Fresh[6702], Fresh[6701], Fresh[6700]}), .outt ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, new_AGEMA_signal_3147, n2067}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2230 ( .ina ({new_AGEMA_signal_1040, new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2699}), .inb ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, new_AGEMA_signal_2925, n2077}), .clk ( clk ), .rnd ({Fresh[6719], Fresh[6718], Fresh[6717], Fresh[6716], Fresh[6715], Fresh[6714], Fresh[6713], Fresh[6712], Fresh[6711], Fresh[6710]}), .outt ({new_AGEMA_signal_3152, new_AGEMA_signal_3151, new_AGEMA_signal_3150, n2078}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2250 ( .ina ({new_AGEMA_signal_2618, new_AGEMA_signal_2617, new_AGEMA_signal_2616, n2091}), .inb ({new_AGEMA_signal_2930, new_AGEMA_signal_2929, new_AGEMA_signal_2928, n2158}), .clk ( clk ), .rnd ({Fresh[6729], Fresh[6728], Fresh[6727], Fresh[6726], Fresh[6725], Fresh[6724], Fresh[6723], Fresh[6722], Fresh[6721], Fresh[6720]}), .outt ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, new_AGEMA_signal_3153, n2097}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2257 ( .ina ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, new_AGEMA_signal_2931, n2095}), .inb ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, new_AGEMA_signal_2181, n2094}), .clk ( clk ), .rnd ({Fresh[6739], Fresh[6738], Fresh[6737], Fresh[6736], Fresh[6735], Fresh[6734], Fresh[6733], Fresh[6732], Fresh[6731], Fresh[6730]}), .outt ({new_AGEMA_signal_3158, new_AGEMA_signal_3157, new_AGEMA_signal_3156, n2096}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2275 ( .ina ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .inb ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, new_AGEMA_signal_3159, n2117}), .clk ( clk ), .rnd ({Fresh[6749], Fresh[6748], Fresh[6747], Fresh[6746], Fresh[6745], Fresh[6744], Fresh[6743], Fresh[6742], Fresh[6741], Fresh[6740]}), .outt ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, new_AGEMA_signal_3321, n2128}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2285 ( .ina ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, new_AGEMA_signal_2937, n2123}), .inb ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, new_AGEMA_signal_1695, n2122}), .clk ( clk ), .rnd ({Fresh[6759], Fresh[6758], Fresh[6757], Fresh[6756], Fresh[6755], Fresh[6754], Fresh[6753], Fresh[6752], Fresh[6751], Fresh[6750]}), .outt ({new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162, n2124}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2301 ( .ina ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, new_AGEMA_signal_2634, n2543}), .inb ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, new_AGEMA_signal_2637, n2135}), .clk ( clk ), .rnd ({Fresh[6769], Fresh[6768], Fresh[6767], Fresh[6766], Fresh[6765], Fresh[6764], Fresh[6763], Fresh[6762], Fresh[6761], Fresh[6760]}), .outt ({new_AGEMA_signal_2942, new_AGEMA_signal_2941, new_AGEMA_signal_2940, n2148}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2310 ( .ina ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, new_AGEMA_signal_1713, n2220}), .inb ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, new_AGEMA_signal_2943, n2141}), .clk ( clk ), .rnd ({Fresh[6779], Fresh[6778], Fresh[6777], Fresh[6776], Fresh[6775], Fresh[6774], Fresh[6773], Fresh[6772], Fresh[6771], Fresh[6770]}), .outt ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, new_AGEMA_signal_3165, n2142}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2325 ( .ina ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, new_AGEMA_signal_2646, n2159}), .inb ({new_AGEMA_signal_2930, new_AGEMA_signal_2929, new_AGEMA_signal_2928, n2158}), .clk ( clk ), .rnd ({Fresh[6789], Fresh[6788], Fresh[6787], Fresh[6786], Fresh[6785], Fresh[6784], Fresh[6783], Fresh[6782], Fresh[6781], Fresh[6780]}), .outt ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, new_AGEMA_signal_3168, n2168}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2332 ( .ina ({new_AGEMA_signal_2948, new_AGEMA_signal_2947, new_AGEMA_signal_2946, n2166}), .inb ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, new_AGEMA_signal_2652, n2165}), .clk ( clk ), .rnd ({Fresh[6799], Fresh[6798], Fresh[6797], Fresh[6796], Fresh[6795], Fresh[6794], Fresh[6793], Fresh[6792], Fresh[6791], Fresh[6790]}), .outt ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, new_AGEMA_signal_3171, n2167}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2347 ( .ina ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, new_AGEMA_signal_2223, n2181}), .inb ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, new_AGEMA_signal_2949, n2180}), .clk ( clk ), .rnd ({Fresh[6809], Fresh[6808], Fresh[6807], Fresh[6806], Fresh[6805], Fresh[6804], Fresh[6803], Fresh[6802], Fresh[6801], Fresh[6800]}), .outt ({new_AGEMA_signal_3176, new_AGEMA_signal_3175, new_AGEMA_signal_3174, n2184}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2361 ( .ina ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, new_AGEMA_signal_2229, n2195}), .inb ({new_AGEMA_signal_2954, new_AGEMA_signal_2953, new_AGEMA_signal_2952, n2194}), .clk ( clk ), .rnd ({Fresh[6819], Fresh[6818], Fresh[6817], Fresh[6816], Fresh[6815], Fresh[6814], Fresh[6813], Fresh[6812], Fresh[6811], Fresh[6810]}), .outt ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, new_AGEMA_signal_3177, n2197}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2373 ( .ina ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}), .inb ({new_AGEMA_signal_3182, new_AGEMA_signal_3181, new_AGEMA_signal_3180, n2204}), .clk ( clk ), .rnd ({Fresh[6829], Fresh[6828], Fresh[6827], Fresh[6826], Fresh[6825], Fresh[6824], Fresh[6823], Fresh[6822], Fresh[6821], Fresh[6820]}), .outt ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, new_AGEMA_signal_3339, n2205}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2390 ( .ina ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, n2828}), .inb ({new_AGEMA_signal_2960, new_AGEMA_signal_2959, new_AGEMA_signal_2958, n2225}), .clk ( clk ), .rnd ({Fresh[6839], Fresh[6838], Fresh[6837], Fresh[6836], Fresh[6835], Fresh[6834], Fresh[6833], Fresh[6832], Fresh[6831], Fresh[6830]}), .outt ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, new_AGEMA_signal_3183, n2232}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2395 ( .ina ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, new_AGEMA_signal_2673, n2230}), .inb ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}), .clk ( clk ), .rnd ({Fresh[6849], Fresh[6848], Fresh[6847], Fresh[6846], Fresh[6845], Fresh[6844], Fresh[6843], Fresh[6842], Fresh[6841], Fresh[6840]}), .outt ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, new_AGEMA_signal_2961, n2231}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2401 ( .ina ({new_AGEMA_signal_1763, new_AGEMA_signal_1762, new_AGEMA_signal_1761, n2237}), .inb ({new_AGEMA_signal_3188, new_AGEMA_signal_3187, new_AGEMA_signal_3186, n2236}), .clk ( clk ), .rnd ({Fresh[6859], Fresh[6858], Fresh[6857], Fresh[6856], Fresh[6855], Fresh[6854], Fresh[6853], Fresh[6852], Fresh[6851], Fresh[6850]}), .outt ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, new_AGEMA_signal_3345, n2239}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2413 ( .ina ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, new_AGEMA_signal_2256, n2248}), .inb ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, new_AGEMA_signal_2967, n2247}), .clk ( clk ), .rnd ({Fresh[6869], Fresh[6868], Fresh[6867], Fresh[6866], Fresh[6865], Fresh[6864], Fresh[6863], Fresh[6862], Fresh[6861], Fresh[6860]}), .outt ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, new_AGEMA_signal_3189, n2250}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2428 ( .ina ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .inb ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, new_AGEMA_signal_2973, n2264}), .clk ( clk ), .rnd ({Fresh[6879], Fresh[6878], Fresh[6877], Fresh[6876], Fresh[6875], Fresh[6874], Fresh[6873], Fresh[6872], Fresh[6871], Fresh[6870]}), .outt ({new_AGEMA_signal_3194, new_AGEMA_signal_3193, new_AGEMA_signal_3192, n2276}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2439 ( .ina ({new_AGEMA_signal_2978, new_AGEMA_signal_2977, new_AGEMA_signal_2976, n2271}), .inb ({new_AGEMA_signal_2276, new_AGEMA_signal_2275, new_AGEMA_signal_2274, n2270}), .clk ( clk ), .rnd ({Fresh[6889], Fresh[6888], Fresh[6887], Fresh[6886], Fresh[6885], Fresh[6884], Fresh[6883], Fresh[6882], Fresh[6881], Fresh[6880]}), .outt ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, new_AGEMA_signal_3195, n2272}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2454 ( .ina ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, new_AGEMA_signal_2697, n2286}), .inb ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, new_AGEMA_signal_2700, n2285}), .clk ( clk ), .rnd ({Fresh[6899], Fresh[6898], Fresh[6897], Fresh[6896], Fresh[6895], Fresh[6894], Fresh[6893], Fresh[6892], Fresh[6891], Fresh[6890]}), .outt ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, new_AGEMA_signal_2979, n2306}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2468 ( .ina ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, new_AGEMA_signal_2985, n2295}), .inb ({new_AGEMA_signal_1808, new_AGEMA_signal_1807, new_AGEMA_signal_1806, n2294}), .clk ( clk ), .rnd ({Fresh[6909], Fresh[6908], Fresh[6907], Fresh[6906], Fresh[6905], Fresh[6904], Fresh[6903], Fresh[6902], Fresh[6901], Fresh[6900]}), .outt ({new_AGEMA_signal_3200, new_AGEMA_signal_3199, new_AGEMA_signal_3198, n2296}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2489 ( .ina ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, new_AGEMA_signal_2301, n2323}), .inb ({new_AGEMA_signal_2990, new_AGEMA_signal_2989, new_AGEMA_signal_2988, n2322}), .clk ( clk ), .rnd ({Fresh[6919], Fresh[6918], Fresh[6917], Fresh[6916], Fresh[6915], Fresh[6914], Fresh[6913], Fresh[6912], Fresh[6911], Fresh[6910]}), .outt ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, new_AGEMA_signal_3201, n2324}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2500 ( .ina ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, new_AGEMA_signal_2307, n2334}), .inb ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, new_AGEMA_signal_2991, n2333}), .clk ( clk ), .rnd ({Fresh[6929], Fresh[6928], Fresh[6927], Fresh[6926], Fresh[6925], Fresh[6924], Fresh[6923], Fresh[6922], Fresh[6921], Fresh[6920]}), .outt ({new_AGEMA_signal_3206, new_AGEMA_signal_3205, new_AGEMA_signal_3204, n2337}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2511 ( .ina ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, new_AGEMA_signal_2997, n2345}), .inb ({new_AGEMA_signal_1835, new_AGEMA_signal_1834, new_AGEMA_signal_1833, n2344}), .clk ( clk ), .rnd ({Fresh[6939], Fresh[6938], Fresh[6937], Fresh[6936], Fresh[6935], Fresh[6934], Fresh[6933], Fresh[6932], Fresh[6931], Fresh[6930]}), .outt ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, new_AGEMA_signal_3207, n2350}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2528 ( .ina ({new_AGEMA_signal_3002, new_AGEMA_signal_3001, new_AGEMA_signal_3000, n2361}), .inb ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, new_AGEMA_signal_2325, n2360}), .clk ( clk ), .rnd ({Fresh[6949], Fresh[6948], Fresh[6947], Fresh[6946], Fresh[6945], Fresh[6944], Fresh[6943], Fresh[6942], Fresh[6941], Fresh[6940]}), .outt ({new_AGEMA_signal_3212, new_AGEMA_signal_3211, new_AGEMA_signal_3210, n2362}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2550 ( .ina ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, new_AGEMA_signal_1854, n2467}), .inb ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, new_AGEMA_signal_2739, n2388}), .clk ( clk ), .rnd ({Fresh[6959], Fresh[6958], Fresh[6957], Fresh[6956], Fresh[6955], Fresh[6954], Fresh[6953], Fresh[6952], Fresh[6951], Fresh[6950]}), .outt ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003, n2389}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2557 ( .ina ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, new_AGEMA_signal_1863, n2394}), .inb ({new_AGEMA_signal_3008, new_AGEMA_signal_3007, new_AGEMA_signal_3006, n2393}), .clk ( clk ), .rnd ({Fresh[6969], Fresh[6968], Fresh[6967], Fresh[6966], Fresh[6965], Fresh[6964], Fresh[6963], Fresh[6962], Fresh[6961], Fresh[6960]}), .outt ({new_AGEMA_signal_3218, new_AGEMA_signal_3217, new_AGEMA_signal_3216, n2397}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2568 ( .ina ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, new_AGEMA_signal_2343, n2406}), .inb ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, new_AGEMA_signal_2745, n2405}), .clk ( clk ), .rnd ({Fresh[6979], Fresh[6978], Fresh[6977], Fresh[6976], Fresh[6975], Fresh[6974], Fresh[6973], Fresh[6972], Fresh[6971], Fresh[6970]}), .outt ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, new_AGEMA_signal_3009, n2411}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2580 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, new_AGEMA_signal_2754, n2419}), .clk ( clk ), .rnd ({Fresh[6989], Fresh[6988], Fresh[6987], Fresh[6986], Fresh[6985], Fresh[6984], Fresh[6983], Fresh[6982], Fresh[6981], Fresh[6980]}), .outt ({new_AGEMA_signal_3020, new_AGEMA_signal_3019, new_AGEMA_signal_3018, n2420}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2593 ( .ina ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, new_AGEMA_signal_3021, n2436}), .inb ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, new_AGEMA_signal_2364, n2435}), .clk ( clk ), .rnd ({Fresh[6999], Fresh[6998], Fresh[6997], Fresh[6996], Fresh[6995], Fresh[6994], Fresh[6993], Fresh[6992], Fresh[6991], Fresh[6990]}), .outt ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, new_AGEMA_signal_3225, n2440}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2614 ( .ina ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_3032, new_AGEMA_signal_3031, new_AGEMA_signal_3030, n2461}), .clk ( clk ), .rnd ({Fresh[7009], Fresh[7008], Fresh[7007], Fresh[7006], Fresh[7005], Fresh[7004], Fresh[7003], Fresh[7002], Fresh[7001], Fresh[7000]}), .outt ({new_AGEMA_signal_3230, new_AGEMA_signal_3229, new_AGEMA_signal_3228, n2516}) ) ;
    mux2_HPC1 #(.security_order(3), .pipeline(0)) U2621 ( .ins ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .inb ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, new_AGEMA_signal_2772, n2469}), .ina ({new_AGEMA_signal_1448, new_AGEMA_signal_1447, new_AGEMA_signal_1446, n2468}), .clk ( clk ), .rnd ({Fresh[7019], Fresh[7018], Fresh[7017], Fresh[7016], Fresh[7015], Fresh[7014], Fresh[7013], Fresh[7012], Fresh[7011], Fresh[7010]}), .outt ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, new_AGEMA_signal_3033, n2471}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2636 ( .ina ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}), .inb ({new_AGEMA_signal_3038, new_AGEMA_signal_3037, new_AGEMA_signal_3036, n2484}), .clk ( clk ), .rnd ({Fresh[7029], Fresh[7028], Fresh[7027], Fresh[7026], Fresh[7025], Fresh[7024], Fresh[7023], Fresh[7022], Fresh[7021], Fresh[7020]}), .outt ({new_AGEMA_signal_3236, new_AGEMA_signal_3235, new_AGEMA_signal_3234, n2485}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2644 ( .ina ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .inb ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, new_AGEMA_signal_2781, n2491}), .clk ( clk ), .rnd ({Fresh[7039], Fresh[7038], Fresh[7037], Fresh[7036], Fresh[7035], Fresh[7034], Fresh[7033], Fresh[7032], Fresh[7031], Fresh[7030]}), .outt ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, new_AGEMA_signal_3039, n2502}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2651 ( .ina ({new_AGEMA_signal_3044, new_AGEMA_signal_3043, new_AGEMA_signal_3042, n2500}), .inb ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, new_AGEMA_signal_1923, n2499}), .clk ( clk ), .rnd ({Fresh[7049], Fresh[7048], Fresh[7047], Fresh[7046], Fresh[7045], Fresh[7044], Fresh[7043], Fresh[7042], Fresh[7041], Fresh[7040]}), .outt ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, new_AGEMA_signal_3237, n2501}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2657 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, new_AGEMA_signal_3240, n2508}), .clk ( clk ), .rnd ({Fresh[7059], Fresh[7058], Fresh[7057], Fresh[7056], Fresh[7055], Fresh[7054], Fresh[7053], Fresh[7052], Fresh[7051], Fresh[7050]}), .outt ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, new_AGEMA_signal_3387, n2509}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2671 ( .ina ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, n2785}), .inb ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, new_AGEMA_signal_3243, n2526}), .clk ( clk ), .rnd ({Fresh[7069], Fresh[7068], Fresh[7067], Fresh[7066], Fresh[7065], Fresh[7064], Fresh[7063], Fresh[7062], Fresh[7061], Fresh[7060]}), .outt ({new_AGEMA_signal_3392, new_AGEMA_signal_3391, new_AGEMA_signal_3390, n2527}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2680 ( .ina ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, new_AGEMA_signal_3051, n2539}), .inb ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, new_AGEMA_signal_1071, n2538}), .clk ( clk ), .rnd ({Fresh[7079], Fresh[7078], Fresh[7077], Fresh[7076], Fresh[7075], Fresh[7074], Fresh[7073], Fresh[7072], Fresh[7071], Fresh[7070]}), .outt ({new_AGEMA_signal_3248, new_AGEMA_signal_3247, new_AGEMA_signal_3246, n2550}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2685 ( .ina ({new_AGEMA_signal_3056, new_AGEMA_signal_3055, new_AGEMA_signal_3054, n2548}), .inb ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, new_AGEMA_signal_2418, n2547}), .clk ( clk ), .rnd ({Fresh[7089], Fresh[7088], Fresh[7087], Fresh[7086], Fresh[7085], Fresh[7084], Fresh[7083], Fresh[7082], Fresh[7081], Fresh[7080]}), .outt ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, new_AGEMA_signal_3249, n2549}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2701 ( .ina ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, new_AGEMA_signal_3057, n2568}), .inb ({new_AGEMA_signal_3062, new_AGEMA_signal_3061, new_AGEMA_signal_3060, n2567}), .clk ( clk ), .rnd ({Fresh[7099], Fresh[7098], Fresh[7097], Fresh[7096], Fresh[7095], Fresh[7094], Fresh[7093], Fresh[7092], Fresh[7091], Fresh[7090]}), .outt ({new_AGEMA_signal_3254, new_AGEMA_signal_3253, new_AGEMA_signal_3252, n2569}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2712 ( .ina ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, new_AGEMA_signal_3063, n2583}), .inb ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, new_AGEMA_signal_2445, n2582}), .clk ( clk ), .rnd ({Fresh[7109], Fresh[7108], Fresh[7107], Fresh[7106], Fresh[7105], Fresh[7104], Fresh[7103], Fresh[7102], Fresh[7101], Fresh[7100]}), .outt ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, new_AGEMA_signal_3255, n2584}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2729 ( .ina ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, new_AGEMA_signal_2451, n2605}), .inb ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, new_AGEMA_signal_2814, n2604}), .clk ( clk ), .rnd ({Fresh[7119], Fresh[7118], Fresh[7117], Fresh[7116], Fresh[7115], Fresh[7114], Fresh[7113], Fresh[7112], Fresh[7111], Fresh[7110]}), .outt ({new_AGEMA_signal_3068, new_AGEMA_signal_3067, new_AGEMA_signal_3066, n2606}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2740 ( .ina ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .inb ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, new_AGEMA_signal_3069, n2621}), .clk ( clk ), .rnd ({Fresh[7129], Fresh[7128], Fresh[7127], Fresh[7126], Fresh[7125], Fresh[7124], Fresh[7123], Fresh[7122], Fresh[7121], Fresh[7120]}), .outt ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, new_AGEMA_signal_3261, n2622}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2747 ( .ina ({new_AGEMA_signal_3074, new_AGEMA_signal_3073, new_AGEMA_signal_3072, n2633}), .inb ({new_AGEMA_signal_1976, new_AGEMA_signal_1975, new_AGEMA_signal_1974, n2632}), .clk ( clk ), .rnd ({Fresh[7139], Fresh[7138], Fresh[7137], Fresh[7136], Fresh[7135], Fresh[7134], Fresh[7133], Fresh[7132], Fresh[7131], Fresh[7130]}), .outt ({new_AGEMA_signal_3266, new_AGEMA_signal_3265, new_AGEMA_signal_3264, n2634}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2761 ( .ina ({new_AGEMA_signal_3080, new_AGEMA_signal_3079, new_AGEMA_signal_3078, n2656}), .inb ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, new_AGEMA_signal_2472, n2655}), .clk ( clk ), .rnd ({Fresh[7149], Fresh[7148], Fresh[7147], Fresh[7146], Fresh[7145], Fresh[7144], Fresh[7143], Fresh[7142], Fresh[7141], Fresh[7140]}), .outt ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, new_AGEMA_signal_3267, n2657}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2783 ( .ina ({new_AGEMA_signal_3092, new_AGEMA_signal_3091, new_AGEMA_signal_3090, n2696}), .inb ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, new_AGEMA_signal_2481, n2695}), .clk ( clk ), .rnd ({Fresh[7159], Fresh[7158], Fresh[7157], Fresh[7156], Fresh[7155], Fresh[7154], Fresh[7153], Fresh[7152], Fresh[7151], Fresh[7150]}), .outt ({new_AGEMA_signal_3272, new_AGEMA_signal_3271, new_AGEMA_signal_3270, n2697}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2795 ( .ina ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .inb ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, new_AGEMA_signal_3093, n2718}), .clk ( clk ), .rnd ({Fresh[7169], Fresh[7168], Fresh[7167], Fresh[7166], Fresh[7165], Fresh[7164], Fresh[7163], Fresh[7162], Fresh[7161], Fresh[7160]}), .outt ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, new_AGEMA_signal_3273, n2808}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2802 ( .ina ({new_AGEMA_signal_3098, new_AGEMA_signal_3097, new_AGEMA_signal_3096, n2730}), .inb ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, n2809}), .clk ( clk ), .rnd ({Fresh[7179], Fresh[7178], Fresh[7177], Fresh[7176], Fresh[7175], Fresh[7174], Fresh[7173], Fresh[7172], Fresh[7171], Fresh[7170]}), .outt ({new_AGEMA_signal_3278, new_AGEMA_signal_3277, new_AGEMA_signal_3276, n2747}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2810 ( .ina ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, new_AGEMA_signal_3099, n2745}), .inb ({new_AGEMA_signal_3104, new_AGEMA_signal_3103, new_AGEMA_signal_3102, n2744}), .clk ( clk ), .rnd ({Fresh[7189], Fresh[7188], Fresh[7187], Fresh[7186], Fresh[7185], Fresh[7184], Fresh[7183], Fresh[7182], Fresh[7181], Fresh[7180]}), .outt ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, new_AGEMA_signal_3279, n2746}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2818 ( .ina ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, new_AGEMA_signal_3105, n2759}), .inb ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, new_AGEMA_signal_2853, n2758}), .clk ( clk ), .rnd ({Fresh[7199], Fresh[7198], Fresh[7197], Fresh[7196], Fresh[7195], Fresh[7194], Fresh[7193], Fresh[7192], Fresh[7191], Fresh[7190]}), .outt ({new_AGEMA_signal_3284, new_AGEMA_signal_3283, new_AGEMA_signal_3282, n2804}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2824 ( .ina ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, new_AGEMA_signal_3108, n2771}), .inb ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, new_AGEMA_signal_2505, n2770}), .clk ( clk ), .rnd ({Fresh[7209], Fresh[7208], Fresh[7207], Fresh[7206], Fresh[7205], Fresh[7204], Fresh[7203], Fresh[7202], Fresh[7201], Fresh[7200]}), .outt ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, new_AGEMA_signal_3285, n2802}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2838 ( .ina ({new_AGEMA_signal_2864, new_AGEMA_signal_2863, new_AGEMA_signal_2862, n2798}), .inb ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, new_AGEMA_signal_2865, n2797}), .clk ( clk ), .rnd ({Fresh[7219], Fresh[7218], Fresh[7217], Fresh[7216], Fresh[7215], Fresh[7214], Fresh[7213], Fresh[7212], Fresh[7211], Fresh[7210]}), .outt ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, new_AGEMA_signal_3111, n2799}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2852 ( .ina ({new_AGEMA_signal_3116, new_AGEMA_signal_3115, new_AGEMA_signal_3114, n2826}), .inb ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, new_AGEMA_signal_2040, n2825}), .clk ( clk ), .rnd ({Fresh[7229], Fresh[7228], Fresh[7227], Fresh[7226], Fresh[7225], Fresh[7224], Fresh[7223], Fresh[7222], Fresh[7221], Fresh[7220]}), .outt ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, new_AGEMA_signal_3291, n2827}) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2002 ( .ina ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, new_AGEMA_signal_2871, n1934}), .inb ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, new_AGEMA_signal_3117, n1933}), .clk ( clk ), .rnd ({Fresh[7239], Fresh[7238], Fresh[7237], Fresh[7236], Fresh[7235], Fresh[7234], Fresh[7233], Fresh[7232], Fresh[7231], Fresh[7230]}), .outt ({new_AGEMA_signal_3296, new_AGEMA_signal_3295, new_AGEMA_signal_3294, n1935}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2054 ( .ina ({new_AGEMA_signal_3122, new_AGEMA_signal_3121, new_AGEMA_signal_3120, n1958}), .inb ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, new_AGEMA_signal_1263, n1957}), .clk ( clk ), .rnd ({Fresh[7249], Fresh[7248], Fresh[7247], Fresh[7246], Fresh[7245], Fresh[7244], Fresh[7243], Fresh[7242], Fresh[7241], Fresh[7240]}), .outt ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, new_AGEMA_signal_3297, n1959}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2109 ( .ina ({new_AGEMA_signal_3128, new_AGEMA_signal_3127, new_AGEMA_signal_3126, n1982}), .inb ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, new_AGEMA_signal_2895, n1981}), .clk ( clk ), .rnd ({Fresh[7259], Fresh[7258], Fresh[7257], Fresh[7256], Fresh[7255], Fresh[7254], Fresh[7253], Fresh[7252], Fresh[7251], Fresh[7250]}), .outt ({new_AGEMA_signal_3302, new_AGEMA_signal_3301, new_AGEMA_signal_3300, n1983}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2149 ( .ina ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, new_AGEMA_signal_2577, n2012}), .inb ({new_AGEMA_signal_3134, new_AGEMA_signal_3133, new_AGEMA_signal_3132, n2011}), .clk ( clk ), .rnd ({Fresh[7269], Fresh[7268], Fresh[7267], Fresh[7266], Fresh[7265], Fresh[7264], Fresh[7263], Fresh[7262], Fresh[7261], Fresh[7260]}), .outt ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, new_AGEMA_signal_3303, n2014}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2166 ( .ina ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, new_AGEMA_signal_1323, n2026}), .inb ({new_AGEMA_signal_2906, new_AGEMA_signal_2905, new_AGEMA_signal_2904, n2025}), .clk ( clk ), .rnd ({Fresh[7279], Fresh[7278], Fresh[7277], Fresh[7276], Fresh[7275], Fresh[7274], Fresh[7273], Fresh[7272], Fresh[7271], Fresh[7270]}), .outt ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, new_AGEMA_signal_3135, n2029}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2180 ( .ina ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .inb ({new_AGEMA_signal_3140, new_AGEMA_signal_3139, new_AGEMA_signal_3138, n2036}), .clk ( clk ), .rnd ({Fresh[7289], Fresh[7288], Fresh[7287], Fresh[7286], Fresh[7285], Fresh[7284], Fresh[7283], Fresh[7282], Fresh[7281], Fresh[7280]}), .outt ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, new_AGEMA_signal_3309, n2037}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2197 ( .ina ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, new_AGEMA_signal_1629, n2050}), .inb ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, new_AGEMA_signal_3141, n2049}), .clk ( clk ), .rnd ({Fresh[7299], Fresh[7298], Fresh[7297], Fresh[7296], Fresh[7295], Fresh[7294], Fresh[7293], Fresh[7292], Fresh[7291], Fresh[7290]}), .outt ({new_AGEMA_signal_3314, new_AGEMA_signal_3313, new_AGEMA_signal_3312, n2052}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2219 ( .ina ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, new_AGEMA_signal_3147, n2067}), .inb ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, new_AGEMA_signal_2604, n2652}), .clk ( clk ), .rnd ({Fresh[7309], Fresh[7308], Fresh[7307], Fresh[7306], Fresh[7305], Fresh[7304], Fresh[7303], Fresh[7302], Fresh[7301], Fresh[7300]}), .outt ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, new_AGEMA_signal_3315, n2070}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2258 ( .ina ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, new_AGEMA_signal_3153, n2097}), .inb ({new_AGEMA_signal_3158, new_AGEMA_signal_3157, new_AGEMA_signal_3156, n2096}), .clk ( clk ), .rnd ({Fresh[7319], Fresh[7318], Fresh[7317], Fresh[7316], Fresh[7315], Fresh[7314], Fresh[7313], Fresh[7312], Fresh[7311], Fresh[7310]}), .outt ({new_AGEMA_signal_3320, new_AGEMA_signal_3319, new_AGEMA_signal_3318, n2098}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2287 ( .ina ({new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162, n2124}), .inb ({new_AGEMA_signal_1700, new_AGEMA_signal_1699, new_AGEMA_signal_1698, n2811}), .clk ( clk ), .rnd ({Fresh[7329], Fresh[7328], Fresh[7327], Fresh[7326], Fresh[7325], Fresh[7324], Fresh[7323], Fresh[7322], Fresh[7321], Fresh[7320]}), .outt ({new_AGEMA_signal_3326, new_AGEMA_signal_3325, new_AGEMA_signal_3324, n2125}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2311 ( .ina ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, new_AGEMA_signal_2640, n2143}), .inb ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, new_AGEMA_signal_3165, n2142}), .clk ( clk ), .rnd ({Fresh[7339], Fresh[7338], Fresh[7337], Fresh[7336], Fresh[7335], Fresh[7334], Fresh[7333], Fresh[7332], Fresh[7331], Fresh[7330]}), .outt ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, new_AGEMA_signal_3327, n2145}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2333 ( .ina ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, new_AGEMA_signal_3168, n2168}), .inb ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, new_AGEMA_signal_3171, n2167}), .clk ( clk ), .rnd ({Fresh[7349], Fresh[7348], Fresh[7347], Fresh[7346], Fresh[7345], Fresh[7344], Fresh[7343], Fresh[7342], Fresh[7341], Fresh[7340]}), .outt ({new_AGEMA_signal_3332, new_AGEMA_signal_3331, new_AGEMA_signal_3330, n2169}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2350 ( .ina ({new_AGEMA_signal_3176, new_AGEMA_signal_3175, new_AGEMA_signal_3174, n2184}), .inb ({new_AGEMA_signal_1376, new_AGEMA_signal_1375, new_AGEMA_signal_1374, n2183}), .clk ( clk ), .rnd ({Fresh[7359], Fresh[7358], Fresh[7357], Fresh[7356], Fresh[7355], Fresh[7354], Fresh[7353], Fresh[7352], Fresh[7351], Fresh[7350]}), .outt ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, new_AGEMA_signal_3333, n2185}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2365 ( .ina ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, new_AGEMA_signal_3177, n2197}), .inb ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, new_AGEMA_signal_1743, n2196}), .clk ( clk ), .rnd ({Fresh[7369], Fresh[7368], Fresh[7367], Fresh[7366], Fresh[7365], Fresh[7364], Fresh[7363], Fresh[7362], Fresh[7361], Fresh[7360]}), .outt ({new_AGEMA_signal_3338, new_AGEMA_signal_3337, new_AGEMA_signal_3336, n2198}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2396 ( .ina ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, new_AGEMA_signal_3183, n2232}), .inb ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, new_AGEMA_signal_2961, n2231}), .clk ( clk ), .rnd ({Fresh[7379], Fresh[7378], Fresh[7377], Fresh[7376], Fresh[7375], Fresh[7374], Fresh[7373], Fresh[7372], Fresh[7371], Fresh[7370]}), .outt ({new_AGEMA_signal_3344, new_AGEMA_signal_3343, new_AGEMA_signal_3342, n2312}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2404 ( .ina ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, new_AGEMA_signal_3345, n2239}), .inb ({new_AGEMA_signal_1766, new_AGEMA_signal_1765, new_AGEMA_signal_1764, n2238}), .clk ( clk ), .rnd ({Fresh[7389], Fresh[7388], Fresh[7387], Fresh[7386], Fresh[7385], Fresh[7384], Fresh[7383], Fresh[7382], Fresh[7381], Fresh[7380]}), .outt ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, new_AGEMA_signal_3459, n2258}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2415 ( .ina ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, new_AGEMA_signal_3189, n2250}), .inb ({new_AGEMA_signal_2264, new_AGEMA_signal_2263, new_AGEMA_signal_2262, n2249}), .clk ( clk ), .rnd ({Fresh[7399], Fresh[7398], Fresh[7397], Fresh[7396], Fresh[7395], Fresh[7394], Fresh[7393], Fresh[7392], Fresh[7391], Fresh[7390]}), .outt ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, new_AGEMA_signal_3348, n2251}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2440 ( .ina ({new_AGEMA_signal_2690, new_AGEMA_signal_2689, new_AGEMA_signal_2688, n2273}), .inb ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, new_AGEMA_signal_3195, n2272}), .clk ( clk ), .rnd ({Fresh[7409], Fresh[7408], Fresh[7407], Fresh[7406], Fresh[7405], Fresh[7404], Fresh[7403], Fresh[7402], Fresh[7401], Fresh[7400]}), .outt ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, new_AGEMA_signal_3351, n2274}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2469 ( .ina ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, new_AGEMA_signal_2709, n2297}), .inb ({new_AGEMA_signal_3200, new_AGEMA_signal_3199, new_AGEMA_signal_3198, n2296}), .clk ( clk ), .rnd ({Fresh[7419], Fresh[7418], Fresh[7417], Fresh[7416], Fresh[7415], Fresh[7414], Fresh[7413], Fresh[7412], Fresh[7411], Fresh[7410]}), .outt ({new_AGEMA_signal_3356, new_AGEMA_signal_3355, new_AGEMA_signal_3354, n2302}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2490 ( .ina ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, new_AGEMA_signal_3201, n2324}), .inb ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2772}), .clk ( clk ), .rnd ({Fresh[7429], Fresh[7428], Fresh[7427], Fresh[7426], Fresh[7425], Fresh[7424], Fresh[7423], Fresh[7422], Fresh[7421], Fresh[7420]}), .outt ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, new_AGEMA_signal_3357, n2339}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2503 ( .ina ({new_AGEMA_signal_3206, new_AGEMA_signal_3205, new_AGEMA_signal_3204, n2337}), .inb ({new_AGEMA_signal_2996, new_AGEMA_signal_2995, new_AGEMA_signal_2994, n2336}), .clk ( clk ), .rnd ({Fresh[7439], Fresh[7438], Fresh[7437], Fresh[7436], Fresh[7435], Fresh[7434], Fresh[7433], Fresh[7432], Fresh[7431], Fresh[7430]}), .outt ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, new_AGEMA_signal_3360, n2338}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2515 ( .ina ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, new_AGEMA_signal_3207, n2350}), .inb ({new_AGEMA_signal_1838, new_AGEMA_signal_1837, new_AGEMA_signal_1836, n2349}), .clk ( clk ), .rnd ({Fresh[7449], Fresh[7448], Fresh[7447], Fresh[7446], Fresh[7445], Fresh[7444], Fresh[7443], Fresh[7442], Fresh[7441], Fresh[7440]}), .outt ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, new_AGEMA_signal_3363, n2351}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2529 ( .ina ({new_AGEMA_signal_1424, new_AGEMA_signal_1423, new_AGEMA_signal_1422, n2363}), .inb ({new_AGEMA_signal_3212, new_AGEMA_signal_3211, new_AGEMA_signal_3210, n2362}), .clk ( clk ), .rnd ({Fresh[7459], Fresh[7458], Fresh[7457], Fresh[7456], Fresh[7455], Fresh[7454], Fresh[7453], Fresh[7452], Fresh[7451], Fresh[7450]}), .outt ({new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366, n2365}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2551 ( .ina ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003, n2389}), .inb ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .rnd ({Fresh[7469], Fresh[7468], Fresh[7467], Fresh[7466], Fresh[7465], Fresh[7464], Fresh[7463], Fresh[7462], Fresh[7461], Fresh[7460]}), .outt ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, new_AGEMA_signal_3213, n2399}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2560 ( .ina ({new_AGEMA_signal_3218, new_AGEMA_signal_3217, new_AGEMA_signal_3216, n2397}), .inb ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, new_AGEMA_signal_1869, n2396}), .clk ( clk ), .rnd ({Fresh[7479], Fresh[7478], Fresh[7477], Fresh[7476], Fresh[7475], Fresh[7474], Fresh[7473], Fresh[7472], Fresh[7471], Fresh[7470]}), .outt ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, new_AGEMA_signal_3369, n2398}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2572 ( .ina ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, new_AGEMA_signal_3009, n2411}), .inb ({new_AGEMA_signal_3014, new_AGEMA_signal_3013, new_AGEMA_signal_3012, n2410}), .clk ( clk ), .rnd ({Fresh[7489], Fresh[7488], Fresh[7487], Fresh[7486], Fresh[7485], Fresh[7484], Fresh[7483], Fresh[7482], Fresh[7481], Fresh[7480]}), .outt ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, new_AGEMA_signal_3219, n2423}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2581 ( .ina ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, new_AGEMA_signal_3015, n2421}), .inb ({new_AGEMA_signal_3020, new_AGEMA_signal_3019, new_AGEMA_signal_3018, n2420}), .clk ( clk ), .rnd ({Fresh[7499], Fresh[7498], Fresh[7497], Fresh[7496], Fresh[7495], Fresh[7494], Fresh[7493], Fresh[7492], Fresh[7491], Fresh[7490]}), .outt ({new_AGEMA_signal_3224, new_AGEMA_signal_3223, new_AGEMA_signal_3222, n2422}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2596 ( .ina ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, new_AGEMA_signal_3225, n2440}), .inb ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, new_AGEMA_signal_2367, n2439}), .clk ( clk ), .rnd ({Fresh[7509], Fresh[7508], Fresh[7507], Fresh[7506], Fresh[7505], Fresh[7504], Fresh[7503], Fresh[7502], Fresh[7501], Fresh[7500]}), .outt ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, new_AGEMA_signal_3375, n2441}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2623 ( .ina ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, new_AGEMA_signal_3033, n2471}), .inb ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, new_AGEMA_signal_1899, n2470}), .clk ( clk ), .rnd ({Fresh[7519], Fresh[7518], Fresh[7517], Fresh[7516], Fresh[7515], Fresh[7514], Fresh[7513], Fresh[7512], Fresh[7511], Fresh[7510]}), .outt ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, new_AGEMA_signal_3231, n2479}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2637 ( .ina ({new_AGEMA_signal_3236, new_AGEMA_signal_3235, new_AGEMA_signal_3234, n2485}), .inb ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .clk ( clk ), .rnd ({Fresh[7529], Fresh[7528], Fresh[7527], Fresh[7526], Fresh[7525], Fresh[7524], Fresh[7523], Fresh[7522], Fresh[7521], Fresh[7520]}), .outt ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, new_AGEMA_signal_3381, n2512}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2652 ( .ina ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, new_AGEMA_signal_3039, n2502}), .inb ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, new_AGEMA_signal_3237, n2501}), .clk ( clk ), .rnd ({Fresh[7539], Fresh[7538], Fresh[7537], Fresh[7536], Fresh[7535], Fresh[7534], Fresh[7533], Fresh[7532], Fresh[7531], Fresh[7530]}), .outt ({new_AGEMA_signal_3386, new_AGEMA_signal_3385, new_AGEMA_signal_3384, n2510}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2686 ( .ina ({new_AGEMA_signal_3248, new_AGEMA_signal_3247, new_AGEMA_signal_3246, n2550}), .inb ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, new_AGEMA_signal_3249, n2549}), .clk ( clk ), .rnd ({Fresh[7549], Fresh[7548], Fresh[7547], Fresh[7546], Fresh[7545], Fresh[7544], Fresh[7543], Fresh[7542], Fresh[7541], Fresh[7540]}), .outt ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, new_AGEMA_signal_3393, n2552}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2702 ( .ina ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2570}), .inb ({new_AGEMA_signal_3254, new_AGEMA_signal_3253, new_AGEMA_signal_3252, n2569}), .clk ( clk ), .rnd ({Fresh[7559], Fresh[7558], Fresh[7557], Fresh[7556], Fresh[7555], Fresh[7554], Fresh[7553], Fresh[7552], Fresh[7551], Fresh[7550]}), .outt ({new_AGEMA_signal_3398, new_AGEMA_signal_3397, new_AGEMA_signal_3396, n2593}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2713 ( .ina ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, new_AGEMA_signal_2439, n2585}), .inb ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, new_AGEMA_signal_3255, n2584}), .clk ( clk ), .rnd ({Fresh[7569], Fresh[7568], Fresh[7567], Fresh[7566], Fresh[7565], Fresh[7564], Fresh[7563], Fresh[7562], Fresh[7561], Fresh[7560]}), .outt ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, new_AGEMA_signal_3399, n2589}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2730 ( .ina ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, new_AGEMA_signal_1953, n2607}), .inb ({new_AGEMA_signal_3068, new_AGEMA_signal_3067, new_AGEMA_signal_3066, n2606}), .clk ( clk ), .rnd ({Fresh[7579], Fresh[7578], Fresh[7577], Fresh[7576], Fresh[7575], Fresh[7574], Fresh[7573], Fresh[7572], Fresh[7571], Fresh[7570]}), .outt ({new_AGEMA_signal_3260, new_AGEMA_signal_3259, new_AGEMA_signal_3258, n2608}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2748 ( .ina ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .inb ({new_AGEMA_signal_3266, new_AGEMA_signal_3265, new_AGEMA_signal_3264, n2634}), .clk ( clk ), .rnd ({Fresh[7589], Fresh[7588], Fresh[7587], Fresh[7586], Fresh[7585], Fresh[7584], Fresh[7583], Fresh[7582], Fresh[7581], Fresh[7580]}), .outt ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, new_AGEMA_signal_3405, n2636}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2762 ( .ina ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, new_AGEMA_signal_2550, n2658}), .inb ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, new_AGEMA_signal_3267, n2657}), .clk ( clk ), .rnd ({Fresh[7599], Fresh[7598], Fresh[7597], Fresh[7596], Fresh[7595], Fresh[7594], Fresh[7593], Fresh[7592], Fresh[7591], Fresh[7590]}), .outt ({new_AGEMA_signal_3410, new_AGEMA_signal_3409, new_AGEMA_signal_3408, n2659}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2784 ( .ina ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, new_AGEMA_signal_2835, n2698}), .inb ({new_AGEMA_signal_3272, new_AGEMA_signal_3271, new_AGEMA_signal_3270, n2697}), .clk ( clk ), .rnd ({Fresh[7609], Fresh[7608], Fresh[7607], Fresh[7606], Fresh[7605], Fresh[7604], Fresh[7603], Fresh[7602], Fresh[7601], Fresh[7600]}), .outt ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, new_AGEMA_signal_3411, n2702}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2811 ( .ina ({new_AGEMA_signal_3278, new_AGEMA_signal_3277, new_AGEMA_signal_3276, n2747}), .inb ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, new_AGEMA_signal_3279, n2746}), .clk ( clk ), .rnd ({Fresh[7619], Fresh[7618], Fresh[7617], Fresh[7616], Fresh[7615], Fresh[7614], Fresh[7613], Fresh[7612], Fresh[7611], Fresh[7610]}), .outt ({new_AGEMA_signal_3416, new_AGEMA_signal_3415, new_AGEMA_signal_3414, n2806}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2839 ( .ina ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, new_AGEMA_signal_2859, n2800}), .inb ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, new_AGEMA_signal_3111, n2799}), .clk ( clk ), .rnd ({Fresh[7629], Fresh[7628], Fresh[7627], Fresh[7626], Fresh[7625], Fresh[7624], Fresh[7623], Fresh[7622], Fresh[7621], Fresh[7620]}), .outt ({new_AGEMA_signal_3290, new_AGEMA_signal_3289, new_AGEMA_signal_3288, n2801}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2853 ( .ina ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, n2828}), .inb ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, new_AGEMA_signal_3291, n2827}), .clk ( clk ), .rnd ({Fresh[7639], Fresh[7638], Fresh[7637], Fresh[7636], Fresh[7635], Fresh[7634], Fresh[7633], Fresh[7632], Fresh[7631], Fresh[7630]}), .outt ({new_AGEMA_signal_3422, new_AGEMA_signal_3421, new_AGEMA_signal_3420, n2829}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2003 ( .ina ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, new_AGEMA_signal_2526, n1936}), .inb ({new_AGEMA_signal_3296, new_AGEMA_signal_3295, new_AGEMA_signal_3294, n1935}), .clk ( clk ), .rnd ({Fresh[7649], Fresh[7648], Fresh[7647], Fresh[7646], Fresh[7645], Fresh[7644], Fresh[7643], Fresh[7642], Fresh[7641], Fresh[7640]}), .outt ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, new_AGEMA_signal_3423, n1941}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2059 ( .ina ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, new_AGEMA_signal_3297, n1959}), .inb ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, new_AGEMA_signal_2550, n2658}), .clk ( clk ), .rnd ({Fresh[7659], Fresh[7658], Fresh[7657], Fresh[7656], Fresh[7655], Fresh[7654], Fresh[7653], Fresh[7652], Fresh[7651], Fresh[7650]}), .outt ({new_AGEMA_signal_3428, new_AGEMA_signal_3427, new_AGEMA_signal_3426, n1960}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2110 ( .ina ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, new_AGEMA_signal_3123, n1984}), .inb ({new_AGEMA_signal_3302, new_AGEMA_signal_3301, new_AGEMA_signal_3300, n1983}), .clk ( clk ), .rnd ({Fresh[7669], Fresh[7668], Fresh[7667], Fresh[7666], Fresh[7665], Fresh[7664], Fresh[7663], Fresh[7662], Fresh[7661], Fresh[7660]}), .outt ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, new_AGEMA_signal_3429, n1988}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2153 ( .ina ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, new_AGEMA_signal_3303, n2014}), .inb ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, new_AGEMA_signal_2121, n2013}), .clk ( clk ), .rnd ({Fresh[7679], Fresh[7678], Fresh[7677], Fresh[7676], Fresh[7675], Fresh[7674], Fresh[7673], Fresh[7672], Fresh[7671], Fresh[7670]}), .outt ({new_AGEMA_signal_3434, new_AGEMA_signal_3433, new_AGEMA_signal_3432, n2015}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2169 ( .ina ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, new_AGEMA_signal_3135, n2029}), .inb ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, new_AGEMA_signal_1329, n2028}), .clk ( clk ), .rnd ({Fresh[7689], Fresh[7688], Fresh[7687], Fresh[7686], Fresh[7685], Fresh[7684], Fresh[7683], Fresh[7682], Fresh[7681], Fresh[7680]}), .outt ({new_AGEMA_signal_3308, new_AGEMA_signal_3307, new_AGEMA_signal_3306, n2030}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2200 ( .ina ({new_AGEMA_signal_3314, new_AGEMA_signal_3313, new_AGEMA_signal_3312, n2052}), .inb ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, new_AGEMA_signal_2139, n2051}), .clk ( clk ), .rnd ({Fresh[7699], Fresh[7698], Fresh[7697], Fresh[7696], Fresh[7695], Fresh[7694], Fresh[7693], Fresh[7692], Fresh[7691], Fresh[7690]}), .outt ({new_AGEMA_signal_3440, new_AGEMA_signal_3439, new_AGEMA_signal_3438, n2053}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2222 ( .ina ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, new_AGEMA_signal_3315, n2070}), .inb ({new_AGEMA_signal_2156, new_AGEMA_signal_2155, new_AGEMA_signal_2154, n2069}), .clk ( clk ), .rnd ({Fresh[7709], Fresh[7708], Fresh[7707], Fresh[7706], Fresh[7705], Fresh[7704], Fresh[7703], Fresh[7702], Fresh[7701], Fresh[7700]}), .outt ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, new_AGEMA_signal_3441, n2071}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2259 ( .ina ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, new_AGEMA_signal_2613, n2099}), .inb ({new_AGEMA_signal_3320, new_AGEMA_signal_3319, new_AGEMA_signal_3318, n2098}), .clk ( clk ), .rnd ({Fresh[7719], Fresh[7718], Fresh[7717], Fresh[7716], Fresh[7715], Fresh[7714], Fresh[7713], Fresh[7712], Fresh[7711], Fresh[7710]}), .outt ({new_AGEMA_signal_3446, new_AGEMA_signal_3445, new_AGEMA_signal_3444, n2103}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2288 ( .ina ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, new_AGEMA_signal_1353, n2544}), .inb ({new_AGEMA_signal_3326, new_AGEMA_signal_3325, new_AGEMA_signal_3324, n2125}), .clk ( clk ), .rnd ({Fresh[7729], Fresh[7728], Fresh[7727], Fresh[7726], Fresh[7725], Fresh[7724], Fresh[7723], Fresh[7722], Fresh[7721], Fresh[7720]}), .outt ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, new_AGEMA_signal_3447, n2126}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2314 ( .ina ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, new_AGEMA_signal_3327, n2145}), .inb ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, new_AGEMA_signal_2205, n2144}), .clk ( clk ), .rnd ({Fresh[7739], Fresh[7738], Fresh[7737], Fresh[7736], Fresh[7735], Fresh[7734], Fresh[7733], Fresh[7732], Fresh[7731], Fresh[7730]}), .outt ({new_AGEMA_signal_3452, new_AGEMA_signal_3451, new_AGEMA_signal_3450, n2146}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2334 ( .ina ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, new_AGEMA_signal_2211, n2170}), .inb ({new_AGEMA_signal_3332, new_AGEMA_signal_3331, new_AGEMA_signal_3330, n2169}), .clk ( clk ), .rnd ({Fresh[7749], Fresh[7748], Fresh[7747], Fresh[7746], Fresh[7745], Fresh[7744], Fresh[7743], Fresh[7742], Fresh[7741], Fresh[7740]}), .outt ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, new_AGEMA_signal_3453, n2173}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2351 ( .ina ({new_AGEMA_signal_1370, new_AGEMA_signal_1369, new_AGEMA_signal_1368, n2186}), .inb ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, new_AGEMA_signal_3333, n2185}), .clk ( clk ), .rnd ({Fresh[7759], Fresh[7758], Fresh[7757], Fresh[7756], Fresh[7755], Fresh[7754], Fresh[7753], Fresh[7752], Fresh[7751], Fresh[7750]}), .outt ({new_AGEMA_signal_3458, new_AGEMA_signal_3457, new_AGEMA_signal_3456, n2187}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2416 ( .ina ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .inb ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, new_AGEMA_signal_3348, n2251}), .clk ( clk ), .rnd ({Fresh[7769], Fresh[7768], Fresh[7767], Fresh[7766], Fresh[7765], Fresh[7764], Fresh[7763], Fresh[7762], Fresh[7761], Fresh[7760]}), .outt ({new_AGEMA_signal_3464, new_AGEMA_signal_3463, new_AGEMA_signal_3462, n2256}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2441 ( .ina ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, new_AGEMA_signal_3351, n2274}), .inb ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .rnd ({Fresh[7779], Fresh[7778], Fresh[7777], Fresh[7776], Fresh[7775], Fresh[7774], Fresh[7773], Fresh[7772], Fresh[7771], Fresh[7770]}), .outt ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, new_AGEMA_signal_3465, n2275}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2474 ( .ina ({new_AGEMA_signal_3356, new_AGEMA_signal_3355, new_AGEMA_signal_3354, n2302}), .inb ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, new_AGEMA_signal_2715, n2301}), .clk ( clk ), .rnd ({Fresh[7789], Fresh[7788], Fresh[7787], Fresh[7786], Fresh[7785], Fresh[7784], Fresh[7783], Fresh[7782], Fresh[7781], Fresh[7780]}), .outt ({new_AGEMA_signal_3470, new_AGEMA_signal_3469, new_AGEMA_signal_3468, n2303}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2504 ( .ina ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, new_AGEMA_signal_3357, n2339}), .inb ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, new_AGEMA_signal_3360, n2338}), .clk ( clk ), .rnd ({Fresh[7799], Fresh[7798], Fresh[7797], Fresh[7796], Fresh[7795], Fresh[7794], Fresh[7793], Fresh[7792], Fresh[7791], Fresh[7790]}), .outt ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, new_AGEMA_signal_3471, n2382}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2516 ( .ina ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, new_AGEMA_signal_3363, n2351}), .inb ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .clk ( clk ), .rnd ({Fresh[7809], Fresh[7808], Fresh[7807], Fresh[7806], Fresh[7805], Fresh[7804], Fresh[7803], Fresh[7802], Fresh[7801], Fresh[7800]}), .outt ({new_AGEMA_signal_3476, new_AGEMA_signal_3475, new_AGEMA_signal_3474, n2380}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2531 ( .ina ({new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366, n2365}), .inb ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, new_AGEMA_signal_1851, n2364}), .clk ( clk ), .rnd ({Fresh[7819], Fresh[7818], Fresh[7817], Fresh[7816], Fresh[7815], Fresh[7814], Fresh[7813], Fresh[7812], Fresh[7811], Fresh[7810]}), .outt ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, new_AGEMA_signal_3477, n2366}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2561 ( .ina ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, new_AGEMA_signal_3213, n2399}), .inb ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, new_AGEMA_signal_3369, n2398}), .clk ( clk ), .rnd ({Fresh[7829], Fresh[7828], Fresh[7827], Fresh[7826], Fresh[7825], Fresh[7824], Fresh[7823], Fresh[7822], Fresh[7821], Fresh[7820]}), .outt ({new_AGEMA_signal_3482, new_AGEMA_signal_3481, new_AGEMA_signal_3480, n2425}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2582 ( .ina ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, new_AGEMA_signal_3219, n2423}), .inb ({new_AGEMA_signal_3224, new_AGEMA_signal_3223, new_AGEMA_signal_3222, n2422}), .clk ( clk ), .rnd ({Fresh[7839], Fresh[7838], Fresh[7837], Fresh[7836], Fresh[7835], Fresh[7834], Fresh[7833], Fresh[7832], Fresh[7831], Fresh[7830]}), .outt ({new_AGEMA_signal_3374, new_AGEMA_signal_3373, new_AGEMA_signal_3372, n2424}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2597 ( .ina ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .inb ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, new_AGEMA_signal_3375, n2441}), .clk ( clk ), .rnd ({Fresh[7849], Fresh[7848], Fresh[7847], Fresh[7846], Fresh[7845], Fresh[7844], Fresh[7843], Fresh[7842], Fresh[7841], Fresh[7840]}), .outt ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, new_AGEMA_signal_3483, n2451}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2631 ( .ina ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, new_AGEMA_signal_3231, n2479}), .inb ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, new_AGEMA_signal_2775, n2478}), .clk ( clk ), .rnd ({Fresh[7859], Fresh[7858], Fresh[7857], Fresh[7856], Fresh[7855], Fresh[7854], Fresh[7853], Fresh[7852], Fresh[7851], Fresh[7850]}), .outt ({new_AGEMA_signal_3380, new_AGEMA_signal_3379, new_AGEMA_signal_3378, n2514}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2658 ( .ina ({new_AGEMA_signal_3386, new_AGEMA_signal_3385, new_AGEMA_signal_3384, n2510}), .inb ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, new_AGEMA_signal_3387, n2509}), .clk ( clk ), .rnd ({Fresh[7869], Fresh[7868], Fresh[7867], Fresh[7866], Fresh[7865], Fresh[7864], Fresh[7863], Fresh[7862], Fresh[7861], Fresh[7860]}), .outt ({new_AGEMA_signal_3488, new_AGEMA_signal_3487, new_AGEMA_signal_3486, n2511}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2688 ( .ina ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, new_AGEMA_signal_3393, n2552}), .inb ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, new_AGEMA_signal_2421, n2551}), .clk ( clk ), .rnd ({Fresh[7879], Fresh[7878], Fresh[7877], Fresh[7876], Fresh[7875], Fresh[7874], Fresh[7873], Fresh[7872], Fresh[7871], Fresh[7870]}), .outt ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, new_AGEMA_signal_3489, n2671}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2716 ( .ina ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, new_AGEMA_signal_3399, n2589}), .inb ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, new_AGEMA_signal_2448, n2588}), .clk ( clk ), .rnd ({Fresh[7889], Fresh[7888], Fresh[7887], Fresh[7886], Fresh[7885], Fresh[7884], Fresh[7883], Fresh[7882], Fresh[7881], Fresh[7880]}), .outt ({new_AGEMA_signal_3494, new_AGEMA_signal_3493, new_AGEMA_signal_3492, n2590}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2731 ( .ina ({new_AGEMA_signal_3260, new_AGEMA_signal_3259, new_AGEMA_signal_3258, n2608}), .inb ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .clk ( clk ), .rnd ({Fresh[7899], Fresh[7898], Fresh[7897], Fresh[7896], Fresh[7895], Fresh[7894], Fresh[7893], Fresh[7892], Fresh[7891], Fresh[7890]}), .outt ({new_AGEMA_signal_3404, new_AGEMA_signal_3403, new_AGEMA_signal_3402, n2623}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2763 ( .ina ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, new_AGEMA_signal_3075, n2660}), .inb ({new_AGEMA_signal_3410, new_AGEMA_signal_3409, new_AGEMA_signal_3408, n2659}), .clk ( clk ), .rnd ({Fresh[7909], Fresh[7908], Fresh[7907], Fresh[7906], Fresh[7905], Fresh[7904], Fresh[7903], Fresh[7902], Fresh[7901], Fresh[7900]}), .outt ({new_AGEMA_signal_3500, new_AGEMA_signal_3499, new_AGEMA_signal_3498, n2667}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2786 ( .ina ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, new_AGEMA_signal_3411, n2702}), .inb ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, new_AGEMA_signal_1995, n2701}), .clk ( clk ), .rnd ({Fresh[7919], Fresh[7918], Fresh[7917], Fresh[7916], Fresh[7915], Fresh[7914], Fresh[7913], Fresh[7912], Fresh[7911], Fresh[7910]}), .outt ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, new_AGEMA_signal_3501, n2703}) ) ;
    mux2_HPC1 #(.security_order(3), .pipeline(0)) U2840 ( .ins ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .inb ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, new_AGEMA_signal_3285, n2802}), .ina ({new_AGEMA_signal_3290, new_AGEMA_signal_3289, new_AGEMA_signal_3288, n2801}), .clk ( clk ), .rnd ({Fresh[7929], Fresh[7928], Fresh[7927], Fresh[7926], Fresh[7925], Fresh[7924], Fresh[7923], Fresh[7922], Fresh[7921], Fresh[7920]}), .outt ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, new_AGEMA_signal_3417, n2803}) ) ;

    /* cells in depth 17 */

    /* cells in depth 18 */
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2016 ( .ina ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, new_AGEMA_signal_3423, n1941}), .inb ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, new_AGEMA_signal_2877, n1940}), .clk ( clk ), .rnd ({Fresh[7939], Fresh[7938], Fresh[7937], Fresh[7936], Fresh[7935], Fresh[7934], Fresh[7933], Fresh[7932], Fresh[7931], Fresh[7930]}), .outt ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, new_AGEMA_signal_3507, n2019}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2060 ( .ina ({new_AGEMA_signal_2882, new_AGEMA_signal_2881, new_AGEMA_signal_2880, n1961}), .inb ({new_AGEMA_signal_3428, new_AGEMA_signal_3427, new_AGEMA_signal_3426, n1960}), .clk ( clk ), .rnd ({Fresh[7949], Fresh[7948], Fresh[7947], Fresh[7946], Fresh[7945], Fresh[7944], Fresh[7943], Fresh[7942], Fresh[7941], Fresh[7940]}), .outt ({new_AGEMA_signal_3512, new_AGEMA_signal_3511, new_AGEMA_signal_3510, n2002}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2116 ( .ina ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, new_AGEMA_signal_3429, n1988}), .inb ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, new_AGEMA_signal_2571, n1987}), .clk ( clk ), .rnd ({Fresh[7959], Fresh[7958], Fresh[7957], Fresh[7956], Fresh[7955], Fresh[7954], Fresh[7953], Fresh[7952], Fresh[7951], Fresh[7950]}), .outt ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, new_AGEMA_signal_3513, n1989}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2154 ( .ina ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, n2828}), .inb ({new_AGEMA_signal_3434, new_AGEMA_signal_3433, new_AGEMA_signal_3432, n2015}), .clk ( clk ), .rnd ({Fresh[7969], Fresh[7968], Fresh[7967], Fresh[7966], Fresh[7965], Fresh[7964], Fresh[7963], Fresh[7962], Fresh[7961], Fresh[7960]}), .outt ({new_AGEMA_signal_3518, new_AGEMA_signal_3517, new_AGEMA_signal_3516, n2016}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2170 ( .ina ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .inb ({new_AGEMA_signal_3308, new_AGEMA_signal_3307, new_AGEMA_signal_3306, n2030}), .clk ( clk ), .rnd ({Fresh[7979], Fresh[7978], Fresh[7977], Fresh[7976], Fresh[7975], Fresh[7974], Fresh[7973], Fresh[7972], Fresh[7971], Fresh[7970]}), .outt ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, new_AGEMA_signal_3435, n2038}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2201 ( .ina ({new_AGEMA_signal_2912, new_AGEMA_signal_2911, new_AGEMA_signal_2910, n2054}), .inb ({new_AGEMA_signal_3440, new_AGEMA_signal_3439, new_AGEMA_signal_3438, n2053}), .clk ( clk ), .rnd ({Fresh[7989], Fresh[7988], Fresh[7987], Fresh[7986], Fresh[7985], Fresh[7984], Fresh[7983], Fresh[7982], Fresh[7981], Fresh[7980]}), .outt ({new_AGEMA_signal_3524, new_AGEMA_signal_3523, new_AGEMA_signal_3522, n2111}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2223 ( .ina ({new_AGEMA_signal_3146, new_AGEMA_signal_3145, new_AGEMA_signal_3144, n2072}), .inb ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, new_AGEMA_signal_3441, n2071}), .clk ( clk ), .rnd ({Fresh[7999], Fresh[7998], Fresh[7997], Fresh[7996], Fresh[7995], Fresh[7994], Fresh[7993], Fresh[7992], Fresh[7991], Fresh[7990]}), .outt ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, new_AGEMA_signal_3525, n2079}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2263 ( .ina ({new_AGEMA_signal_3446, new_AGEMA_signal_3445, new_AGEMA_signal_3444, n2103}), .inb ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, new_AGEMA_signal_2625, n2102}), .clk ( clk ), .rnd ({Fresh[8009], Fresh[8008], Fresh[8007], Fresh[8006], Fresh[8005], Fresh[8004], Fresh[8003], Fresh[8002], Fresh[8001], Fresh[8000]}), .outt ({new_AGEMA_signal_3530, new_AGEMA_signal_3529, new_AGEMA_signal_3528, n2104}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2289 ( .ina ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .inb ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, new_AGEMA_signal_3447, n2126}), .clk ( clk ), .rnd ({Fresh[8019], Fresh[8018], Fresh[8017], Fresh[8016], Fresh[8015], Fresh[8014], Fresh[8013], Fresh[8012], Fresh[8011], Fresh[8010]}), .outt ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, new_AGEMA_signal_3531, n2127}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2315 ( .ina ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, n2828}), .inb ({new_AGEMA_signal_3452, new_AGEMA_signal_3451, new_AGEMA_signal_3450, n2146}), .clk ( clk ), .rnd ({Fresh[8029], Fresh[8028], Fresh[8027], Fresh[8026], Fresh[8025], Fresh[8024], Fresh[8023], Fresh[8022], Fresh[8021], Fresh[8020]}), .outt ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, new_AGEMA_signal_3534, n2147}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2336 ( .ina ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, new_AGEMA_signal_3453, n2173}), .inb ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, new_AGEMA_signal_2220, n2172}), .clk ( clk ), .rnd ({Fresh[8039], Fresh[8038], Fresh[8037], Fresh[8036], Fresh[8035], Fresh[8034], Fresh[8033], Fresh[8032], Fresh[8031], Fresh[8030]}), .outt ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, new_AGEMA_signal_3537, n2208}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2352 ( .ina ({new_AGEMA_signal_3458, new_AGEMA_signal_3457, new_AGEMA_signal_3456, n2187}), .inb ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .rnd ({Fresh[8049], Fresh[8048], Fresh[8047], Fresh[8046], Fresh[8045], Fresh[8044], Fresh[8043], Fresh[8042], Fresh[8041], Fresh[8040]}), .outt ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, new_AGEMA_signal_3540, n2199}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2420 ( .ina ({new_AGEMA_signal_3464, new_AGEMA_signal_3463, new_AGEMA_signal_3462, n2256}), .inb ({new_AGEMA_signal_2972, new_AGEMA_signal_2971, new_AGEMA_signal_2970, n2255}), .clk ( clk ), .rnd ({Fresh[8059], Fresh[8058], Fresh[8057], Fresh[8056], Fresh[8055], Fresh[8054], Fresh[8053], Fresh[8052], Fresh[8051], Fresh[8050]}), .outt ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, new_AGEMA_signal_3543, n2257}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2442 ( .ina ({new_AGEMA_signal_3194, new_AGEMA_signal_3193, new_AGEMA_signal_3192, n2276}), .inb ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, new_AGEMA_signal_3465, n2275}), .clk ( clk ), .rnd ({Fresh[8069], Fresh[8068], Fresh[8067], Fresh[8066], Fresh[8065], Fresh[8064], Fresh[8063], Fresh[8062], Fresh[8061], Fresh[8060]}), .outt ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, new_AGEMA_signal_3546, n2281}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2475 ( .ina ({new_AGEMA_signal_2984, new_AGEMA_signal_2983, new_AGEMA_signal_2982, n2304}), .inb ({new_AGEMA_signal_3470, new_AGEMA_signal_3469, new_AGEMA_signal_3468, n2303}), .clk ( clk ), .rnd ({Fresh[8079], Fresh[8078], Fresh[8077], Fresh[8076], Fresh[8075], Fresh[8074], Fresh[8073], Fresh[8072], Fresh[8071], Fresh[8070]}), .outt ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, new_AGEMA_signal_3549, n2305}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2532 ( .ina ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, new_AGEMA_signal_2316, n2367}), .inb ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, new_AGEMA_signal_3477, n2366}), .clk ( clk ), .rnd ({Fresh[8089], Fresh[8088], Fresh[8087], Fresh[8086], Fresh[8085], Fresh[8084], Fresh[8083], Fresh[8082], Fresh[8081], Fresh[8080]}), .outt ({new_AGEMA_signal_3554, new_AGEMA_signal_3553, new_AGEMA_signal_3552, n2368}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2583 ( .ina ({new_AGEMA_signal_3482, new_AGEMA_signal_3481, new_AGEMA_signal_3480, n2425}), .inb ({new_AGEMA_signal_3374, new_AGEMA_signal_3373, new_AGEMA_signal_3372, n2424}), .clk ( clk ), .rnd ({Fresh[8099], Fresh[8098], Fresh[8097], Fresh[8096], Fresh[8095], Fresh[8094], Fresh[8093], Fresh[8092], Fresh[8091], Fresh[8090]}), .outt ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, new_AGEMA_signal_3555, n2426}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2605 ( .ina ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, new_AGEMA_signal_3483, n2451}), .inb ({new_AGEMA_signal_3026, new_AGEMA_signal_3025, new_AGEMA_signal_3024, n2450}), .clk ( clk ), .rnd ({Fresh[8109], Fresh[8108], Fresh[8107], Fresh[8106], Fresh[8105], Fresh[8104], Fresh[8103], Fresh[8102], Fresh[8101], Fresh[8100]}), .outt ({new_AGEMA_signal_3560, new_AGEMA_signal_3559, new_AGEMA_signal_3558, n2457}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2659 ( .ina ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, new_AGEMA_signal_3381, n2512}), .inb ({new_AGEMA_signal_3488, new_AGEMA_signal_3487, new_AGEMA_signal_3486, n2511}), .clk ( clk ), .rnd ({Fresh[8119], Fresh[8118], Fresh[8117], Fresh[8116], Fresh[8115], Fresh[8114], Fresh[8113], Fresh[8112], Fresh[8111], Fresh[8110]}), .outt ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, new_AGEMA_signal_3561, n2513}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2717 ( .ina ({new_AGEMA_signal_2810, new_AGEMA_signal_2809, new_AGEMA_signal_2808, n2591}), .inb ({new_AGEMA_signal_3494, new_AGEMA_signal_3493, new_AGEMA_signal_3492, n2590}), .clk ( clk ), .rnd ({Fresh[8129], Fresh[8128], Fresh[8127], Fresh[8126], Fresh[8125], Fresh[8124], Fresh[8123], Fresh[8122], Fresh[8121], Fresh[8120]}), .outt ({new_AGEMA_signal_3566, new_AGEMA_signal_3565, new_AGEMA_signal_3564, n2592}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2741 ( .ina ({new_AGEMA_signal_3404, new_AGEMA_signal_3403, new_AGEMA_signal_3402, n2623}), .inb ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, new_AGEMA_signal_3261, n2622}), .clk ( clk ), .rnd ({Fresh[8139], Fresh[8138], Fresh[8137], Fresh[8136], Fresh[8135], Fresh[8134], Fresh[8133], Fresh[8132], Fresh[8131], Fresh[8130]}), .outt ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, new_AGEMA_signal_3495, n2637}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2767 ( .ina ({new_AGEMA_signal_3500, new_AGEMA_signal_3499, new_AGEMA_signal_3498, n2667}), .inb ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, new_AGEMA_signal_3081, n2666}), .clk ( clk ), .rnd ({Fresh[8149], Fresh[8148], Fresh[8147], Fresh[8146], Fresh[8145], Fresh[8144], Fresh[8143], Fresh[8142], Fresh[8141], Fresh[8140]}), .outt ({new_AGEMA_signal_3572, new_AGEMA_signal_3571, new_AGEMA_signal_3570, n2668}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2787 ( .ina ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, new_AGEMA_signal_3087, n2704}), .inb ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, new_AGEMA_signal_3501, n2703}), .clk ( clk ), .rnd ({Fresh[8159], Fresh[8158], Fresh[8157], Fresh[8156], Fresh[8155], Fresh[8154], Fresh[8153], Fresh[8152], Fresh[8151], Fresh[8150]}), .outt ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, new_AGEMA_signal_3573, n2705}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2841 ( .ina ({new_AGEMA_signal_3284, new_AGEMA_signal_3283, new_AGEMA_signal_3282, n2804}), .inb ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, new_AGEMA_signal_3417, n2803}), .clk ( clk ), .rnd ({Fresh[8169], Fresh[8168], Fresh[8167], Fresh[8166], Fresh[8165], Fresh[8164], Fresh[8163], Fresh[8162], Fresh[8161], Fresh[8160]}), .outt ({new_AGEMA_signal_3506, new_AGEMA_signal_3505, new_AGEMA_signal_3504, n2805}) ) ;

    /* cells in depth 19 */

    /* cells in depth 20 */
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2117 ( .ina ({new_AGEMA_signal_2888, new_AGEMA_signal_2887, new_AGEMA_signal_2886, n1990}), .inb ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, new_AGEMA_signal_3513, n1989}), .clk ( clk ), .rnd ({Fresh[8179], Fresh[8178], Fresh[8177], Fresh[8176], Fresh[8175], Fresh[8174], Fresh[8173], Fresh[8172], Fresh[8171], Fresh[8170]}), .outt ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, new_AGEMA_signal_3579, n2000}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2181 ( .ina ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, new_AGEMA_signal_3435, n2038}), .inb ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, new_AGEMA_signal_3309, n2037}), .clk ( clk ), .rnd ({Fresh[8189], Fresh[8188], Fresh[8187], Fresh[8186], Fresh[8185], Fresh[8184], Fresh[8183], Fresh[8182], Fresh[8181], Fresh[8180]}), .outt ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, new_AGEMA_signal_3519, n2113}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2231 ( .ina ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, new_AGEMA_signal_3525, n2079}), .inb ({new_AGEMA_signal_3152, new_AGEMA_signal_3151, new_AGEMA_signal_3150, n2078}), .clk ( clk ), .rnd ({Fresh[8199], Fresh[8198], Fresh[8197], Fresh[8196], Fresh[8195], Fresh[8194], Fresh[8193], Fresh[8192], Fresh[8191], Fresh[8190]}), .outt ({new_AGEMA_signal_3584, new_AGEMA_signal_3583, new_AGEMA_signal_3582, n2109}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2264 ( .ina ({new_AGEMA_signal_2612, new_AGEMA_signal_2611, new_AGEMA_signal_2610, n2105}), .inb ({new_AGEMA_signal_3530, new_AGEMA_signal_3529, new_AGEMA_signal_3528, n2104}), .clk ( clk ), .rnd ({Fresh[8209], Fresh[8208], Fresh[8207], Fresh[8206], Fresh[8205], Fresh[8204], Fresh[8203], Fresh[8202], Fresh[8201], Fresh[8200]}), .outt ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, new_AGEMA_signal_3585, n2107}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2290 ( .ina ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, new_AGEMA_signal_3321, n2128}), .inb ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, new_AGEMA_signal_3531, n2127}), .clk ( clk ), .rnd ({Fresh[8219], Fresh[8218], Fresh[8217], Fresh[8216], Fresh[8215], Fresh[8214], Fresh[8213], Fresh[8212], Fresh[8211], Fresh[8210]}), .outt ({new_AGEMA_signal_3590, new_AGEMA_signal_3589, new_AGEMA_signal_3588, n2212}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2316 ( .ina ({new_AGEMA_signal_2942, new_AGEMA_signal_2941, new_AGEMA_signal_2940, n2148}), .inb ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, new_AGEMA_signal_3534, n2147}), .clk ( clk ), .rnd ({Fresh[8229], Fresh[8228], Fresh[8227], Fresh[8226], Fresh[8225], Fresh[8224], Fresh[8223], Fresh[8222], Fresh[8221], Fresh[8220]}), .outt ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, new_AGEMA_signal_3591, n2149}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2366 ( .ina ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, new_AGEMA_signal_3540, n2199}), .inb ({new_AGEMA_signal_3338, new_AGEMA_signal_3337, new_AGEMA_signal_3336, n2198}), .clk ( clk ), .rnd ({Fresh[8239], Fresh[8238], Fresh[8237], Fresh[8236], Fresh[8235], Fresh[8234], Fresh[8233], Fresh[8232], Fresh[8231], Fresh[8230]}), .outt ({new_AGEMA_signal_3596, new_AGEMA_signal_3595, new_AGEMA_signal_3594, n2206}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2421 ( .ina ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, new_AGEMA_signal_3459, n2258}), .inb ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, new_AGEMA_signal_3543, n2257}), .clk ( clk ), .rnd ({Fresh[8249], Fresh[8248], Fresh[8247], Fresh[8246], Fresh[8245], Fresh[8244], Fresh[8243], Fresh[8242], Fresh[8241], Fresh[8240]}), .outt ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, new_AGEMA_signal_3597, n2310}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2447 ( .ina ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, new_AGEMA_signal_3546, n2281}), .inb ({new_AGEMA_signal_2696, new_AGEMA_signal_2695, new_AGEMA_signal_2694, n2280}), .clk ( clk ), .rnd ({Fresh[8259], Fresh[8258], Fresh[8257], Fresh[8256], Fresh[8255], Fresh[8254], Fresh[8253], Fresh[8252], Fresh[8251], Fresh[8250]}), .outt ({new_AGEMA_signal_3602, new_AGEMA_signal_3601, new_AGEMA_signal_3600, n2308}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2476 ( .ina ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, new_AGEMA_signal_2979, n2306}), .inb ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, new_AGEMA_signal_3549, n2305}), .clk ( clk ), .rnd ({Fresh[8269], Fresh[8268], Fresh[8267], Fresh[8266], Fresh[8265], Fresh[8264], Fresh[8263], Fresh[8262], Fresh[8261], Fresh[8260]}), .outt ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, new_AGEMA_signal_3603, n2307}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2533 ( .ina ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .inb ({new_AGEMA_signal_3554, new_AGEMA_signal_3553, new_AGEMA_signal_3552, n2368}), .clk ( clk ), .rnd ({Fresh[8279], Fresh[8278], Fresh[8277], Fresh[8276], Fresh[8275], Fresh[8274], Fresh[8273], Fresh[8272], Fresh[8271], Fresh[8270]}), .outt ({new_AGEMA_signal_3608, new_AGEMA_signal_3607, new_AGEMA_signal_3606, n2370}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2611 ( .ina ({new_AGEMA_signal_3560, new_AGEMA_signal_3559, new_AGEMA_signal_3558, n2457}), .inb ({new_AGEMA_signal_3029, new_AGEMA_signal_3028, new_AGEMA_signal_3027, n2456}), .clk ( clk ), .rnd ({Fresh[8289], Fresh[8288], Fresh[8287], Fresh[8286], Fresh[8285], Fresh[8284], Fresh[8283], Fresh[8282], Fresh[8281], Fresh[8280]}), .outt ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, new_AGEMA_signal_3609, n2530}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2660 ( .ina ({new_AGEMA_signal_3380, new_AGEMA_signal_3379, new_AGEMA_signal_3378, n2514}), .inb ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, new_AGEMA_signal_3561, n2513}), .clk ( clk ), .rnd ({Fresh[8299], Fresh[8298], Fresh[8297], Fresh[8296], Fresh[8295], Fresh[8294], Fresh[8293], Fresh[8292], Fresh[8291], Fresh[8290]}), .outt ({new_AGEMA_signal_3614, new_AGEMA_signal_3613, new_AGEMA_signal_3612, n2515}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2718 ( .ina ({new_AGEMA_signal_3398, new_AGEMA_signal_3397, new_AGEMA_signal_3396, n2593}), .inb ({new_AGEMA_signal_3566, new_AGEMA_signal_3565, new_AGEMA_signal_3564, n2592}), .clk ( clk ), .rnd ({Fresh[8309], Fresh[8308], Fresh[8307], Fresh[8306], Fresh[8305], Fresh[8304], Fresh[8303], Fresh[8302], Fresh[8301], Fresh[8300]}), .outt ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, new_AGEMA_signal_3615, n2639}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2749 ( .ina ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, new_AGEMA_signal_3495, n2637}), .inb ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, new_AGEMA_signal_3405, n2636}), .clk ( clk ), .rnd ({Fresh[8319], Fresh[8318], Fresh[8317], Fresh[8316], Fresh[8315], Fresh[8314], Fresh[8313], Fresh[8312], Fresh[8311], Fresh[8310]}), .outt ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, new_AGEMA_signal_3567, n2638}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2788 ( .ina ({new_AGEMA_signal_3086, new_AGEMA_signal_3085, new_AGEMA_signal_3084, n2706}), .inb ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, new_AGEMA_signal_3573, n2705}), .clk ( clk ), .rnd ({Fresh[8329], Fresh[8328], Fresh[8327], Fresh[8326], Fresh[8325], Fresh[8324], Fresh[8323], Fresh[8322], Fresh[8321], Fresh[8320]}), .outt ({new_AGEMA_signal_3620, new_AGEMA_signal_3619, new_AGEMA_signal_3618, n2832}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2842 ( .ina ({new_AGEMA_signal_3416, new_AGEMA_signal_3415, new_AGEMA_signal_3414, n2806}), .inb ({new_AGEMA_signal_3506, new_AGEMA_signal_3505, new_AGEMA_signal_3504, n2805}), .clk ( clk ), .rnd ({Fresh[8339], Fresh[8338], Fresh[8337], Fresh[8336], Fresh[8335], Fresh[8334], Fresh[8333], Fresh[8332], Fresh[8331], Fresh[8330]}), .outt ({new_AGEMA_signal_3578, new_AGEMA_signal_3577, new_AGEMA_signal_3576, n2807}) ) ;

    /* cells in depth 21 */

    /* cells in depth 22 */
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2129 ( .ina ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, new_AGEMA_signal_3579, n2000}), .inb ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, new_AGEMA_signal_3129, n1999}), .clk ( clk ), .rnd ({Fresh[8349], Fresh[8348], Fresh[8347], Fresh[8346], Fresh[8345], Fresh[8344], Fresh[8343], Fresh[8342], Fresh[8341], Fresh[8340]}), .outt ({new_AGEMA_signal_3626, new_AGEMA_signal_3625, new_AGEMA_signal_3624, n2001}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2267 ( .ina ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, new_AGEMA_signal_3585, n2107}), .inb ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, new_AGEMA_signal_2187, n2106}), .clk ( clk ), .rnd ({Fresh[8359], Fresh[8358], Fresh[8357], Fresh[8356], Fresh[8355], Fresh[8354], Fresh[8353], Fresh[8352], Fresh[8351], Fresh[8350]}), .outt ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, new_AGEMA_signal_3627, n2108}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2317 ( .ina ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, new_AGEMA_signal_1707, n2150}), .inb ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, new_AGEMA_signal_3591, n2149}), .clk ( clk ), .rnd ({Fresh[8369], Fresh[8368], Fresh[8367], Fresh[8366], Fresh[8365], Fresh[8364], Fresh[8363], Fresh[8362], Fresh[8361], Fresh[8360]}), .outt ({new_AGEMA_signal_3632, new_AGEMA_signal_3631, new_AGEMA_signal_3630, n2153}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2374 ( .ina ({new_AGEMA_signal_3596, new_AGEMA_signal_3595, new_AGEMA_signal_3594, n2206}), .inb ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, new_AGEMA_signal_3339, n2205}), .clk ( clk ), .rnd ({Fresh[8379], Fresh[8378], Fresh[8377], Fresh[8376], Fresh[8375], Fresh[8374], Fresh[8373], Fresh[8372], Fresh[8371], Fresh[8370]}), .outt ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, new_AGEMA_signal_3633, n2207}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2477 ( .ina ({new_AGEMA_signal_3602, new_AGEMA_signal_3601, new_AGEMA_signal_3600, n2308}), .inb ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, new_AGEMA_signal_3603, n2307}), .clk ( clk ), .rnd ({Fresh[8389], Fresh[8388], Fresh[8387], Fresh[8386], Fresh[8385], Fresh[8384], Fresh[8383], Fresh[8382], Fresh[8381], Fresh[8380]}), .outt ({new_AGEMA_signal_3638, new_AGEMA_signal_3637, new_AGEMA_signal_3636, n2309}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2535 ( .ina ({new_AGEMA_signal_3608, new_AGEMA_signal_3607, new_AGEMA_signal_3606, n2370}), .inb ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, new_AGEMA_signal_2736, n2369}), .clk ( clk ), .rnd ({Fresh[8399], Fresh[8398], Fresh[8397], Fresh[8396], Fresh[8395], Fresh[8394], Fresh[8393], Fresh[8392], Fresh[8391], Fresh[8390]}), .outt ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, new_AGEMA_signal_3639, n2373}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2661 ( .ina ({new_AGEMA_signal_3230, new_AGEMA_signal_3229, new_AGEMA_signal_3228, n2516}), .inb ({new_AGEMA_signal_3614, new_AGEMA_signal_3613, new_AGEMA_signal_3612, n2515}), .clk ( clk ), .rnd ({Fresh[8409], Fresh[8408], Fresh[8407], Fresh[8406], Fresh[8405], Fresh[8404], Fresh[8403], Fresh[8402], Fresh[8401], Fresh[8400]}), .outt ({new_AGEMA_signal_3644, new_AGEMA_signal_3643, new_AGEMA_signal_3642, n2528}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2750 ( .ina ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, new_AGEMA_signal_3615, n2639}), .inb ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, new_AGEMA_signal_3567, n2638}), .clk ( clk ), .rnd ({Fresh[8419], Fresh[8418], Fresh[8417], Fresh[8416], Fresh[8415], Fresh[8414], Fresh[8413], Fresh[8412], Fresh[8411], Fresh[8410]}), .outt ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, new_AGEMA_signal_3645, n2669}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2843 ( .ina ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, new_AGEMA_signal_3273, n2808}), .inb ({new_AGEMA_signal_3578, new_AGEMA_signal_3577, new_AGEMA_signal_3576, n2807}), .clk ( clk ), .rnd ({Fresh[8429], Fresh[8428], Fresh[8427], Fresh[8426], Fresh[8425], Fresh[8424], Fresh[8423], Fresh[8422], Fresh[8421], Fresh[8420]}), .outt ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, new_AGEMA_signal_3621, n2830}) ) ;

    /* cells in depth 23 */

    /* cells in depth 24 */
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2130 ( .ina ({new_AGEMA_signal_3512, new_AGEMA_signal_3511, new_AGEMA_signal_3510, n2002}), .inb ({new_AGEMA_signal_3626, new_AGEMA_signal_3625, new_AGEMA_signal_3624, n2001}), .clk ( clk ), .rnd ({Fresh[8439], Fresh[8438], Fresh[8437], Fresh[8436], Fresh[8435], Fresh[8434], Fresh[8433], Fresh[8432], Fresh[8431], Fresh[8430]}), .outt ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, new_AGEMA_signal_3651, n2017}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2268 ( .ina ({new_AGEMA_signal_3584, new_AGEMA_signal_3583, new_AGEMA_signal_3582, n2109}), .inb ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, new_AGEMA_signal_3627, n2108}), .clk ( clk ), .rnd ({Fresh[8449], Fresh[8448], Fresh[8447], Fresh[8446], Fresh[8445], Fresh[8444], Fresh[8443], Fresh[8442], Fresh[8441], Fresh[8440]}), .outt ({new_AGEMA_signal_3656, new_AGEMA_signal_3655, new_AGEMA_signal_3654, n2110}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2319 ( .ina ({new_AGEMA_signal_3632, new_AGEMA_signal_3631, new_AGEMA_signal_3630, n2153}), .inb ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, new_AGEMA_signal_2208, n2152}), .clk ( clk ), .rnd ({Fresh[8459], Fresh[8458], Fresh[8457], Fresh[8456], Fresh[8455], Fresh[8454], Fresh[8453], Fresh[8452], Fresh[8451], Fresh[8450]}), .outt ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, new_AGEMA_signal_3657, n2154}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2375 ( .ina ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, new_AGEMA_signal_3537, n2208}), .inb ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, new_AGEMA_signal_3633, n2207}), .clk ( clk ), .rnd ({Fresh[8469], Fresh[8468], Fresh[8467], Fresh[8466], Fresh[8465], Fresh[8464], Fresh[8463], Fresh[8462], Fresh[8461], Fresh[8460]}), .outt ({new_AGEMA_signal_3662, new_AGEMA_signal_3661, new_AGEMA_signal_3660, n2209}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2478 ( .ina ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, new_AGEMA_signal_3597, n2310}), .inb ({new_AGEMA_signal_3638, new_AGEMA_signal_3637, new_AGEMA_signal_3636, n2309}), .clk ( clk ), .rnd ({Fresh[8479], Fresh[8478], Fresh[8477], Fresh[8476], Fresh[8475], Fresh[8474], Fresh[8473], Fresh[8472], Fresh[8471], Fresh[8470]}), .outt ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, new_AGEMA_signal_3663, n2311}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2537 ( .ina ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, new_AGEMA_signal_3639, n2373}), .inb ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, new_AGEMA_signal_2328, n2372}), .clk ( clk ), .rnd ({Fresh[8489], Fresh[8488], Fresh[8487], Fresh[8486], Fresh[8485], Fresh[8484], Fresh[8483], Fresh[8482], Fresh[8481], Fresh[8480]}), .outt ({new_AGEMA_signal_3668, new_AGEMA_signal_3667, new_AGEMA_signal_3666, n2374}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2672 ( .ina ({new_AGEMA_signal_3644, new_AGEMA_signal_3643, new_AGEMA_signal_3642, n2528}), .inb ({new_AGEMA_signal_3392, new_AGEMA_signal_3391, new_AGEMA_signal_3390, n2527}), .clk ( clk ), .rnd ({Fresh[8499], Fresh[8498], Fresh[8497], Fresh[8496], Fresh[8495], Fresh[8494], Fresh[8493], Fresh[8492], Fresh[8491], Fresh[8490]}), .outt ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, new_AGEMA_signal_3669, n2529}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2768 ( .ina ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, new_AGEMA_signal_3645, n2669}), .inb ({new_AGEMA_signal_3572, new_AGEMA_signal_3571, new_AGEMA_signal_3570, n2668}), .clk ( clk ), .rnd ({Fresh[8509], Fresh[8508], Fresh[8507], Fresh[8506], Fresh[8505], Fresh[8504], Fresh[8503], Fresh[8502], Fresh[8501], Fresh[8500]}), .outt ({new_AGEMA_signal_3674, new_AGEMA_signal_3673, new_AGEMA_signal_3672, n2670}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2854 ( .ina ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, new_AGEMA_signal_3621, n2830}), .inb ({new_AGEMA_signal_3422, new_AGEMA_signal_3421, new_AGEMA_signal_3420, n2829}), .clk ( clk ), .rnd ({Fresh[8519], Fresh[8518], Fresh[8517], Fresh[8516], Fresh[8515], Fresh[8514], Fresh[8513], Fresh[8512], Fresh[8511], Fresh[8510]}), .outt ({new_AGEMA_signal_3650, new_AGEMA_signal_3649, new_AGEMA_signal_3648, n2831}) ) ;

    /* cells in depth 25 */

    /* cells in depth 26 */
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2155 ( .ina ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, new_AGEMA_signal_3651, n2017}), .inb ({new_AGEMA_signal_3518, new_AGEMA_signal_3517, new_AGEMA_signal_3516, n2016}), .clk ( clk ), .rnd ({Fresh[8529], Fresh[8528], Fresh[8527], Fresh[8526], Fresh[8525], Fresh[8524], Fresh[8523], Fresh[8522], Fresh[8521], Fresh[8520]}), .outt ({new_AGEMA_signal_3680, new_AGEMA_signal_3679, new_AGEMA_signal_3678, n2018}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2269 ( .ina ({new_AGEMA_signal_3524, new_AGEMA_signal_3523, new_AGEMA_signal_3522, n2111}), .inb ({new_AGEMA_signal_3656, new_AGEMA_signal_3655, new_AGEMA_signal_3654, n2110}), .clk ( clk ), .rnd ({Fresh[8539], Fresh[8538], Fresh[8537], Fresh[8536], Fresh[8535], Fresh[8534], Fresh[8533], Fresh[8532], Fresh[8531], Fresh[8530]}), .outt ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, new_AGEMA_signal_3681, n2112}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2320 ( .ina ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, new_AGEMA_signal_2193, n2155}), .inb ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, new_AGEMA_signal_3657, n2154}), .clk ( clk ), .rnd ({Fresh[8549], Fresh[8548], Fresh[8547], Fresh[8546], Fresh[8545], Fresh[8544], Fresh[8543], Fresh[8542], Fresh[8541], Fresh[8540]}), .outt ({new_AGEMA_signal_3686, new_AGEMA_signal_3685, new_AGEMA_signal_3684, n2210}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2479 ( .ina ({new_AGEMA_signal_3344, new_AGEMA_signal_3343, new_AGEMA_signal_3342, n2312}), .inb ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, new_AGEMA_signal_3663, n2311}), .clk ( clk ), .rnd ({Fresh[8559], Fresh[8558], Fresh[8557], Fresh[8556], Fresh[8555], Fresh[8554], Fresh[8553], Fresh[8552], Fresh[8551], Fresh[8550]}), .outt ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, new_AGEMA_signal_3687, N470}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2538 ( .ina ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, new_AGEMA_signal_1839, n2375}), .inb ({new_AGEMA_signal_3668, new_AGEMA_signal_3667, new_AGEMA_signal_3666, n2374}), .clk ( clk ), .rnd ({Fresh[8569], Fresh[8568], Fresh[8567], Fresh[8566], Fresh[8565], Fresh[8564], Fresh[8563], Fresh[8562], Fresh[8561], Fresh[8560]}), .outt ({new_AGEMA_signal_3692, new_AGEMA_signal_3691, new_AGEMA_signal_3690, n2378}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2673 ( .ina ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, new_AGEMA_signal_3609, n2530}), .inb ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, new_AGEMA_signal_3669, n2529}), .clk ( clk ), .rnd ({Fresh[8579], Fresh[8578], Fresh[8577], Fresh[8576], Fresh[8575], Fresh[8574], Fresh[8573], Fresh[8572], Fresh[8571], Fresh[8570]}), .outt ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, new_AGEMA_signal_3693, N639}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2769 ( .ina ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, new_AGEMA_signal_3489, n2671}), .inb ({new_AGEMA_signal_3674, new_AGEMA_signal_3673, new_AGEMA_signal_3672, n2670}), .clk ( clk ), .rnd ({Fresh[8589], Fresh[8588], Fresh[8587], Fresh[8586], Fresh[8585], Fresh[8584], Fresh[8583], Fresh[8582], Fresh[8581], Fresh[8580]}), .outt ({new_AGEMA_signal_3698, new_AGEMA_signal_3697, new_AGEMA_signal_3696, N723}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2855 ( .ina ({new_AGEMA_signal_3620, new_AGEMA_signal_3619, new_AGEMA_signal_3618, n2832}), .inb ({new_AGEMA_signal_3650, new_AGEMA_signal_3649, new_AGEMA_signal_3648, n2831}), .clk ( clk ), .rnd ({Fresh[8599], Fresh[8598], Fresh[8597], Fresh[8596], Fresh[8595], Fresh[8594], Fresh[8593], Fresh[8592], Fresh[8591], Fresh[8590]}), .outt ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, new_AGEMA_signal_3675, N789}) ) ;

    /* cells in depth 27 */

    /* cells in depth 28 */
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2156 ( .ina ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, new_AGEMA_signal_3507, n2019}), .inb ({new_AGEMA_signal_3680, new_AGEMA_signal_3679, new_AGEMA_signal_3678, n2018}), .clk ( clk ), .rnd ({Fresh[8609], Fresh[8608], Fresh[8607], Fresh[8606], Fresh[8605], Fresh[8604], Fresh[8603], Fresh[8602], Fresh[8601], Fresh[8600]}), .outt ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, new_AGEMA_signal_3699, N169}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2270 ( .ina ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, new_AGEMA_signal_3519, n2113}), .inb ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, new_AGEMA_signal_3681, n2112}), .clk ( clk ), .rnd ({Fresh[8619], Fresh[8618], Fresh[8617], Fresh[8616], Fresh[8615], Fresh[8614], Fresh[8613], Fresh[8612], Fresh[8611], Fresh[8610]}), .outt ({new_AGEMA_signal_3704, new_AGEMA_signal_3703, new_AGEMA_signal_3702, N277}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2376 ( .ina ({new_AGEMA_signal_3686, new_AGEMA_signal_3685, new_AGEMA_signal_3684, n2210}), .inb ({new_AGEMA_signal_3662, new_AGEMA_signal_3661, new_AGEMA_signal_3660, n2209}), .clk ( clk ), .rnd ({Fresh[8629], Fresh[8628], Fresh[8627], Fresh[8626], Fresh[8625], Fresh[8624], Fresh[8623], Fresh[8622], Fresh[8621], Fresh[8620]}), .outt ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, new_AGEMA_signal_3705, n2211}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2540 ( .ina ({new_AGEMA_signal_3692, new_AGEMA_signal_3691, new_AGEMA_signal_3690, n2378}), .inb ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, new_AGEMA_signal_2331, n2377}), .clk ( clk ), .rnd ({Fresh[8639], Fresh[8638], Fresh[8637], Fresh[8636], Fresh[8635], Fresh[8634], Fresh[8633], Fresh[8632], Fresh[8631], Fresh[8630]}), .outt ({new_AGEMA_signal_3710, new_AGEMA_signal_3709, new_AGEMA_signal_3708, n2379}) ) ;

    /* cells in depth 29 */

    /* cells in depth 30 */
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2377 ( .ina ({new_AGEMA_signal_3590, new_AGEMA_signal_3589, new_AGEMA_signal_3588, n2212}), .inb ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, new_AGEMA_signal_3705, n2211}), .clk ( clk ), .rnd ({Fresh[8649], Fresh[8648], Fresh[8647], Fresh[8646], Fresh[8645], Fresh[8644], Fresh[8643], Fresh[8642], Fresh[8641], Fresh[8640]}), .outt ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, new_AGEMA_signal_3711, N379}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2541 ( .ina ({new_AGEMA_signal_3476, new_AGEMA_signal_3475, new_AGEMA_signal_3474, n2380}), .inb ({new_AGEMA_signal_3710, new_AGEMA_signal_3709, new_AGEMA_signal_3708, n2379}), .clk ( clk ), .rnd ({Fresh[8659], Fresh[8658], Fresh[8657], Fresh[8656], Fresh[8655], Fresh[8654], Fresh[8653], Fresh[8652], Fresh[8651], Fresh[8650]}), .outt ({new_AGEMA_signal_3716, new_AGEMA_signal_3715, new_AGEMA_signal_3714, n2381}) ) ;

    /* cells in depth 31 */

    /* cells in depth 32 */
    nor_HPC1 #(.security_order(3), .pipeline(0)) U2542 ( .ina ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, new_AGEMA_signal_3471, n2382}), .inb ({new_AGEMA_signal_3716, new_AGEMA_signal_3715, new_AGEMA_signal_3714, n2381}), .clk ( clk ), .rnd ({Fresh[8669], Fresh[8668], Fresh[8667], Fresh[8666], Fresh[8665], Fresh[8664], Fresh[8663], Fresh[8662], Fresh[8661], Fresh[8660]}), .outt ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, new_AGEMA_signal_3717, n2427}) ) ;

    /* cells in depth 33 */

    /* cells in depth 34 */
    nand_HPC1 #(.security_order(3), .pipeline(0)) U2584 ( .ina ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, new_AGEMA_signal_3717, n2427}), .inb ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, new_AGEMA_signal_3555, n2426}), .clk ( clk ), .rnd ({Fresh[8679], Fresh[8678], Fresh[8677], Fresh[8676], Fresh[8675], Fresh[8674], Fresh[8673], Fresh[8672], Fresh[8671], Fresh[8670]}), .outt ({new_AGEMA_signal_3722, new_AGEMA_signal_3721, new_AGEMA_signal_3720, N563}) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(0)) SO_reg_7_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, new_AGEMA_signal_3699, N169}), .Q ({SO_s3[7], SO_s2[7], SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) SO_reg_6_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_3704, new_AGEMA_signal_3703, new_AGEMA_signal_3702, N277}), .Q ({SO_s3[6], SO_s2[6], SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) SO_reg_5_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, new_AGEMA_signal_3711, N379}), .Q ({SO_s3[5], SO_s2[5], SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) SO_reg_4_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, new_AGEMA_signal_3687, N470}), .Q ({SO_s3[4], SO_s2[4], SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) SO_reg_3_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_3722, new_AGEMA_signal_3721, new_AGEMA_signal_3720, N563}), .Q ({SO_s3[3], SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) SO_reg_2_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, new_AGEMA_signal_3693, N639}), .Q ({SO_s3[2], SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) SO_reg_1_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_3698, new_AGEMA_signal_3697, new_AGEMA_signal_3696, N723}), .Q ({SO_s3[1], SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) SO_reg_0_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, new_AGEMA_signal_3675, N789}), .Q ({SO_s3[0], SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
