/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module sbox_HPC2_AIG_ClockGating_d2 (X_s0, clk, X_s1, X_s2, Fresh, rst, Y_s0, Y_s1, Y_s2, Synch);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input rst ;
    input [101:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output Synch ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_169 ;
    wire signal_170 ;
    wire signal_171 ;
    wire signal_172 ;
    wire signal_173 ;
    wire signal_174 ;
    wire signal_175 ;
    wire signal_176 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_182 ;
    wire signal_183 ;
    wire signal_184 ;
    wire signal_185 ;
    wire signal_186 ;
    wire signal_187 ;
    wire signal_188 ;
    wire signal_189 ;
    wire signal_190 ;
    wire signal_191 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_674 ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_136 ( .a ({X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s2[4], X_s1[4], X_s0[4]}), .c ({signal_280, signal_279, signal_151}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_137 ( .a ({X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_284, signal_283, signal_152}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_138 ( .a ({X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s2[1], X_s1[1], X_s0[1]}), .c ({signal_288, signal_287, signal_153}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_139 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_290, signal_289, signal_154}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_140 ( .a ({X_s2[3], X_s1[3], X_s0[3]}), .b ({X_s2[1], X_s1[1], X_s0[1]}), .c ({signal_294, signal_293, signal_155}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_141 ( .a ({X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s2[5], X_s1[5], X_s0[5]}), .c ({signal_300, signal_299, signal_156}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_142 ( .a ({X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_302, signal_301, signal_157}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_143 ( .a ({X_s2[5], X_s1[5], X_s0[5]}), .b ({X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_304, signal_303, signal_158}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_144 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_308, signal_307, signal_159}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_145 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_310, signal_309, signal_160}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_146 ( .a ({signal_280, signal_279, signal_151}), .b ({signal_294, signal_293, signal_155}), .c ({signal_312, signal_311, signal_161}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_147 ( .a ({X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_300, signal_299, signal_156}), .c ({signal_314, signal_313, signal_162}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_148 ( .a ({signal_288, signal_287, signal_153}), .b ({signal_290, signal_289, signal_154}), .c ({signal_316, signal_315, signal_163}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_149 ( .a ({signal_294, signal_293, signal_155}), .b ({signal_302, signal_301, signal_157}), .c ({signal_318, signal_317, signal_164}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_150 ( .a ({signal_294, signal_293, signal_155}), .b ({signal_304, signal_303, signal_158}), .c ({signal_320, signal_319, signal_165}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_151 ( .a ({signal_300, signal_299, signal_156}), .b ({signal_308, signal_307, signal_159}), .c ({signal_322, signal_321, signal_166}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_152 ( .a ({signal_300, signal_299, signal_156}), .b ({signal_310, signal_309, signal_160}), .c ({signal_324, signal_323, signal_167}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_153 ( .a ({signal_280, signal_279, signal_151}), .b ({signal_304, signal_303, signal_158}), .c ({signal_326, signal_325, signal_168}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_160 ( .a ({X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_312, signal_311, signal_161}), .c ({signal_340, signal_339, signal_175}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_161 ( .a ({signal_300, signal_299, signal_156}), .b ({signal_312, signal_311, signal_161}), .c ({signal_342, signal_341, signal_176}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_162 ( .a ({signal_302, signal_301, signal_157}), .b ({signal_312, signal_311, signal_161}), .c ({signal_344, signal_343, signal_177}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_163 ( .a ({signal_314, signal_313, signal_162}), .b ({signal_320, signal_319, signal_165}), .c ({signal_346, signal_345, signal_178}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_164 ( .a ({signal_280, signal_279, signal_151}), .b ({signal_322, signal_321, signal_166}), .c ({signal_348, signal_347, signal_179}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_165 ( .a ({signal_284, signal_283, signal_152}), .b ({signal_324, signal_323, signal_167}), .c ({signal_350, signal_349, signal_180}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_166 ( .a ({signal_288, signal_287, signal_153}), .b ({signal_320, signal_319, signal_165}), .c ({signal_352, signal_351, signal_181}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_170 ( .a ({signal_284, signal_283, signal_152}), .b ({signal_342, signal_341, signal_176}), .c ({signal_360, signal_359, signal_185}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_171 ( .a ({signal_346, signal_345, signal_178}), .b ({signal_348, signal_347, signal_179}), .c ({signal_362, signal_361, signal_186}) ) ;
    ClockGatingController #(9) cell_268 ( .clk (clk), .rst (rst), .GatedClk (signal_674), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_154 ( .a ({signal_312, signal_311, signal_161}), .b ({signal_316, signal_315, signal_163}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_328, signal_327, signal_169}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_155 ( .a ({X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_322, signal_321, signal_166}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({signal_330, signal_329, signal_170}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_156 ( .a ({signal_288, signal_287, signal_153}), .b ({signal_320, signal_319, signal_165}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_332, signal_331, signal_171}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_157 ( .a ({signal_314, signal_313, signal_162}), .b ({signal_324, signal_323, signal_167}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({signal_334, signal_333, signal_172}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_158 ( .a ({signal_280, signal_279, signal_151}), .b ({signal_318, signal_317, signal_164}), .clk (clk), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_336, signal_335, signal_173}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_159 ( .a ({signal_290, signal_289, signal_154}), .b ({signal_326, signal_325, signal_168}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({signal_338, signal_337, signal_174}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_167 ( .a ({signal_340, signal_339, signal_175}), .b ({signal_350, signal_349, signal_180}), .clk (clk), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_354, signal_353, signal_182}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_168 ( .a ({signal_346, signal_345, signal_178}), .b ({signal_348, signal_347, signal_179}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({signal_356, signal_355, signal_183}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_169 ( .a ({signal_284, signal_283, signal_152}), .b ({signal_342, signal_341, signal_176}), .clk (clk), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({signal_358, signal_357, signal_184}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_172 ( .a ({signal_344, signal_343, signal_177}), .b ({signal_328, signal_327, signal_169}), .c ({signal_364, signal_363, signal_187}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_173 ( .a ({signal_328, signal_327, signal_169}), .b ({signal_330, signal_329, signal_170}), .c ({signal_366, signal_365, signal_188}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_174 ( .a ({signal_352, signal_351, signal_181}), .b ({signal_332, signal_331, signal_171}), .c ({signal_368, signal_367, signal_189}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_175 ( .a ({signal_336, signal_335, signal_173}), .b ({signal_338, signal_337, signal_174}), .c ({signal_370, signal_369, signal_190}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_176 ( .a ({signal_332, signal_331, signal_171}), .b ({signal_356, signal_355, signal_183}), .c ({signal_372, signal_371, signal_191}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_177 ( .a ({signal_336, signal_335, signal_173}), .b ({signal_358, signal_357, signal_184}), .c ({signal_374, signal_373, signal_192}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_178 ( .a ({signal_354, signal_353, signal_182}), .b ({signal_364, signal_363, signal_187}), .c ({signal_376, signal_375, signal_193}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_179 ( .a ({signal_360, signal_359, signal_185}), .b ({signal_366, signal_365, signal_188}), .c ({signal_378, signal_377, signal_194}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_180 ( .a ({signal_334, signal_333, signal_172}), .b ({signal_368, signal_367, signal_189}), .c ({signal_380, signal_379, signal_195}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_181 ( .a ({signal_372, signal_371, signal_191}), .b ({signal_374, signal_373, signal_192}), .c ({signal_382, signal_381, signal_196}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_182 ( .a ({signal_370, signal_369, signal_190}), .b ({signal_376, signal_375, signal_193}), .c ({signal_384, signal_383, signal_197}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_183 ( .a ({signal_374, signal_373, signal_192}), .b ({signal_378, signal_377, signal_194}), .c ({signal_386, signal_385, signal_198}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_184 ( .a ({signal_370, signal_369, signal_190}), .b ({signal_380, signal_379, signal_195}), .c ({signal_388, signal_387, signal_199}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_187 ( .a ({signal_362, signal_361, signal_186}), .b ({signal_382, signal_381, signal_196}), .c ({signal_394, signal_393, signal_202}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_188 ( .a ({signal_384, signal_383, signal_197}), .b ({signal_386, signal_385, signal_198}), .c ({signal_396, signal_395, signal_203}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_190 ( .a ({signal_388, signal_387, signal_199}), .b ({signal_394, signal_393, signal_202}), .c ({signal_400, signal_399, signal_205}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_185 ( .a ({signal_384, signal_383, signal_197}), .b ({signal_388, signal_387, signal_199}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({signal_390, signal_389, signal_200}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_186 ( .a ({signal_386, signal_385, signal_198}), .b ({signal_388, signal_387, signal_199}), .clk (clk), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_392, signal_391, signal_201}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_189 ( .a ({signal_384, signal_383, signal_197}), .b ({signal_394, signal_393, signal_202}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({signal_398, signal_397, signal_204}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_191 ( .a ({signal_386, signal_385, signal_198}), .b ({signal_390, signal_389, signal_200}), .c ({signal_402, signal_401, signal_206}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_192 ( .a ({signal_394, signal_393, signal_202}), .b ({signal_390, signal_389, signal_200}), .c ({signal_404, signal_403, signal_207}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_193 ( .a ({signal_390, signal_389, signal_200}), .b ({signal_396, signal_395, signal_203}), .c ({signal_406, signal_405, signal_208}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_198 ( .a ({signal_390, signal_389, signal_200}), .b ({signal_400, signal_399, signal_205}), .c ({signal_416, signal_415, signal_213}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_194 ( .a ({signal_396, signal_395, signal_203}), .b ({signal_404, signal_403, signal_207}), .clk (clk), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({signal_408, signal_407, signal_209}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_195 ( .a ({signal_400, signal_399, signal_205}), .b ({signal_402, signal_401, signal_206}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({signal_410, signal_409, signal_210}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_196 ( .a ({signal_396, signal_395, signal_203}), .b ({signal_398, signal_397, signal_204}), .clk (clk), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({signal_412, signal_411, signal_211}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_197 ( .a ({signal_392, signal_391, signal_201}), .b ({signal_400, signal_399, signal_205}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({signal_414, signal_413, signal_212}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_199 ( .a ({signal_386, signal_385, signal_198}), .b ({signal_408, signal_407, signal_209}), .c ({signal_418, signal_417, signal_214}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_200 ( .a ({signal_406, signal_405, signal_208}), .b ({signal_412, signal_411, signal_211}), .c ({signal_420, signal_419, signal_215}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_201 ( .a ({signal_394, signal_393, signal_202}), .b ({signal_410, signal_409, signal_210}), .c ({signal_422, signal_421, signal_216}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_202 ( .a ({signal_414, signal_413, signal_212}), .b ({signal_416, signal_415, signal_213}), .c ({signal_424, signal_423, signal_217}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_211 ( .a ({signal_420, signal_419, signal_215}), .b ({signal_424, signal_423, signal_217}), .c ({signal_442, signal_441, signal_226}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_212 ( .a ({signal_418, signal_417, signal_214}), .b ({signal_422, signal_421, signal_216}), .c ({signal_444, signal_443, signal_227}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_213 ( .a ({signal_418, signal_417, signal_214}), .b ({signal_420, signal_419, signal_215}), .c ({signal_446, signal_445, signal_228}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_214 ( .a ({signal_422, signal_421, signal_216}), .b ({signal_424, signal_423, signal_217}), .c ({signal_448, signal_447, signal_229}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_223 ( .a ({signal_442, signal_441, signal_226}), .b ({signal_444, signal_443, signal_227}), .c ({signal_466, signal_465, signal_238}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_203 ( .a ({signal_340, signal_339, signal_175}), .b ({signal_424, signal_423, signal_217}), .clk (clk), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({signal_426, signal_425, signal_218}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_204 ( .a ({X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_422, signal_421, signal_216}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({signal_428, signal_427, signal_219}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_205 ( .a ({signal_314, signal_313, signal_162}), .b ({signal_420, signal_419, signal_215}), .clk (clk), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({signal_430, signal_429, signal_220}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_206 ( .a ({signal_346, signal_345, signal_178}), .b ({signal_418, signal_417, signal_214}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({signal_432, signal_431, signal_221}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_207 ( .a ({signal_350, signal_349, signal_180}), .b ({signal_424, signal_423, signal_217}), .clk (clk), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_434, signal_433, signal_222}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_208 ( .a ({signal_322, signal_321, signal_166}), .b ({signal_422, signal_421, signal_216}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({signal_436, signal_435, signal_223}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_209 ( .a ({signal_324, signal_323, signal_167}), .b ({signal_420, signal_419, signal_215}), .clk (clk), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({signal_438, signal_437, signal_224}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_210 ( .a ({signal_348, signal_347, signal_179}), .b ({signal_418, signal_417, signal_214}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({signal_440, signal_439, signal_225}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_215 ( .a ({signal_312, signal_311, signal_161}), .b ({signal_448, signal_447, signal_229}), .clk (clk), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({signal_450, signal_449, signal_230}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_216 ( .a ({signal_320, signal_319, signal_165}), .b ({signal_446, signal_445, signal_228}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({signal_452, signal_451, signal_231}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_217 ( .a ({signal_318, signal_317, signal_164}), .b ({signal_444, signal_443, signal_227}), .clk (clk), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({signal_454, signal_453, signal_232}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_218 ( .a ({signal_342, signal_341, signal_176}), .b ({signal_442, signal_441, signal_226}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({signal_456, signal_455, signal_233}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_219 ( .a ({signal_316, signal_315, signal_163}), .b ({signal_448, signal_447, signal_229}), .clk (clk), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({signal_458, signal_457, signal_234}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_220 ( .a ({signal_288, signal_287, signal_153}), .b ({signal_446, signal_445, signal_228}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({signal_460, signal_459, signal_235}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_221 ( .a ({signal_280, signal_279, signal_151}), .b ({signal_444, signal_443, signal_227}), .clk (clk), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_462, signal_461, signal_236}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_222 ( .a ({signal_284, signal_283, signal_152}), .b ({signal_442, signal_441, signal_226}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({signal_464, signal_463, signal_237}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_224 ( .a ({signal_430, signal_429, signal_220}), .b ({signal_434, signal_433, signal_222}), .c ({signal_468, signal_467, signal_239}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_225 ( .a ({signal_432, signal_431, signal_221}), .b ({signal_438, signal_437, signal_224}), .c ({signal_470, signal_469, signal_240}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_226 ( .a ({signal_428, signal_427, signal_219}), .b ({signal_432, signal_431, signal_221}), .c ({signal_472, signal_471, signal_241}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_227 ( .a ({signal_326, signal_325, signal_168}), .b ({signal_466, signal_465, signal_238}), .clk (clk), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({signal_474, signal_473, signal_242}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(0)) cell_228 ( .a ({signal_290, signal_289, signal_154}), .b ({signal_466, signal_465, signal_238}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({signal_476, signal_475, signal_243}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_229 ( .a ({signal_428, signal_427, signal_219}), .b ({signal_450, signal_449, signal_230}), .c ({signal_478, signal_477, signal_244}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_230 ( .a ({signal_426, signal_425, signal_218}), .b ({signal_458, signal_457, signal_234}), .c ({signal_480, signal_479, signal_245}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_231 ( .a ({signal_456, signal_455, signal_233}), .b ({signal_460, signal_459, signal_235}), .c ({signal_482, signal_481, signal_246}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_232 ( .a ({signal_452, signal_451, signal_231}), .b ({signal_462, signal_461, signal_236}), .c ({signal_484, signal_483, signal_247}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_233 ( .a ({signal_454, signal_453, signal_232}), .b ({signal_462, signal_461, signal_236}), .c ({signal_486, signal_485, signal_248}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_234 ( .a ({signal_458, signal_457, signal_234}), .b ({signal_468, signal_467, signal_239}), .c ({signal_488, signal_487, signal_249}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_235 ( .a ({signal_436, signal_435, signal_223}), .b ({signal_468, signal_467, signal_239}), .c ({signal_490, signal_489, signal_250}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_236 ( .a ({signal_460, signal_459, signal_235}), .b ({signal_470, signal_469, signal_240}), .c ({signal_492, signal_491, signal_251}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_237 ( .a ({signal_462, signal_461, signal_236}), .b ({signal_476, signal_475, signal_243}), .c ({signal_494, signal_493, signal_252}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_238 ( .a ({signal_476, signal_475, signal_243}), .b ({signal_484, signal_483, signal_247}), .c ({signal_496, signal_495, signal_253}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_239 ( .a ({signal_450, signal_449, signal_230}), .b ({signal_480, signal_479, signal_245}), .c ({signal_498, signal_497, signal_254}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_240 ( .a ({signal_454, signal_453, signal_232}), .b ({signal_474, signal_473, signal_242}), .c ({signal_500, signal_499, signal_255}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_241 ( .a ({signal_474, signal_473, signal_242}), .b ({signal_482, signal_481, signal_246}), .c ({signal_502, signal_501, signal_256}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_242 ( .a ({signal_440, signal_439, signal_225}), .b ({signal_478, signal_477, signal_244}), .c ({signal_504, signal_503, signal_257}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_243 ( .a ({signal_464, signal_463, signal_237}), .b ({signal_482, signal_481, signal_246}), .c ({signal_506, signal_505, signal_258}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_244 ( .a ({signal_472, signal_471, signal_241}), .b ({signal_480, signal_479, signal_245}), .c ({signal_508, signal_507, signal_259}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_245 ( .a ({signal_478, signal_477, signal_244}), .b ({signal_492, signal_491, signal_251}), .c ({signal_510, signal_509, signal_260}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_246 ( .a ({signal_430, signal_429, signal_220}), .b ({signal_494, signal_493, signal_252}), .c ({signal_512, signal_511, signal_261}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_247 ( .a ({signal_434, signal_433, signal_222}), .b ({signal_494, signal_493, signal_252}), .c ({signal_514, signal_513, signal_262}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_248 ( .a ({signal_468, signal_467, signal_239}), .b ({signal_494, signal_493, signal_252}), .c ({signal_516, signal_515, signal_263}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_249 ( .a ({signal_468, signal_467, signal_239}), .b ({signal_498, signal_497, signal_254}), .c ({signal_518, signal_517, signal_264}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_250 ( .a ({signal_488, signal_487, signal_249}), .b ({signal_500, signal_499, signal_255}), .c ({signal_520, signal_519, signal_265}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_251 ( .a ({signal_496, signal_495, signal_253}), .b ({signal_502, signal_501, signal_256}), .c ({signal_522, signal_521, signal_266}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_252 ( .a ({signal_498, signal_497, signal_254}), .b ({signal_500, signal_499, signal_255}), .c ({signal_524, signal_523, signal_267}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_253 ( .a ({signal_470, signal_469, signal_240}), .b ({signal_502, signal_501, signal_256}), .c ({signal_526, signal_525, signal_268}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_254 ( .a ({signal_486, signal_485, signal_248}), .b ({signal_504, signal_503, signal_257}), .c ({signal_528, signal_527, signal_269}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_255 ( .a ({signal_490, signal_489, signal_250}), .b ({signal_504, signal_503, signal_257}), .c ({signal_530, signal_529, signal_270}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_256 ( .a ({signal_496, signal_495, signal_253}), .b ({signal_510, signal_509, signal_260}), .c ({signal_532, signal_531, signal_271}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_257 ( .a ({signal_532, signal_531, signal_271}), .b ({signal_534, signal_533, signal_150}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_258 ( .a ({signal_496, signal_495, signal_253}), .b ({signal_520, signal_519, signal_265}), .c ({signal_536, signal_535, signal_143}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_259 ( .a ({signal_514, signal_513, signal_262}), .b ({signal_524, signal_523, signal_267}), .c ({signal_538, signal_537, signal_272}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_260 ( .a ({signal_506, signal_505, signal_258}), .b ({signal_528, signal_527, signal_269}), .c ({signal_540, signal_539, signal_273}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_261 ( .a ({signal_496, signal_495, signal_253}), .b ({signal_518, signal_517, signal_264}), .c ({signal_542, signal_541, signal_146}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_262 ( .a ({signal_508, signal_507, signal_259}), .b ({signal_516, signal_515, signal_263}), .c ({signal_544, signal_543, signal_147}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_263 ( .a ({signal_522, signal_521, signal_266}), .b ({signal_530, signal_529, signal_270}), .c ({signal_546, signal_545, signal_148}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) cell_264 ( .a ({signal_512, signal_511, signal_261}), .b ({signal_526, signal_525, signal_268}), .c ({signal_548, signal_547, signal_274}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_265 ( .a ({signal_538, signal_537, signal_272}), .b ({signal_550, signal_549, signal_144}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_266 ( .a ({signal_540, signal_539, signal_273}), .b ({signal_552, signal_551, signal_145}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) cell_267 ( .a ({signal_548, signal_547, signal_274}), .b ({signal_554, signal_553, signal_149}) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(0)) cell_0 ( .clk (signal_674), .D ({signal_536, signal_535, signal_143}), .Q ({Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_1 ( .clk (signal_674), .D ({signal_550, signal_549, signal_144}), .Q ({Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_2 ( .clk (signal_674), .D ({signal_552, signal_551, signal_145}), .Q ({Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_3 ( .clk (signal_674), .D ({signal_542, signal_541, signal_146}), .Q ({Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_4 ( .clk (signal_674), .D ({signal_544, signal_543, signal_147}), .Q ({Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_5 ( .clk (signal_674), .D ({signal_546, signal_545, signal_148}), .Q ({Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_6 ( .clk (signal_674), .D ({signal_554, signal_553, signal_149}), .Q ({Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) cell_7 ( .clk (signal_674), .D ({signal_534, signal_533, signal_150}), .Q ({Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
