
module AES ( plaintext, key, reset, clk, ciphertext, done );
  (* AGEMA = "secure" *) input [127:0] plaintext;
  (* AGEMA = "secure" *) input [127:0] key;
  (* AGEMA = "clock" *)  input clk;
  (* AGEMA = "reset" *)  input reset;

  output [127:0] ciphertext;
  output done;

  wire   AKSRnotDone, LastRoundorDone, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         RoundReg_Inst_ff_SDE_0_next_state,
         RoundReg_Inst_ff_SDE_0_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_1_next_state,
         RoundReg_Inst_ff_SDE_1_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_2_next_state,
         RoundReg_Inst_ff_SDE_2_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_3_next_state,
         RoundReg_Inst_ff_SDE_3_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_4_next_state,
         RoundReg_Inst_ff_SDE_4_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_5_next_state,
         RoundReg_Inst_ff_SDE_5_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_6_next_state,
         RoundReg_Inst_ff_SDE_6_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_7_next_state,
         RoundReg_Inst_ff_SDE_7_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_8_next_state,
         RoundReg_Inst_ff_SDE_8_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_9_next_state,
         RoundReg_Inst_ff_SDE_9_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_10_next_state,
         RoundReg_Inst_ff_SDE_10_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_11_next_state,
         RoundReg_Inst_ff_SDE_11_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_12_next_state,
         RoundReg_Inst_ff_SDE_12_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_13_next_state,
         RoundReg_Inst_ff_SDE_13_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_14_next_state,
         RoundReg_Inst_ff_SDE_14_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_15_next_state,
         RoundReg_Inst_ff_SDE_15_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_16_next_state,
         RoundReg_Inst_ff_SDE_16_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_17_next_state,
         RoundReg_Inst_ff_SDE_17_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_18_next_state,
         RoundReg_Inst_ff_SDE_18_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_19_next_state,
         RoundReg_Inst_ff_SDE_19_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_20_next_state,
         RoundReg_Inst_ff_SDE_20_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_21_next_state,
         RoundReg_Inst_ff_SDE_21_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_22_next_state,
         RoundReg_Inst_ff_SDE_22_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_23_next_state,
         RoundReg_Inst_ff_SDE_23_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_24_next_state,
         RoundReg_Inst_ff_SDE_24_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_25_next_state,
         RoundReg_Inst_ff_SDE_25_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_26_next_state,
         RoundReg_Inst_ff_SDE_26_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_27_next_state,
         RoundReg_Inst_ff_SDE_27_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_28_next_state,
         RoundReg_Inst_ff_SDE_28_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_29_next_state,
         RoundReg_Inst_ff_SDE_29_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_30_next_state,
         RoundReg_Inst_ff_SDE_30_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_31_next_state,
         RoundReg_Inst_ff_SDE_31_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_32_next_state,
         RoundReg_Inst_ff_SDE_32_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_33_next_state,
         RoundReg_Inst_ff_SDE_33_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_34_next_state,
         RoundReg_Inst_ff_SDE_34_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_35_next_state,
         RoundReg_Inst_ff_SDE_35_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_36_next_state,
         RoundReg_Inst_ff_SDE_36_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_37_next_state,
         RoundReg_Inst_ff_SDE_37_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_38_next_state,
         RoundReg_Inst_ff_SDE_38_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_39_next_state,
         RoundReg_Inst_ff_SDE_39_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_40_next_state,
         RoundReg_Inst_ff_SDE_40_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_41_next_state,
         RoundReg_Inst_ff_SDE_41_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_42_next_state,
         RoundReg_Inst_ff_SDE_42_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_43_next_state,
         RoundReg_Inst_ff_SDE_43_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_44_next_state,
         RoundReg_Inst_ff_SDE_44_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_45_next_state,
         RoundReg_Inst_ff_SDE_45_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_46_next_state,
         RoundReg_Inst_ff_SDE_46_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_47_next_state,
         RoundReg_Inst_ff_SDE_47_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_48_next_state,
         RoundReg_Inst_ff_SDE_48_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_49_next_state,
         RoundReg_Inst_ff_SDE_49_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_50_next_state,
         RoundReg_Inst_ff_SDE_50_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_51_next_state,
         RoundReg_Inst_ff_SDE_51_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_52_next_state,
         RoundReg_Inst_ff_SDE_52_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_53_next_state,
         RoundReg_Inst_ff_SDE_53_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_54_next_state,
         RoundReg_Inst_ff_SDE_54_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_55_next_state,
         RoundReg_Inst_ff_SDE_55_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_56_next_state,
         RoundReg_Inst_ff_SDE_56_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_57_next_state,
         RoundReg_Inst_ff_SDE_57_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_58_next_state,
         RoundReg_Inst_ff_SDE_58_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_59_next_state,
         RoundReg_Inst_ff_SDE_59_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_60_next_state,
         RoundReg_Inst_ff_SDE_60_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_61_next_state,
         RoundReg_Inst_ff_SDE_61_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_62_next_state,
         RoundReg_Inst_ff_SDE_62_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_63_next_state,
         RoundReg_Inst_ff_SDE_63_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_64_next_state,
         RoundReg_Inst_ff_SDE_64_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_65_next_state,
         RoundReg_Inst_ff_SDE_65_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_66_next_state,
         RoundReg_Inst_ff_SDE_66_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_67_next_state,
         RoundReg_Inst_ff_SDE_67_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_68_next_state,
         RoundReg_Inst_ff_SDE_68_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_69_next_state,
         RoundReg_Inst_ff_SDE_69_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_70_next_state,
         RoundReg_Inst_ff_SDE_70_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_71_next_state,
         RoundReg_Inst_ff_SDE_71_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_72_next_state,
         RoundReg_Inst_ff_SDE_72_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_73_next_state,
         RoundReg_Inst_ff_SDE_73_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_74_next_state,
         RoundReg_Inst_ff_SDE_74_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_75_next_state,
         RoundReg_Inst_ff_SDE_75_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_76_next_state,
         RoundReg_Inst_ff_SDE_76_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_77_next_state,
         RoundReg_Inst_ff_SDE_77_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_78_next_state,
         RoundReg_Inst_ff_SDE_78_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_79_next_state,
         RoundReg_Inst_ff_SDE_79_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_80_next_state,
         RoundReg_Inst_ff_SDE_80_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_81_next_state,
         RoundReg_Inst_ff_SDE_81_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_82_next_state,
         RoundReg_Inst_ff_SDE_82_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_83_next_state,
         RoundReg_Inst_ff_SDE_83_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_84_next_state,
         RoundReg_Inst_ff_SDE_84_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_85_next_state,
         RoundReg_Inst_ff_SDE_85_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_86_next_state,
         RoundReg_Inst_ff_SDE_86_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_87_next_state,
         RoundReg_Inst_ff_SDE_87_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_88_next_state,
         RoundReg_Inst_ff_SDE_88_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_89_next_state,
         RoundReg_Inst_ff_SDE_89_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_90_next_state,
         RoundReg_Inst_ff_SDE_90_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_91_next_state,
         RoundReg_Inst_ff_SDE_91_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_92_next_state,
         RoundReg_Inst_ff_SDE_92_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_93_next_state,
         RoundReg_Inst_ff_SDE_93_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_94_next_state,
         RoundReg_Inst_ff_SDE_94_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_95_next_state,
         RoundReg_Inst_ff_SDE_95_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_96_next_state,
         RoundReg_Inst_ff_SDE_96_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_97_next_state,
         RoundReg_Inst_ff_SDE_97_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_98_next_state,
         RoundReg_Inst_ff_SDE_98_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_99_next_state,
         RoundReg_Inst_ff_SDE_99_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_100_next_state,
         RoundReg_Inst_ff_SDE_100_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_101_next_state,
         RoundReg_Inst_ff_SDE_101_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_102_next_state,
         RoundReg_Inst_ff_SDE_102_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_103_next_state,
         RoundReg_Inst_ff_SDE_103_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_104_next_state,
         RoundReg_Inst_ff_SDE_104_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_105_next_state,
         RoundReg_Inst_ff_SDE_105_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_106_next_state,
         RoundReg_Inst_ff_SDE_106_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_107_next_state,
         RoundReg_Inst_ff_SDE_107_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_108_next_state,
         RoundReg_Inst_ff_SDE_108_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_109_next_state,
         RoundReg_Inst_ff_SDE_109_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_110_next_state,
         RoundReg_Inst_ff_SDE_110_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_111_next_state,
         RoundReg_Inst_ff_SDE_111_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_112_next_state,
         RoundReg_Inst_ff_SDE_112_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_113_next_state,
         RoundReg_Inst_ff_SDE_113_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_114_next_state,
         RoundReg_Inst_ff_SDE_114_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_115_next_state,
         RoundReg_Inst_ff_SDE_115_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_116_next_state,
         RoundReg_Inst_ff_SDE_116_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_117_next_state,
         RoundReg_Inst_ff_SDE_117_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_118_next_state,
         RoundReg_Inst_ff_SDE_118_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_119_next_state,
         RoundReg_Inst_ff_SDE_119_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_120_next_state,
         RoundReg_Inst_ff_SDE_120_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_121_next_state,
         RoundReg_Inst_ff_SDE_121_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_122_next_state,
         RoundReg_Inst_ff_SDE_122_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_123_next_state,
         RoundReg_Inst_ff_SDE_123_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_124_next_state,
         RoundReg_Inst_ff_SDE_124_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_125_next_state,
         RoundReg_Inst_ff_SDE_125_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_126_next_state,
         RoundReg_Inst_ff_SDE_126_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_127_next_state,
         RoundReg_Inst_ff_SDE_127_current_state_reg_QN, MuxSboxIn_n7,
         MuxSboxIn_n6, MuxSboxIn_n5, SubBytesIns_Inst_Sbox_0_L29,
         SubBytesIns_Inst_Sbox_0_L28, SubBytesIns_Inst_Sbox_0_L27,
         SubBytesIns_Inst_Sbox_0_L26, SubBytesIns_Inst_Sbox_0_L25,
         SubBytesIns_Inst_Sbox_0_L24, SubBytesIns_Inst_Sbox_0_L23,
         SubBytesIns_Inst_Sbox_0_L22, SubBytesIns_Inst_Sbox_0_L21,
         SubBytesIns_Inst_Sbox_0_L20, SubBytesIns_Inst_Sbox_0_L19,
         SubBytesIns_Inst_Sbox_0_L18, SubBytesIns_Inst_Sbox_0_L17,
         SubBytesIns_Inst_Sbox_0_L16, SubBytesIns_Inst_Sbox_0_L15,
         SubBytesIns_Inst_Sbox_0_L14, SubBytesIns_Inst_Sbox_0_L13,
         SubBytesIns_Inst_Sbox_0_L12, SubBytesIns_Inst_Sbox_0_L11,
         SubBytesIns_Inst_Sbox_0_L10, SubBytesIns_Inst_Sbox_0_L9,
         SubBytesIns_Inst_Sbox_0_L8, SubBytesIns_Inst_Sbox_0_L7,
         SubBytesIns_Inst_Sbox_0_L6, SubBytesIns_Inst_Sbox_0_L5,
         SubBytesIns_Inst_Sbox_0_L4, SubBytesIns_Inst_Sbox_0_L3,
         SubBytesIns_Inst_Sbox_0_L2, SubBytesIns_Inst_Sbox_0_L1,
         SubBytesIns_Inst_Sbox_0_L0, SubBytesIns_Inst_Sbox_0_M63,
         SubBytesIns_Inst_Sbox_0_M62, SubBytesIns_Inst_Sbox_0_M61,
         SubBytesIns_Inst_Sbox_0_M60, SubBytesIns_Inst_Sbox_0_M59,
         SubBytesIns_Inst_Sbox_0_M58, SubBytesIns_Inst_Sbox_0_M57,
         SubBytesIns_Inst_Sbox_0_M56, SubBytesIns_Inst_Sbox_0_M55,
         SubBytesIns_Inst_Sbox_0_M54, SubBytesIns_Inst_Sbox_0_M53,
         SubBytesIns_Inst_Sbox_0_M52, SubBytesIns_Inst_Sbox_0_M51,
         SubBytesIns_Inst_Sbox_0_M50, SubBytesIns_Inst_Sbox_0_M49,
         SubBytesIns_Inst_Sbox_0_M48, SubBytesIns_Inst_Sbox_0_M47,
         SubBytesIns_Inst_Sbox_0_M46, SubBytesIns_Inst_Sbox_0_M45,
         SubBytesIns_Inst_Sbox_0_M44, SubBytesIns_Inst_Sbox_0_M43,
         SubBytesIns_Inst_Sbox_0_M42, SubBytesIns_Inst_Sbox_0_M41,
         SubBytesIns_Inst_Sbox_0_M40, SubBytesIns_Inst_Sbox_0_M39,
         SubBytesIns_Inst_Sbox_0_M38, SubBytesIns_Inst_Sbox_0_M37,
         SubBytesIns_Inst_Sbox_0_M36, SubBytesIns_Inst_Sbox_0_M35,
         SubBytesIns_Inst_Sbox_0_M34, SubBytesIns_Inst_Sbox_0_M33,
         SubBytesIns_Inst_Sbox_0_M32, SubBytesIns_Inst_Sbox_0_M31,
         SubBytesIns_Inst_Sbox_0_M30, SubBytesIns_Inst_Sbox_0_M29,
         SubBytesIns_Inst_Sbox_0_M28, SubBytesIns_Inst_Sbox_0_M27,
         SubBytesIns_Inst_Sbox_0_M26, SubBytesIns_Inst_Sbox_0_M25,
         SubBytesIns_Inst_Sbox_0_M24, SubBytesIns_Inst_Sbox_0_M23,
         SubBytesIns_Inst_Sbox_0_M22, SubBytesIns_Inst_Sbox_0_M21,
         SubBytesIns_Inst_Sbox_0_M20, SubBytesIns_Inst_Sbox_0_M19,
         SubBytesIns_Inst_Sbox_0_M18, SubBytesIns_Inst_Sbox_0_M17,
         SubBytesIns_Inst_Sbox_0_M16, SubBytesIns_Inst_Sbox_0_M15,
         SubBytesIns_Inst_Sbox_0_M14, SubBytesIns_Inst_Sbox_0_M13,
         SubBytesIns_Inst_Sbox_0_M12, SubBytesIns_Inst_Sbox_0_M11,
         SubBytesIns_Inst_Sbox_0_M10, SubBytesIns_Inst_Sbox_0_M9,
         SubBytesIns_Inst_Sbox_0_M8, SubBytesIns_Inst_Sbox_0_M7,
         SubBytesIns_Inst_Sbox_0_M6, SubBytesIns_Inst_Sbox_0_M5,
         SubBytesIns_Inst_Sbox_0_M4, SubBytesIns_Inst_Sbox_0_M3,
         SubBytesIns_Inst_Sbox_0_M2, SubBytesIns_Inst_Sbox_0_M1,
         SubBytesIns_Inst_Sbox_0_T27, SubBytesIns_Inst_Sbox_0_T26,
         SubBytesIns_Inst_Sbox_0_T25, SubBytesIns_Inst_Sbox_0_T24,
         SubBytesIns_Inst_Sbox_0_T23, SubBytesIns_Inst_Sbox_0_T22,
         SubBytesIns_Inst_Sbox_0_T21, SubBytesIns_Inst_Sbox_0_T20,
         SubBytesIns_Inst_Sbox_0_T19, SubBytesIns_Inst_Sbox_0_T18,
         SubBytesIns_Inst_Sbox_0_T17, SubBytesIns_Inst_Sbox_0_T16,
         SubBytesIns_Inst_Sbox_0_T15, SubBytesIns_Inst_Sbox_0_T14,
         SubBytesIns_Inst_Sbox_0_T13, SubBytesIns_Inst_Sbox_0_T12,
         SubBytesIns_Inst_Sbox_0_T11, SubBytesIns_Inst_Sbox_0_T10,
         SubBytesIns_Inst_Sbox_0_T9, SubBytesIns_Inst_Sbox_0_T8,
         SubBytesIns_Inst_Sbox_0_T7, SubBytesIns_Inst_Sbox_0_T6,
         SubBytesIns_Inst_Sbox_0_T5, SubBytesIns_Inst_Sbox_0_T4,
         SubBytesIns_Inst_Sbox_0_T3, SubBytesIns_Inst_Sbox_0_T2,
         SubBytesIns_Inst_Sbox_0_T1, SubBytesIns_Inst_Sbox_1_L29,
         SubBytesIns_Inst_Sbox_1_L28, SubBytesIns_Inst_Sbox_1_L27,
         SubBytesIns_Inst_Sbox_1_L26, SubBytesIns_Inst_Sbox_1_L25,
         SubBytesIns_Inst_Sbox_1_L24, SubBytesIns_Inst_Sbox_1_L23,
         SubBytesIns_Inst_Sbox_1_L22, SubBytesIns_Inst_Sbox_1_L21,
         SubBytesIns_Inst_Sbox_1_L20, SubBytesIns_Inst_Sbox_1_L19,
         SubBytesIns_Inst_Sbox_1_L18, SubBytesIns_Inst_Sbox_1_L17,
         SubBytesIns_Inst_Sbox_1_L16, SubBytesIns_Inst_Sbox_1_L15,
         SubBytesIns_Inst_Sbox_1_L14, SubBytesIns_Inst_Sbox_1_L13,
         SubBytesIns_Inst_Sbox_1_L12, SubBytesIns_Inst_Sbox_1_L11,
         SubBytesIns_Inst_Sbox_1_L10, SubBytesIns_Inst_Sbox_1_L9,
         SubBytesIns_Inst_Sbox_1_L8, SubBytesIns_Inst_Sbox_1_L7,
         SubBytesIns_Inst_Sbox_1_L6, SubBytesIns_Inst_Sbox_1_L5,
         SubBytesIns_Inst_Sbox_1_L4, SubBytesIns_Inst_Sbox_1_L3,
         SubBytesIns_Inst_Sbox_1_L2, SubBytesIns_Inst_Sbox_1_L1,
         SubBytesIns_Inst_Sbox_1_L0, SubBytesIns_Inst_Sbox_1_M63,
         SubBytesIns_Inst_Sbox_1_M62, SubBytesIns_Inst_Sbox_1_M61,
         SubBytesIns_Inst_Sbox_1_M60, SubBytesIns_Inst_Sbox_1_M59,
         SubBytesIns_Inst_Sbox_1_M58, SubBytesIns_Inst_Sbox_1_M57,
         SubBytesIns_Inst_Sbox_1_M56, SubBytesIns_Inst_Sbox_1_M55,
         SubBytesIns_Inst_Sbox_1_M54, SubBytesIns_Inst_Sbox_1_M53,
         SubBytesIns_Inst_Sbox_1_M52, SubBytesIns_Inst_Sbox_1_M51,
         SubBytesIns_Inst_Sbox_1_M50, SubBytesIns_Inst_Sbox_1_M49,
         SubBytesIns_Inst_Sbox_1_M48, SubBytesIns_Inst_Sbox_1_M47,
         SubBytesIns_Inst_Sbox_1_M46, SubBytesIns_Inst_Sbox_1_M45,
         SubBytesIns_Inst_Sbox_1_M44, SubBytesIns_Inst_Sbox_1_M43,
         SubBytesIns_Inst_Sbox_1_M42, SubBytesIns_Inst_Sbox_1_M41,
         SubBytesIns_Inst_Sbox_1_M40, SubBytesIns_Inst_Sbox_1_M39,
         SubBytesIns_Inst_Sbox_1_M38, SubBytesIns_Inst_Sbox_1_M37,
         SubBytesIns_Inst_Sbox_1_M36, SubBytesIns_Inst_Sbox_1_M35,
         SubBytesIns_Inst_Sbox_1_M34, SubBytesIns_Inst_Sbox_1_M33,
         SubBytesIns_Inst_Sbox_1_M32, SubBytesIns_Inst_Sbox_1_M31,
         SubBytesIns_Inst_Sbox_1_M30, SubBytesIns_Inst_Sbox_1_M29,
         SubBytesIns_Inst_Sbox_1_M28, SubBytesIns_Inst_Sbox_1_M27,
         SubBytesIns_Inst_Sbox_1_M26, SubBytesIns_Inst_Sbox_1_M25,
         SubBytesIns_Inst_Sbox_1_M24, SubBytesIns_Inst_Sbox_1_M23,
         SubBytesIns_Inst_Sbox_1_M22, SubBytesIns_Inst_Sbox_1_M21,
         SubBytesIns_Inst_Sbox_1_M20, SubBytesIns_Inst_Sbox_1_M19,
         SubBytesIns_Inst_Sbox_1_M18, SubBytesIns_Inst_Sbox_1_M17,
         SubBytesIns_Inst_Sbox_1_M16, SubBytesIns_Inst_Sbox_1_M15,
         SubBytesIns_Inst_Sbox_1_M14, SubBytesIns_Inst_Sbox_1_M13,
         SubBytesIns_Inst_Sbox_1_M12, SubBytesIns_Inst_Sbox_1_M11,
         SubBytesIns_Inst_Sbox_1_M10, SubBytesIns_Inst_Sbox_1_M9,
         SubBytesIns_Inst_Sbox_1_M8, SubBytesIns_Inst_Sbox_1_M7,
         SubBytesIns_Inst_Sbox_1_M6, SubBytesIns_Inst_Sbox_1_M5,
         SubBytesIns_Inst_Sbox_1_M4, SubBytesIns_Inst_Sbox_1_M3,
         SubBytesIns_Inst_Sbox_1_M2, SubBytesIns_Inst_Sbox_1_M1,
         SubBytesIns_Inst_Sbox_1_T27, SubBytesIns_Inst_Sbox_1_T26,
         SubBytesIns_Inst_Sbox_1_T25, SubBytesIns_Inst_Sbox_1_T24,
         SubBytesIns_Inst_Sbox_1_T23, SubBytesIns_Inst_Sbox_1_T22,
         SubBytesIns_Inst_Sbox_1_T21, SubBytesIns_Inst_Sbox_1_T20,
         SubBytesIns_Inst_Sbox_1_T19, SubBytesIns_Inst_Sbox_1_T18,
         SubBytesIns_Inst_Sbox_1_T17, SubBytesIns_Inst_Sbox_1_T16,
         SubBytesIns_Inst_Sbox_1_T15, SubBytesIns_Inst_Sbox_1_T14,
         SubBytesIns_Inst_Sbox_1_T13, SubBytesIns_Inst_Sbox_1_T12,
         SubBytesIns_Inst_Sbox_1_T11, SubBytesIns_Inst_Sbox_1_T10,
         SubBytesIns_Inst_Sbox_1_T9, SubBytesIns_Inst_Sbox_1_T8,
         SubBytesIns_Inst_Sbox_1_T7, SubBytesIns_Inst_Sbox_1_T6,
         SubBytesIns_Inst_Sbox_1_T5, SubBytesIns_Inst_Sbox_1_T4,
         SubBytesIns_Inst_Sbox_1_T3, SubBytesIns_Inst_Sbox_1_T2,
         SubBytesIns_Inst_Sbox_1_T1, SubBytesIns_Inst_Sbox_2_L29,
         SubBytesIns_Inst_Sbox_2_L28, SubBytesIns_Inst_Sbox_2_L27,
         SubBytesIns_Inst_Sbox_2_L26, SubBytesIns_Inst_Sbox_2_L25,
         SubBytesIns_Inst_Sbox_2_L24, SubBytesIns_Inst_Sbox_2_L23,
         SubBytesIns_Inst_Sbox_2_L22, SubBytesIns_Inst_Sbox_2_L21,
         SubBytesIns_Inst_Sbox_2_L20, SubBytesIns_Inst_Sbox_2_L19,
         SubBytesIns_Inst_Sbox_2_L18, SubBytesIns_Inst_Sbox_2_L17,
         SubBytesIns_Inst_Sbox_2_L16, SubBytesIns_Inst_Sbox_2_L15,
         SubBytesIns_Inst_Sbox_2_L14, SubBytesIns_Inst_Sbox_2_L13,
         SubBytesIns_Inst_Sbox_2_L12, SubBytesIns_Inst_Sbox_2_L11,
         SubBytesIns_Inst_Sbox_2_L10, SubBytesIns_Inst_Sbox_2_L9,
         SubBytesIns_Inst_Sbox_2_L8, SubBytesIns_Inst_Sbox_2_L7,
         SubBytesIns_Inst_Sbox_2_L6, SubBytesIns_Inst_Sbox_2_L5,
         SubBytesIns_Inst_Sbox_2_L4, SubBytesIns_Inst_Sbox_2_L3,
         SubBytesIns_Inst_Sbox_2_L2, SubBytesIns_Inst_Sbox_2_L1,
         SubBytesIns_Inst_Sbox_2_L0, SubBytesIns_Inst_Sbox_2_M63,
         SubBytesIns_Inst_Sbox_2_M62, SubBytesIns_Inst_Sbox_2_M61,
         SubBytesIns_Inst_Sbox_2_M60, SubBytesIns_Inst_Sbox_2_M59,
         SubBytesIns_Inst_Sbox_2_M58, SubBytesIns_Inst_Sbox_2_M57,
         SubBytesIns_Inst_Sbox_2_M56, SubBytesIns_Inst_Sbox_2_M55,
         SubBytesIns_Inst_Sbox_2_M54, SubBytesIns_Inst_Sbox_2_M53,
         SubBytesIns_Inst_Sbox_2_M52, SubBytesIns_Inst_Sbox_2_M51,
         SubBytesIns_Inst_Sbox_2_M50, SubBytesIns_Inst_Sbox_2_M49,
         SubBytesIns_Inst_Sbox_2_M48, SubBytesIns_Inst_Sbox_2_M47,
         SubBytesIns_Inst_Sbox_2_M46, SubBytesIns_Inst_Sbox_2_M45,
         SubBytesIns_Inst_Sbox_2_M44, SubBytesIns_Inst_Sbox_2_M43,
         SubBytesIns_Inst_Sbox_2_M42, SubBytesIns_Inst_Sbox_2_M41,
         SubBytesIns_Inst_Sbox_2_M40, SubBytesIns_Inst_Sbox_2_M39,
         SubBytesIns_Inst_Sbox_2_M38, SubBytesIns_Inst_Sbox_2_M37,
         SubBytesIns_Inst_Sbox_2_M36, SubBytesIns_Inst_Sbox_2_M35,
         SubBytesIns_Inst_Sbox_2_M34, SubBytesIns_Inst_Sbox_2_M33,
         SubBytesIns_Inst_Sbox_2_M32, SubBytesIns_Inst_Sbox_2_M31,
         SubBytesIns_Inst_Sbox_2_M30, SubBytesIns_Inst_Sbox_2_M29,
         SubBytesIns_Inst_Sbox_2_M28, SubBytesIns_Inst_Sbox_2_M27,
         SubBytesIns_Inst_Sbox_2_M26, SubBytesIns_Inst_Sbox_2_M25,
         SubBytesIns_Inst_Sbox_2_M24, SubBytesIns_Inst_Sbox_2_M23,
         SubBytesIns_Inst_Sbox_2_M22, SubBytesIns_Inst_Sbox_2_M21,
         SubBytesIns_Inst_Sbox_2_M20, SubBytesIns_Inst_Sbox_2_M19,
         SubBytesIns_Inst_Sbox_2_M18, SubBytesIns_Inst_Sbox_2_M17,
         SubBytesIns_Inst_Sbox_2_M16, SubBytesIns_Inst_Sbox_2_M15,
         SubBytesIns_Inst_Sbox_2_M14, SubBytesIns_Inst_Sbox_2_M13,
         SubBytesIns_Inst_Sbox_2_M12, SubBytesIns_Inst_Sbox_2_M11,
         SubBytesIns_Inst_Sbox_2_M10, SubBytesIns_Inst_Sbox_2_M9,
         SubBytesIns_Inst_Sbox_2_M8, SubBytesIns_Inst_Sbox_2_M7,
         SubBytesIns_Inst_Sbox_2_M6, SubBytesIns_Inst_Sbox_2_M5,
         SubBytesIns_Inst_Sbox_2_M4, SubBytesIns_Inst_Sbox_2_M3,
         SubBytesIns_Inst_Sbox_2_M2, SubBytesIns_Inst_Sbox_2_M1,
         SubBytesIns_Inst_Sbox_2_T27, SubBytesIns_Inst_Sbox_2_T26,
         SubBytesIns_Inst_Sbox_2_T25, SubBytesIns_Inst_Sbox_2_T24,
         SubBytesIns_Inst_Sbox_2_T23, SubBytesIns_Inst_Sbox_2_T22,
         SubBytesIns_Inst_Sbox_2_T21, SubBytesIns_Inst_Sbox_2_T20,
         SubBytesIns_Inst_Sbox_2_T19, SubBytesIns_Inst_Sbox_2_T18,
         SubBytesIns_Inst_Sbox_2_T17, SubBytesIns_Inst_Sbox_2_T16,
         SubBytesIns_Inst_Sbox_2_T15, SubBytesIns_Inst_Sbox_2_T14,
         SubBytesIns_Inst_Sbox_2_T13, SubBytesIns_Inst_Sbox_2_T12,
         SubBytesIns_Inst_Sbox_2_T11, SubBytesIns_Inst_Sbox_2_T10,
         SubBytesIns_Inst_Sbox_2_T9, SubBytesIns_Inst_Sbox_2_T8,
         SubBytesIns_Inst_Sbox_2_T7, SubBytesIns_Inst_Sbox_2_T6,
         SubBytesIns_Inst_Sbox_2_T5, SubBytesIns_Inst_Sbox_2_T4,
         SubBytesIns_Inst_Sbox_2_T3, SubBytesIns_Inst_Sbox_2_T2,
         SubBytesIns_Inst_Sbox_2_T1, SubBytesIns_Inst_Sbox_3_L29,
         SubBytesIns_Inst_Sbox_3_L28, SubBytesIns_Inst_Sbox_3_L27,
         SubBytesIns_Inst_Sbox_3_L26, SubBytesIns_Inst_Sbox_3_L25,
         SubBytesIns_Inst_Sbox_3_L24, SubBytesIns_Inst_Sbox_3_L23,
         SubBytesIns_Inst_Sbox_3_L22, SubBytesIns_Inst_Sbox_3_L21,
         SubBytesIns_Inst_Sbox_3_L20, SubBytesIns_Inst_Sbox_3_L19,
         SubBytesIns_Inst_Sbox_3_L18, SubBytesIns_Inst_Sbox_3_L17,
         SubBytesIns_Inst_Sbox_3_L16, SubBytesIns_Inst_Sbox_3_L15,
         SubBytesIns_Inst_Sbox_3_L14, SubBytesIns_Inst_Sbox_3_L13,
         SubBytesIns_Inst_Sbox_3_L12, SubBytesIns_Inst_Sbox_3_L11,
         SubBytesIns_Inst_Sbox_3_L10, SubBytesIns_Inst_Sbox_3_L9,
         SubBytesIns_Inst_Sbox_3_L8, SubBytesIns_Inst_Sbox_3_L7,
         SubBytesIns_Inst_Sbox_3_L6, SubBytesIns_Inst_Sbox_3_L5,
         SubBytesIns_Inst_Sbox_3_L4, SubBytesIns_Inst_Sbox_3_L3,
         SubBytesIns_Inst_Sbox_3_L2, SubBytesIns_Inst_Sbox_3_L1,
         SubBytesIns_Inst_Sbox_3_L0, SubBytesIns_Inst_Sbox_3_M63,
         SubBytesIns_Inst_Sbox_3_M62, SubBytesIns_Inst_Sbox_3_M61,
         SubBytesIns_Inst_Sbox_3_M60, SubBytesIns_Inst_Sbox_3_M59,
         SubBytesIns_Inst_Sbox_3_M58, SubBytesIns_Inst_Sbox_3_M57,
         SubBytesIns_Inst_Sbox_3_M56, SubBytesIns_Inst_Sbox_3_M55,
         SubBytesIns_Inst_Sbox_3_M54, SubBytesIns_Inst_Sbox_3_M53,
         SubBytesIns_Inst_Sbox_3_M52, SubBytesIns_Inst_Sbox_3_M51,
         SubBytesIns_Inst_Sbox_3_M50, SubBytesIns_Inst_Sbox_3_M49,
         SubBytesIns_Inst_Sbox_3_M48, SubBytesIns_Inst_Sbox_3_M47,
         SubBytesIns_Inst_Sbox_3_M46, SubBytesIns_Inst_Sbox_3_M45,
         SubBytesIns_Inst_Sbox_3_M44, SubBytesIns_Inst_Sbox_3_M43,
         SubBytesIns_Inst_Sbox_3_M42, SubBytesIns_Inst_Sbox_3_M41,
         SubBytesIns_Inst_Sbox_3_M40, SubBytesIns_Inst_Sbox_3_M39,
         SubBytesIns_Inst_Sbox_3_M38, SubBytesIns_Inst_Sbox_3_M37,
         SubBytesIns_Inst_Sbox_3_M36, SubBytesIns_Inst_Sbox_3_M35,
         SubBytesIns_Inst_Sbox_3_M34, SubBytesIns_Inst_Sbox_3_M33,
         SubBytesIns_Inst_Sbox_3_M32, SubBytesIns_Inst_Sbox_3_M31,
         SubBytesIns_Inst_Sbox_3_M30, SubBytesIns_Inst_Sbox_3_M29,
         SubBytesIns_Inst_Sbox_3_M28, SubBytesIns_Inst_Sbox_3_M27,
         SubBytesIns_Inst_Sbox_3_M26, SubBytesIns_Inst_Sbox_3_M25,
         SubBytesIns_Inst_Sbox_3_M24, SubBytesIns_Inst_Sbox_3_M23,
         SubBytesIns_Inst_Sbox_3_M22, SubBytesIns_Inst_Sbox_3_M21,
         SubBytesIns_Inst_Sbox_3_M20, SubBytesIns_Inst_Sbox_3_M19,
         SubBytesIns_Inst_Sbox_3_M18, SubBytesIns_Inst_Sbox_3_M17,
         SubBytesIns_Inst_Sbox_3_M16, SubBytesIns_Inst_Sbox_3_M15,
         SubBytesIns_Inst_Sbox_3_M14, SubBytesIns_Inst_Sbox_3_M13,
         SubBytesIns_Inst_Sbox_3_M12, SubBytesIns_Inst_Sbox_3_M11,
         SubBytesIns_Inst_Sbox_3_M10, SubBytesIns_Inst_Sbox_3_M9,
         SubBytesIns_Inst_Sbox_3_M8, SubBytesIns_Inst_Sbox_3_M7,
         SubBytesIns_Inst_Sbox_3_M6, SubBytesIns_Inst_Sbox_3_M5,
         SubBytesIns_Inst_Sbox_3_M4, SubBytesIns_Inst_Sbox_3_M3,
         SubBytesIns_Inst_Sbox_3_M2, SubBytesIns_Inst_Sbox_3_M1,
         SubBytesIns_Inst_Sbox_3_T27, SubBytesIns_Inst_Sbox_3_T26,
         SubBytesIns_Inst_Sbox_3_T25, SubBytesIns_Inst_Sbox_3_T24,
         SubBytesIns_Inst_Sbox_3_T23, SubBytesIns_Inst_Sbox_3_T22,
         SubBytesIns_Inst_Sbox_3_T21, SubBytesIns_Inst_Sbox_3_T20,
         SubBytesIns_Inst_Sbox_3_T19, SubBytesIns_Inst_Sbox_3_T18,
         SubBytesIns_Inst_Sbox_3_T17, SubBytesIns_Inst_Sbox_3_T16,
         SubBytesIns_Inst_Sbox_3_T15, SubBytesIns_Inst_Sbox_3_T14,
         SubBytesIns_Inst_Sbox_3_T13, SubBytesIns_Inst_Sbox_3_T12,
         SubBytesIns_Inst_Sbox_3_T11, SubBytesIns_Inst_Sbox_3_T10,
         SubBytesIns_Inst_Sbox_3_T9, SubBytesIns_Inst_Sbox_3_T8,
         SubBytesIns_Inst_Sbox_3_T7, SubBytesIns_Inst_Sbox_3_T6,
         SubBytesIns_Inst_Sbox_3_T5, SubBytesIns_Inst_Sbox_3_T4,
         SubBytesIns_Inst_Sbox_3_T3, SubBytesIns_Inst_Sbox_3_T2,
         SubBytesIns_Inst_Sbox_3_T1, MixColumnsIns_n64, MixColumnsIns_n63,
         MixColumnsIns_n62, MixColumnsIns_n61, MixColumnsIns_n60,
         MixColumnsIns_n59, MixColumnsIns_n58, MixColumnsIns_n57,
         MixColumnsIns_n56, MixColumnsIns_n55, MixColumnsIns_n54,
         MixColumnsIns_n53, MixColumnsIns_n52, MixColumnsIns_n51,
         MixColumnsIns_n50, MixColumnsIns_n49, MixColumnsIns_n48,
         MixColumnsIns_n47, MixColumnsIns_n46, MixColumnsIns_n45,
         MixColumnsIns_n44, MixColumnsIns_n43, MixColumnsIns_n42,
         MixColumnsIns_n41, MixColumnsIns_n40, MixColumnsIns_n39,
         MixColumnsIns_n38, MixColumnsIns_n37, MixColumnsIns_n36,
         MixColumnsIns_n35, MixColumnsIns_n34, MixColumnsIns_n33,
         MixColumnsIns_n32, MixColumnsIns_n31, MixColumnsIns_n30,
         MixColumnsIns_n29, MixColumnsIns_n28, MixColumnsIns_n27,
         MixColumnsIns_n26, MixColumnsIns_n25, MixColumnsIns_n24,
         MixColumnsIns_n23, MixColumnsIns_n22, MixColumnsIns_n21,
         MixColumnsIns_n20, MixColumnsIns_n19, MixColumnsIns_n18,
         MixColumnsIns_n17, MixColumnsIns_n16, MixColumnsIns_n15,
         MixColumnsIns_n14, MixColumnsIns_n13, MixColumnsIns_n12,
         MixColumnsIns_n11, MixColumnsIns_n10, MixColumnsIns_n9,
         MixColumnsIns_n8, MixColumnsIns_n7, MixColumnsIns_n6,
         MixColumnsIns_n5, MixColumnsIns_n4, MixColumnsIns_n3,
         MixColumnsIns_n2, MixColumnsIns_n1, MuxMCOut_n6, MuxMCOut_n5,
         MuxMCOut_n4, MuxRound_n19, MuxRound_n18, MuxRound_n17, MuxRound_n16,
         MuxRound_n15, MuxRound_n14, MuxRound_n13,
         KeyReg_Inst_ff_SDE_0_next_state,
         KeyReg_Inst_ff_SDE_0_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_1_next_state,
         KeyReg_Inst_ff_SDE_1_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_2_next_state,
         KeyReg_Inst_ff_SDE_2_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_3_next_state,
         KeyReg_Inst_ff_SDE_3_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_4_next_state,
         KeyReg_Inst_ff_SDE_4_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_5_next_state,
         KeyReg_Inst_ff_SDE_5_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_6_next_state,
         KeyReg_Inst_ff_SDE_6_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_7_next_state,
         KeyReg_Inst_ff_SDE_7_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_8_next_state,
         KeyReg_Inst_ff_SDE_8_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_9_next_state,
         KeyReg_Inst_ff_SDE_9_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_10_next_state,
         KeyReg_Inst_ff_SDE_10_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_11_next_state,
         KeyReg_Inst_ff_SDE_11_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_12_next_state,
         KeyReg_Inst_ff_SDE_12_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_13_next_state,
         KeyReg_Inst_ff_SDE_13_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_14_next_state,
         KeyReg_Inst_ff_SDE_14_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_15_next_state,
         KeyReg_Inst_ff_SDE_15_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_16_next_state,
         KeyReg_Inst_ff_SDE_16_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_17_next_state,
         KeyReg_Inst_ff_SDE_17_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_18_next_state,
         KeyReg_Inst_ff_SDE_18_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_19_next_state,
         KeyReg_Inst_ff_SDE_19_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_20_next_state,
         KeyReg_Inst_ff_SDE_20_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_21_next_state,
         KeyReg_Inst_ff_SDE_21_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_22_next_state,
         KeyReg_Inst_ff_SDE_22_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_23_next_state,
         KeyReg_Inst_ff_SDE_23_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_24_next_state,
         KeyReg_Inst_ff_SDE_24_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_25_next_state,
         KeyReg_Inst_ff_SDE_25_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_26_next_state,
         KeyReg_Inst_ff_SDE_26_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_27_next_state,
         KeyReg_Inst_ff_SDE_27_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_28_next_state,
         KeyReg_Inst_ff_SDE_28_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_29_next_state,
         KeyReg_Inst_ff_SDE_29_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_30_next_state,
         KeyReg_Inst_ff_SDE_30_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_31_next_state,
         KeyReg_Inst_ff_SDE_31_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_32_next_state,
         KeyReg_Inst_ff_SDE_32_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_33_next_state,
         KeyReg_Inst_ff_SDE_33_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_34_next_state,
         KeyReg_Inst_ff_SDE_34_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_35_next_state,
         KeyReg_Inst_ff_SDE_35_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_36_next_state,
         KeyReg_Inst_ff_SDE_36_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_37_next_state,
         KeyReg_Inst_ff_SDE_37_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_38_next_state,
         KeyReg_Inst_ff_SDE_38_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_39_next_state,
         KeyReg_Inst_ff_SDE_39_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_40_next_state,
         KeyReg_Inst_ff_SDE_40_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_41_next_state,
         KeyReg_Inst_ff_SDE_41_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_42_next_state,
         KeyReg_Inst_ff_SDE_42_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_43_next_state,
         KeyReg_Inst_ff_SDE_43_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_44_next_state,
         KeyReg_Inst_ff_SDE_44_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_45_next_state,
         KeyReg_Inst_ff_SDE_45_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_46_next_state,
         KeyReg_Inst_ff_SDE_46_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_47_next_state,
         KeyReg_Inst_ff_SDE_47_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_48_next_state,
         KeyReg_Inst_ff_SDE_48_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_49_next_state,
         KeyReg_Inst_ff_SDE_49_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_50_next_state,
         KeyReg_Inst_ff_SDE_50_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_51_next_state,
         KeyReg_Inst_ff_SDE_51_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_52_next_state,
         KeyReg_Inst_ff_SDE_52_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_53_next_state,
         KeyReg_Inst_ff_SDE_53_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_54_next_state,
         KeyReg_Inst_ff_SDE_54_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_55_next_state,
         KeyReg_Inst_ff_SDE_55_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_56_next_state,
         KeyReg_Inst_ff_SDE_56_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_57_next_state,
         KeyReg_Inst_ff_SDE_57_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_58_next_state,
         KeyReg_Inst_ff_SDE_58_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_59_next_state,
         KeyReg_Inst_ff_SDE_59_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_60_next_state,
         KeyReg_Inst_ff_SDE_60_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_61_next_state,
         KeyReg_Inst_ff_SDE_61_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_62_next_state,
         KeyReg_Inst_ff_SDE_62_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_63_next_state,
         KeyReg_Inst_ff_SDE_63_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_64_next_state,
         KeyReg_Inst_ff_SDE_64_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_65_next_state,
         KeyReg_Inst_ff_SDE_65_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_66_next_state,
         KeyReg_Inst_ff_SDE_66_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_67_next_state,
         KeyReg_Inst_ff_SDE_67_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_68_next_state,
         KeyReg_Inst_ff_SDE_68_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_69_next_state,
         KeyReg_Inst_ff_SDE_69_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_70_next_state,
         KeyReg_Inst_ff_SDE_70_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_71_next_state,
         KeyReg_Inst_ff_SDE_71_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_72_next_state,
         KeyReg_Inst_ff_SDE_72_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_73_next_state,
         KeyReg_Inst_ff_SDE_73_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_74_next_state,
         KeyReg_Inst_ff_SDE_74_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_75_next_state,
         KeyReg_Inst_ff_SDE_75_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_76_next_state,
         KeyReg_Inst_ff_SDE_76_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_77_next_state,
         KeyReg_Inst_ff_SDE_77_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_78_next_state,
         KeyReg_Inst_ff_SDE_78_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_79_next_state,
         KeyReg_Inst_ff_SDE_79_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_80_next_state,
         KeyReg_Inst_ff_SDE_80_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_81_next_state,
         KeyReg_Inst_ff_SDE_81_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_82_next_state,
         KeyReg_Inst_ff_SDE_82_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_83_next_state,
         KeyReg_Inst_ff_SDE_83_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_84_next_state,
         KeyReg_Inst_ff_SDE_84_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_85_next_state,
         KeyReg_Inst_ff_SDE_85_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_86_next_state,
         KeyReg_Inst_ff_SDE_86_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_87_next_state,
         KeyReg_Inst_ff_SDE_87_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_88_next_state,
         KeyReg_Inst_ff_SDE_88_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_89_next_state,
         KeyReg_Inst_ff_SDE_89_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_90_next_state,
         KeyReg_Inst_ff_SDE_90_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_91_next_state,
         KeyReg_Inst_ff_SDE_91_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_92_next_state,
         KeyReg_Inst_ff_SDE_92_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_93_next_state,
         KeyReg_Inst_ff_SDE_93_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_94_next_state,
         KeyReg_Inst_ff_SDE_94_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_95_next_state,
         KeyReg_Inst_ff_SDE_95_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_96_next_state,
         KeyReg_Inst_ff_SDE_96_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_97_next_state,
         KeyReg_Inst_ff_SDE_97_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_98_next_state,
         KeyReg_Inst_ff_SDE_98_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_99_next_state,
         KeyReg_Inst_ff_SDE_99_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_100_next_state,
         KeyReg_Inst_ff_SDE_100_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_101_next_state,
         KeyReg_Inst_ff_SDE_101_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_102_next_state,
         KeyReg_Inst_ff_SDE_102_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_103_next_state,
         KeyReg_Inst_ff_SDE_103_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_104_next_state,
         KeyReg_Inst_ff_SDE_104_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_105_next_state,
         KeyReg_Inst_ff_SDE_105_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_106_next_state,
         KeyReg_Inst_ff_SDE_106_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_107_next_state,
         KeyReg_Inst_ff_SDE_107_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_108_next_state,
         KeyReg_Inst_ff_SDE_108_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_109_next_state,
         KeyReg_Inst_ff_SDE_109_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_110_next_state,
         KeyReg_Inst_ff_SDE_110_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_111_next_state,
         KeyReg_Inst_ff_SDE_111_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_112_next_state,
         KeyReg_Inst_ff_SDE_112_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_113_next_state,
         KeyReg_Inst_ff_SDE_113_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_114_next_state,
         KeyReg_Inst_ff_SDE_114_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_115_next_state,
         KeyReg_Inst_ff_SDE_115_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_116_next_state,
         KeyReg_Inst_ff_SDE_116_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_117_next_state,
         KeyReg_Inst_ff_SDE_117_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_118_next_state,
         KeyReg_Inst_ff_SDE_118_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_119_next_state,
         KeyReg_Inst_ff_SDE_119_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_120_next_state,
         KeyReg_Inst_ff_SDE_120_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_121_next_state,
         KeyReg_Inst_ff_SDE_121_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_122_next_state,
         KeyReg_Inst_ff_SDE_122_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_123_next_state,
         KeyReg_Inst_ff_SDE_123_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_124_next_state,
         KeyReg_Inst_ff_SDE_124_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_125_next_state,
         KeyReg_Inst_ff_SDE_125_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_126_next_state,
         KeyReg_Inst_ff_SDE_126_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_127_next_state,
         KeyReg_Inst_ff_SDE_127_current_state_reg_QN, MuxKeyExpansion_n21,
         MuxKeyExpansion_n20, MuxKeyExpansion_n19, MuxKeyExpansion_n18,
         MuxKeyExpansion_n17, MuxKeyExpansion_n16, MuxKeyExpansion_n15,
         MuxKeyExpansion_n14, RoundCounterIns_n10, RoundCounterIns_n9,
         RoundCounterIns_n8, RoundCounterIns_n7, RoundCounterIns_n6,
         RoundCounterIns_n5, RoundCounterIns_n4, RoundCounterIns_n42,
         RoundCounterIns_n1, RoundCounterIns_n2, RoundCounterIns_n44,
         RoundCounterIns_n45, RoundCounterIns_count_reg_0__QN,
         RoundCounterIns_count_reg_2__QN, RoundCounterIns_count_reg_3__QN,
         InRoundCounterIns_n12, InRoundCounterIns_n11, InRoundCounterIns_n10,
         InRoundCounterIns_n9, InRoundCounterIns_n8, InRoundCounterIns_n7,
         InRoundCounterIns_n5, InRoundCounterIns_n4, InRoundCounterIns_n3,
         InRoundCounterIns_n2, InRoundCounterIns_n1, InRoundCounterIns_n6,
         InRoundCounterIns_n39, InRoundCounterIns_n40, InRoundCounterIns_n41,
         InRoundCounterIns_count_reg_0__QN;
  wire   [127:0] RoundOutput;
  wire   [127:0] ShiftRowsOutput;
  wire   [31:0] KSSubBytesInput;
  wire   [31:0] SubBytesInput;
  wire   [3:0] SubBytesOutput;
  wire   [31:0] MixColumnsOutput;
  wire   [31:0] ColumnOutput;
  wire   [127:0] RoundKeyOutput;
  wire   [127:32] RoundKey;
  wire   [7:0] Rcon;
  wire   [127:0] KeyExpansionOutput;
  wire   [3:0] RoundCounter;
  wire   [2:0] InRoundCounter;
  wire   [28:0] MixColumnsIns_DoubleBytes;
  wire   [31:0] KeyExpansionIns_tmp;

  AND2_X1 U323 ( .A1(n45), .A2(n44), .ZN(AKSRnotDone) );
  NOR2_X1 U324 ( .A1(n60), .A2(n49), .ZN(LastRoundorDone) );
  AND2_X1 U325 ( .A1(RoundCounter[0]), .A2(LastRoundorDone), .ZN(done) );
  INV_X1 U326 ( .A(RoundCounter[3]), .ZN(n60) );
  NOR2_X1 U327 ( .A1(InRoundCounter[0]), .A2(InRoundCounter[1]), .ZN(n45) );
  INV_X1 U328 ( .A(RoundCounter[2]), .ZN(n46) );
  NAND2_X1 U329 ( .A1(RoundCounter[1]), .A2(n46), .ZN(n49) );
  NOR2_X1 U330 ( .A1(done), .A2(InRoundCounter[2]), .ZN(n44) );
  INV_X1 U331 ( .A(RoundCounter[1]), .ZN(n55) );
  NAND2_X1 U332 ( .A1(n55), .A2(n46), .ZN(n47) );
  NOR2_X1 U333 ( .A1(RoundCounter[0]), .A2(n47), .ZN(Rcon[0]) );
  NOR2_X1 U334 ( .A1(RoundCounter[0]), .A2(RoundCounter[3]), .ZN(n58) );
  NOR2_X1 U335 ( .A1(n58), .A2(n47), .ZN(Rcon[1]) );
  NOR2_X1 U336 ( .A1(RoundCounter[3]), .A2(n49), .ZN(n48) );
  NOR2_X1 U337 ( .A1(n60), .A2(n47), .ZN(n54) );
  MUX2_X1 U338 ( .A(n48), .B(n54), .S(RoundCounter[0]), .Z(Rcon[2]) );
  INV_X1 U339 ( .A(RoundCounter[0]), .ZN(n50) );
  NOR2_X1 U340 ( .A1(n50), .A2(n49), .ZN(n51) );
  MUX2_X1 U341 ( .A(n51), .B(Rcon[0]), .S(RoundCounter[3]), .Z(Rcon[3]) );
  NAND2_X1 U342 ( .A1(RoundCounter[2]), .A2(n58), .ZN(n52) );
  NOR2_X1 U343 ( .A1(RoundCounter[1]), .A2(n52), .ZN(n53) );
  OR2_X1 U344 ( .A1(n54), .A2(n53), .ZN(Rcon[4]) );
  XNOR2_X1 U345 ( .A(RoundCounter[2]), .B(RoundCounter[3]), .ZN(n57) );
  NAND2_X1 U346 ( .A1(RoundCounter[0]), .A2(n55), .ZN(n56) );
  NOR2_X1 U347 ( .A1(n57), .A2(n56), .ZN(Rcon[5]) );
  INV_X1 U348 ( .A(n58), .ZN(n59) );
  NAND2_X1 U349 ( .A1(RoundCounter[1]), .A2(RoundCounter[2]), .ZN(n61) );
  NOR2_X1 U350 ( .A1(n59), .A2(n61), .ZN(Rcon[6]) );
  NAND2_X1 U351 ( .A1(RoundCounter[0]), .A2(n60), .ZN(n62) );
  NOR2_X1 U352 ( .A1(n62), .A2(n61), .ZN(Rcon[7]) );
  XOR2_X1 U353 ( .A(ciphertext[32]), .B(KSSubBytesInput[16]), .Z(
        ShiftRowsOutput[96]) );
  XOR2_X1 U354 ( .A(ciphertext[4]), .B(RoundKey[100]), .Z(ShiftRowsOutput[68])
         );
  XOR2_X1 U355 ( .A(ciphertext[5]), .B(RoundKey[101]), .Z(ShiftRowsOutput[69])
         );
  XOR2_X1 U356 ( .A(ciphertext[6]), .B(RoundKey[102]), .Z(ShiftRowsOutput[70])
         );
  XOR2_X1 U357 ( .A(ciphertext[7]), .B(RoundKey[103]), .Z(ShiftRowsOutput[71])
         );
  XOR2_X1 U358 ( .A(ciphertext[40]), .B(RoundKey[104]), .Z(ShiftRowsOutput[40]) );
  XOR2_X1 U359 ( .A(ciphertext[41]), .B(RoundKey[105]), .Z(ShiftRowsOutput[41]) );
  XOR2_X1 U360 ( .A(ciphertext[42]), .B(RoundKey[106]), .Z(ShiftRowsOutput[42]) );
  XOR2_X1 U361 ( .A(ciphertext[43]), .B(RoundKey[107]), .Z(ShiftRowsOutput[43]) );
  XOR2_X1 U362 ( .A(ciphertext[44]), .B(RoundKey[108]), .Z(ShiftRowsOutput[44]) );
  XOR2_X1 U363 ( .A(ciphertext[45]), .B(RoundKey[109]), .Z(ShiftRowsOutput[45]) );
  XOR2_X1 U364 ( .A(ciphertext[74]), .B(KSSubBytesInput[10]), .Z(
        ShiftRowsOutput[74]) );
  XOR2_X1 U365 ( .A(ciphertext[46]), .B(RoundKey[110]), .Z(ShiftRowsOutput[46]) );
  XOR2_X1 U366 ( .A(ciphertext[47]), .B(RoundKey[111]), .Z(ShiftRowsOutput[47]) );
  XOR2_X1 U367 ( .A(ciphertext[80]), .B(RoundKey[112]), .Z(ShiftRowsOutput[16]) );
  XOR2_X1 U368 ( .A(ciphertext[81]), .B(RoundKey[113]), .Z(ShiftRowsOutput[17]) );
  XOR2_X1 U369 ( .A(ciphertext[82]), .B(RoundKey[114]), .Z(ShiftRowsOutput[18]) );
  XOR2_X1 U370 ( .A(ciphertext[83]), .B(RoundKey[115]), .Z(ShiftRowsOutput[19]) );
  XOR2_X1 U371 ( .A(ciphertext[84]), .B(RoundKey[116]), .Z(ShiftRowsOutput[20]) );
  XOR2_X1 U372 ( .A(ciphertext[85]), .B(RoundKey[117]), .Z(ShiftRowsOutput[21]) );
  XOR2_X1 U373 ( .A(ciphertext[86]), .B(RoundKey[118]), .Z(ShiftRowsOutput[22]) );
  XOR2_X1 U374 ( .A(ciphertext[87]), .B(RoundKey[119]), .Z(ShiftRowsOutput[23]) );
  XOR2_X1 U375 ( .A(ciphertext[75]), .B(KSSubBytesInput[11]), .Z(
        ShiftRowsOutput[75]) );
  XOR2_X1 U376 ( .A(ciphertext[120]), .B(RoundKey[120]), .Z(
        ShiftRowsOutput[120]) );
  XOR2_X1 U377 ( .A(ciphertext[121]), .B(RoundKey[121]), .Z(
        ShiftRowsOutput[121]) );
  XOR2_X1 U378 ( .A(ciphertext[122]), .B(RoundKey[122]), .Z(
        ShiftRowsOutput[122]) );
  XOR2_X1 U379 ( .A(ciphertext[123]), .B(RoundKey[123]), .Z(
        ShiftRowsOutput[123]) );
  XOR2_X1 U380 ( .A(ciphertext[124]), .B(RoundKey[124]), .Z(
        ShiftRowsOutput[124]) );
  XOR2_X1 U381 ( .A(ciphertext[125]), .B(RoundKey[125]), .Z(
        ShiftRowsOutput[125]) );
  XOR2_X1 U382 ( .A(ciphertext[126]), .B(RoundKey[126]), .Z(
        ShiftRowsOutput[126]) );
  XOR2_X1 U383 ( .A(ciphertext[127]), .B(RoundKey[127]), .Z(
        ShiftRowsOutput[127]) );
  XOR2_X1 U384 ( .A(ciphertext[76]), .B(KSSubBytesInput[12]), .Z(
        ShiftRowsOutput[76]) );
  XOR2_X1 U385 ( .A(ciphertext[77]), .B(KSSubBytesInput[13]), .Z(
        ShiftRowsOutput[77]) );
  XOR2_X1 U386 ( .A(ciphertext[78]), .B(KSSubBytesInput[14]), .Z(
        ShiftRowsOutput[78]) );
  XOR2_X1 U387 ( .A(ciphertext[79]), .B(KSSubBytesInput[15]), .Z(
        ShiftRowsOutput[79]) );
  XOR2_X1 U388 ( .A(ciphertext[112]), .B(KSSubBytesInput[0]), .Z(
        ShiftRowsOutput[48]) );
  XOR2_X1 U389 ( .A(ciphertext[113]), .B(KSSubBytesInput[1]), .Z(
        ShiftRowsOutput[49]) );
  XOR2_X1 U390 ( .A(ciphertext[114]), .B(KSSubBytesInput[2]), .Z(
        ShiftRowsOutput[50]) );
  XOR2_X1 U391 ( .A(ciphertext[115]), .B(KSSubBytesInput[3]), .Z(
        ShiftRowsOutput[51]) );
  XOR2_X1 U392 ( .A(ciphertext[33]), .B(KSSubBytesInput[17]), .Z(
        ShiftRowsOutput[97]) );
  XOR2_X1 U393 ( .A(ciphertext[116]), .B(KSSubBytesInput[4]), .Z(
        ShiftRowsOutput[52]) );
  XOR2_X1 U394 ( .A(ciphertext[117]), .B(KSSubBytesInput[5]), .Z(
        ShiftRowsOutput[53]) );
  XOR2_X1 U395 ( .A(ciphertext[118]), .B(KSSubBytesInput[6]), .Z(
        ShiftRowsOutput[54]) );
  XOR2_X1 U396 ( .A(ciphertext[119]), .B(KSSubBytesInput[7]), .Z(
        ShiftRowsOutput[55]) );
  XOR2_X1 U397 ( .A(ciphertext[24]), .B(KSSubBytesInput[24]), .Z(
        ShiftRowsOutput[24]) );
  XOR2_X1 U398 ( .A(ciphertext[25]), .B(KSSubBytesInput[25]), .Z(
        ShiftRowsOutput[25]) );
  XOR2_X1 U399 ( .A(ciphertext[26]), .B(KSSubBytesInput[26]), .Z(
        ShiftRowsOutput[26]) );
  XOR2_X1 U400 ( .A(ciphertext[27]), .B(KSSubBytesInput[27]), .Z(
        ShiftRowsOutput[27]) );
  XOR2_X1 U401 ( .A(ciphertext[28]), .B(KSSubBytesInput[28]), .Z(
        ShiftRowsOutput[28]) );
  XOR2_X1 U402 ( .A(ciphertext[29]), .B(KSSubBytesInput[29]), .Z(
        ShiftRowsOutput[29]) );
  XOR2_X1 U403 ( .A(ciphertext[34]), .B(KSSubBytesInput[18]), .Z(
        ShiftRowsOutput[98]) );
  XOR2_X1 U404 ( .A(ciphertext[30]), .B(KSSubBytesInput[30]), .Z(
        ShiftRowsOutput[30]) );
  XOR2_X1 U405 ( .A(ciphertext[31]), .B(KSSubBytesInput[31]), .Z(
        ShiftRowsOutput[31]) );
  XOR2_X1 U406 ( .A(ciphertext[64]), .B(RoundKey[32]), .Z(ShiftRowsOutput[0])
         );
  XOR2_X1 U407 ( .A(ciphertext[65]), .B(RoundKey[33]), .Z(ShiftRowsOutput[1])
         );
  XOR2_X1 U408 ( .A(ciphertext[66]), .B(RoundKey[34]), .Z(ShiftRowsOutput[2])
         );
  XOR2_X1 U409 ( .A(ciphertext[67]), .B(RoundKey[35]), .Z(ShiftRowsOutput[3])
         );
  XOR2_X1 U410 ( .A(ciphertext[68]), .B(RoundKey[36]), .Z(ShiftRowsOutput[4])
         );
  XOR2_X1 U411 ( .A(ciphertext[69]), .B(RoundKey[37]), .Z(ShiftRowsOutput[5])
         );
  XOR2_X1 U412 ( .A(ciphertext[70]), .B(RoundKey[38]), .Z(ShiftRowsOutput[6])
         );
  XOR2_X1 U413 ( .A(ciphertext[71]), .B(RoundKey[39]), .Z(ShiftRowsOutput[7])
         );
  XOR2_X1 U414 ( .A(ciphertext[35]), .B(KSSubBytesInput[19]), .Z(
        ShiftRowsOutput[99]) );
  XOR2_X1 U415 ( .A(ciphertext[104]), .B(RoundKey[40]), .Z(
        ShiftRowsOutput[104]) );
  XOR2_X1 U416 ( .A(ciphertext[105]), .B(RoundKey[41]), .Z(
        ShiftRowsOutput[105]) );
  XOR2_X1 U417 ( .A(ciphertext[106]), .B(RoundKey[42]), .Z(
        ShiftRowsOutput[106]) );
  XOR2_X1 U418 ( .A(ciphertext[107]), .B(RoundKey[43]), .Z(
        ShiftRowsOutput[107]) );
  XOR2_X1 U419 ( .A(ciphertext[108]), .B(RoundKey[44]), .Z(
        ShiftRowsOutput[108]) );
  XOR2_X1 U420 ( .A(ciphertext[109]), .B(RoundKey[45]), .Z(
        ShiftRowsOutput[109]) );
  XOR2_X1 U421 ( .A(ciphertext[110]), .B(RoundKey[46]), .Z(
        ShiftRowsOutput[110]) );
  XOR2_X1 U422 ( .A(ciphertext[111]), .B(RoundKey[47]), .Z(
        ShiftRowsOutput[111]) );
  XOR2_X1 U423 ( .A(ciphertext[16]), .B(RoundKey[48]), .Z(ShiftRowsOutput[80])
         );
  XOR2_X1 U424 ( .A(ciphertext[17]), .B(RoundKey[49]), .Z(ShiftRowsOutput[81])
         );
  XOR2_X1 U425 ( .A(ciphertext[36]), .B(KSSubBytesInput[20]), .Z(
        ShiftRowsOutput[100]) );
  XOR2_X1 U426 ( .A(ciphertext[18]), .B(RoundKey[50]), .Z(ShiftRowsOutput[82])
         );
  XOR2_X1 U427 ( .A(ciphertext[19]), .B(RoundKey[51]), .Z(ShiftRowsOutput[83])
         );
  XOR2_X1 U428 ( .A(ciphertext[20]), .B(RoundKey[52]), .Z(ShiftRowsOutput[84])
         );
  XOR2_X1 U429 ( .A(ciphertext[21]), .B(RoundKey[53]), .Z(ShiftRowsOutput[85])
         );
  XOR2_X1 U430 ( .A(ciphertext[22]), .B(RoundKey[54]), .Z(ShiftRowsOutput[86])
         );
  XOR2_X1 U431 ( .A(ciphertext[23]), .B(RoundKey[55]), .Z(ShiftRowsOutput[87])
         );
  XOR2_X1 U432 ( .A(ciphertext[56]), .B(RoundKey[56]), .Z(ShiftRowsOutput[56])
         );
  XOR2_X1 U433 ( .A(ciphertext[57]), .B(RoundKey[57]), .Z(ShiftRowsOutput[57])
         );
  XOR2_X1 U434 ( .A(ciphertext[58]), .B(RoundKey[58]), .Z(ShiftRowsOutput[58])
         );
  XOR2_X1 U435 ( .A(ciphertext[59]), .B(RoundKey[59]), .Z(ShiftRowsOutput[59])
         );
  XOR2_X1 U436 ( .A(ciphertext[37]), .B(KSSubBytesInput[21]), .Z(
        ShiftRowsOutput[101]) );
  XOR2_X1 U437 ( .A(ciphertext[60]), .B(RoundKey[60]), .Z(ShiftRowsOutput[60])
         );
  XOR2_X1 U438 ( .A(ciphertext[61]), .B(RoundKey[61]), .Z(ShiftRowsOutput[61])
         );
  XOR2_X1 U439 ( .A(ciphertext[62]), .B(RoundKey[62]), .Z(ShiftRowsOutput[62])
         );
  XOR2_X1 U440 ( .A(ciphertext[63]), .B(RoundKey[63]), .Z(ShiftRowsOutput[63])
         );
  XOR2_X1 U441 ( .A(ciphertext[96]), .B(RoundKey[64]), .Z(ShiftRowsOutput[32])
         );
  XOR2_X1 U442 ( .A(ciphertext[97]), .B(RoundKey[65]), .Z(ShiftRowsOutput[33])
         );
  XOR2_X1 U443 ( .A(ciphertext[98]), .B(RoundKey[66]), .Z(ShiftRowsOutput[34])
         );
  XOR2_X1 U444 ( .A(ciphertext[99]), .B(RoundKey[67]), .Z(ShiftRowsOutput[35])
         );
  XOR2_X1 U445 ( .A(ciphertext[100]), .B(RoundKey[68]), .Z(ShiftRowsOutput[36]) );
  XOR2_X1 U446 ( .A(ciphertext[101]), .B(RoundKey[69]), .Z(ShiftRowsOutput[37]) );
  XOR2_X1 U447 ( .A(ciphertext[38]), .B(KSSubBytesInput[22]), .Z(
        ShiftRowsOutput[102]) );
  XOR2_X1 U448 ( .A(ciphertext[102]), .B(RoundKey[70]), .Z(ShiftRowsOutput[38]) );
  XOR2_X1 U449 ( .A(ciphertext[103]), .B(RoundKey[71]), .Z(ShiftRowsOutput[39]) );
  XOR2_X1 U450 ( .A(ciphertext[8]), .B(RoundKey[72]), .Z(ShiftRowsOutput[8])
         );
  XOR2_X1 U451 ( .A(ciphertext[9]), .B(RoundKey[73]), .Z(ShiftRowsOutput[9])
         );
  XOR2_X1 U452 ( .A(ciphertext[10]), .B(RoundKey[74]), .Z(ShiftRowsOutput[10])
         );
  XOR2_X1 U453 ( .A(ciphertext[11]), .B(RoundKey[75]), .Z(ShiftRowsOutput[11])
         );
  XOR2_X1 U454 ( .A(ciphertext[12]), .B(RoundKey[76]), .Z(ShiftRowsOutput[12])
         );
  XOR2_X1 U455 ( .A(ciphertext[13]), .B(RoundKey[77]), .Z(ShiftRowsOutput[13])
         );
  XOR2_X1 U456 ( .A(ciphertext[14]), .B(RoundKey[78]), .Z(ShiftRowsOutput[14])
         );
  XOR2_X1 U457 ( .A(ciphertext[15]), .B(RoundKey[79]), .Z(ShiftRowsOutput[15])
         );
  XOR2_X1 U458 ( .A(ciphertext[39]), .B(KSSubBytesInput[23]), .Z(
        ShiftRowsOutput[103]) );
  XOR2_X1 U459 ( .A(ciphertext[48]), .B(RoundKey[80]), .Z(ShiftRowsOutput[112]) );
  XOR2_X1 U460 ( .A(ciphertext[49]), .B(RoundKey[81]), .Z(ShiftRowsOutput[113]) );
  XOR2_X1 U461 ( .A(ciphertext[50]), .B(RoundKey[82]), .Z(ShiftRowsOutput[114]) );
  XOR2_X1 U462 ( .A(ciphertext[51]), .B(RoundKey[83]), .Z(ShiftRowsOutput[115]) );
  XOR2_X1 U463 ( .A(ciphertext[52]), .B(RoundKey[84]), .Z(ShiftRowsOutput[116]) );
  XOR2_X1 U464 ( .A(ciphertext[53]), .B(RoundKey[85]), .Z(ShiftRowsOutput[117]) );
  XOR2_X1 U465 ( .A(ciphertext[54]), .B(RoundKey[86]), .Z(ShiftRowsOutput[118]) );
  XOR2_X1 U466 ( .A(ciphertext[55]), .B(RoundKey[87]), .Z(ShiftRowsOutput[119]) );
  XOR2_X1 U467 ( .A(ciphertext[88]), .B(RoundKey[88]), .Z(ShiftRowsOutput[88])
         );
  XOR2_X1 U468 ( .A(ciphertext[89]), .B(RoundKey[89]), .Z(ShiftRowsOutput[89])
         );
  XOR2_X1 U469 ( .A(ciphertext[72]), .B(KSSubBytesInput[8]), .Z(
        ShiftRowsOutput[72]) );
  XOR2_X1 U470 ( .A(ciphertext[90]), .B(RoundKey[90]), .Z(ShiftRowsOutput[90])
         );
  XOR2_X1 U471 ( .A(ciphertext[91]), .B(RoundKey[91]), .Z(ShiftRowsOutput[91])
         );
  XOR2_X1 U472 ( .A(ciphertext[92]), .B(RoundKey[92]), .Z(ShiftRowsOutput[92])
         );
  XOR2_X1 U473 ( .A(ciphertext[93]), .B(RoundKey[93]), .Z(ShiftRowsOutput[93])
         );
  XOR2_X1 U474 ( .A(ciphertext[94]), .B(RoundKey[94]), .Z(ShiftRowsOutput[94])
         );
  XOR2_X1 U475 ( .A(ciphertext[95]), .B(RoundKey[95]), .Z(ShiftRowsOutput[95])
         );
  XOR2_X1 U476 ( .A(ciphertext[0]), .B(RoundKey[96]), .Z(ShiftRowsOutput[64])
         );
  XOR2_X1 U477 ( .A(ciphertext[1]), .B(RoundKey[97]), .Z(ShiftRowsOutput[65])
         );
  XOR2_X1 U478 ( .A(ciphertext[2]), .B(RoundKey[98]), .Z(ShiftRowsOutput[66])
         );
  XOR2_X1 U479 ( .A(ciphertext[3]), .B(RoundKey[99]), .Z(ShiftRowsOutput[67])
         );
  XOR2_X1 U480 ( .A(ciphertext[73]), .B(KSSubBytesInput[9]), .Z(
        ShiftRowsOutput[73]) );
  INV_X1 RoundReg_Inst_ff_SDE_0_current_state_reg_U1 ( .A(ciphertext[32]), 
        .ZN(RoundReg_Inst_ff_SDE_0_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_0_next_state), .CK(clk), .Q(ciphertext[32]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_0_MUX_inst_U1 ( .A(RoundOutput[0]), .B(
        plaintext[0]), .S(reset), .Z(RoundReg_Inst_ff_SDE_0_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_1_current_state_reg_U1 ( .A(ciphertext[33]), 
        .ZN(RoundReg_Inst_ff_SDE_1_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_1_next_state), .CK(clk), .Q(ciphertext[33]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_1_MUX_inst_U1 ( .A(RoundOutput[1]), .B(
        plaintext[1]), .S(reset), .Z(RoundReg_Inst_ff_SDE_1_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_2_current_state_reg_U1 ( .A(ciphertext[34]), 
        .ZN(RoundReg_Inst_ff_SDE_2_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_2_next_state), .CK(clk), .Q(ciphertext[34]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_2_MUX_inst_U1 ( .A(RoundOutput[2]), .B(
        plaintext[2]), .S(reset), .Z(RoundReg_Inst_ff_SDE_2_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_3_current_state_reg_U1 ( .A(ciphertext[35]), 
        .ZN(RoundReg_Inst_ff_SDE_3_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_3_next_state), .CK(clk), .Q(ciphertext[35]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_3_MUX_inst_U1 ( .A(RoundOutput[3]), .B(
        plaintext[3]), .S(reset), .Z(RoundReg_Inst_ff_SDE_3_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_4_current_state_reg_U1 ( .A(ciphertext[36]), 
        .ZN(RoundReg_Inst_ff_SDE_4_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_4_next_state), .CK(clk), .Q(ciphertext[36]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_4_MUX_inst_U1 ( .A(RoundOutput[4]), .B(
        plaintext[4]), .S(reset), .Z(RoundReg_Inst_ff_SDE_4_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_5_current_state_reg_U1 ( .A(ciphertext[37]), 
        .ZN(RoundReg_Inst_ff_SDE_5_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_5_next_state), .CK(clk), .Q(ciphertext[37]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_5_MUX_inst_U1 ( .A(RoundOutput[5]), .B(
        plaintext[5]), .S(reset), .Z(RoundReg_Inst_ff_SDE_5_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_6_current_state_reg_U1 ( .A(ciphertext[38]), 
        .ZN(RoundReg_Inst_ff_SDE_6_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_6_next_state), .CK(clk), .Q(ciphertext[38]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_6_MUX_inst_U1 ( .A(RoundOutput[6]), .B(
        plaintext[6]), .S(reset), .Z(RoundReg_Inst_ff_SDE_6_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_7_current_state_reg_U1 ( .A(ciphertext[39]), 
        .ZN(RoundReg_Inst_ff_SDE_7_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_7_next_state), .CK(clk), .Q(ciphertext[39]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_7_MUX_inst_U1 ( .A(RoundOutput[7]), .B(
        plaintext[7]), .S(reset), .Z(RoundReg_Inst_ff_SDE_7_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_8_current_state_reg_U1 ( .A(ciphertext[72]), 
        .ZN(RoundReg_Inst_ff_SDE_8_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_8_next_state), .CK(clk), .Q(ciphertext[72]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_8_MUX_inst_U1 ( .A(RoundOutput[8]), .B(
        plaintext[8]), .S(reset), .Z(RoundReg_Inst_ff_SDE_8_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_9_current_state_reg_U1 ( .A(ciphertext[73]), 
        .ZN(RoundReg_Inst_ff_SDE_9_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_9_next_state), .CK(clk), .Q(ciphertext[73]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_9_MUX_inst_U1 ( .A(RoundOutput[9]), .B(
        plaintext[9]), .S(reset), .Z(RoundReg_Inst_ff_SDE_9_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_10_current_state_reg_U1 ( .A(ciphertext[74]), 
        .ZN(RoundReg_Inst_ff_SDE_10_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_10_next_state), .CK(clk), .Q(ciphertext[74]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_10_MUX_inst_U1 ( .A(RoundOutput[10]), .B(
        plaintext[10]), .S(reset), .Z(RoundReg_Inst_ff_SDE_10_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_11_current_state_reg_U1 ( .A(ciphertext[75]), 
        .ZN(RoundReg_Inst_ff_SDE_11_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_11_next_state), .CK(clk), .Q(ciphertext[75]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_11_MUX_inst_U1 ( .A(RoundOutput[11]), .B(
        plaintext[11]), .S(reset), .Z(RoundReg_Inst_ff_SDE_11_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_12_current_state_reg_U1 ( .A(ciphertext[76]), 
        .ZN(RoundReg_Inst_ff_SDE_12_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_12_next_state), .CK(clk), .Q(ciphertext[76]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_12_MUX_inst_U1 ( .A(RoundOutput[12]), .B(
        plaintext[12]), .S(reset), .Z(RoundReg_Inst_ff_SDE_12_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_13_current_state_reg_U1 ( .A(ciphertext[77]), 
        .ZN(RoundReg_Inst_ff_SDE_13_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_13_next_state), .CK(clk), .Q(ciphertext[77]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_13_MUX_inst_U1 ( .A(RoundOutput[13]), .B(
        plaintext[13]), .S(reset), .Z(RoundReg_Inst_ff_SDE_13_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_14_current_state_reg_U1 ( .A(ciphertext[78]), 
        .ZN(RoundReg_Inst_ff_SDE_14_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_14_next_state), .CK(clk), .Q(ciphertext[78]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_14_MUX_inst_U1 ( .A(RoundOutput[14]), .B(
        plaintext[14]), .S(reset), .Z(RoundReg_Inst_ff_SDE_14_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_15_current_state_reg_U1 ( .A(ciphertext[79]), 
        .ZN(RoundReg_Inst_ff_SDE_15_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_15_next_state), .CK(clk), .Q(ciphertext[79]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_15_MUX_inst_U1 ( .A(RoundOutput[15]), .B(
        plaintext[15]), .S(reset), .Z(RoundReg_Inst_ff_SDE_15_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_16_current_state_reg_U1 ( .A(ciphertext[112]), 
        .ZN(RoundReg_Inst_ff_SDE_16_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_16_next_state), .CK(clk), .Q(ciphertext[112]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_16_MUX_inst_U1 ( .A(RoundOutput[16]), .B(
        plaintext[16]), .S(reset), .Z(RoundReg_Inst_ff_SDE_16_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_17_current_state_reg_U1 ( .A(ciphertext[113]), 
        .ZN(RoundReg_Inst_ff_SDE_17_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_17_next_state), .CK(clk), .Q(ciphertext[113]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_17_MUX_inst_U1 ( .A(RoundOutput[17]), .B(
        plaintext[17]), .S(reset), .Z(RoundReg_Inst_ff_SDE_17_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_18_current_state_reg_U1 ( .A(ciphertext[114]), 
        .ZN(RoundReg_Inst_ff_SDE_18_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_18_next_state), .CK(clk), .Q(ciphertext[114]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_18_MUX_inst_U1 ( .A(RoundOutput[18]), .B(
        plaintext[18]), .S(reset), .Z(RoundReg_Inst_ff_SDE_18_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_19_current_state_reg_U1 ( .A(ciphertext[115]), 
        .ZN(RoundReg_Inst_ff_SDE_19_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_19_next_state), .CK(clk), .Q(ciphertext[115]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_19_MUX_inst_U1 ( .A(RoundOutput[19]), .B(
        plaintext[19]), .S(reset), .Z(RoundReg_Inst_ff_SDE_19_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_20_current_state_reg_U1 ( .A(ciphertext[116]), 
        .ZN(RoundReg_Inst_ff_SDE_20_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_20_next_state), .CK(clk), .Q(ciphertext[116]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_20_MUX_inst_U1 ( .A(RoundOutput[20]), .B(
        plaintext[20]), .S(reset), .Z(RoundReg_Inst_ff_SDE_20_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_21_current_state_reg_U1 ( .A(ciphertext[117]), 
        .ZN(RoundReg_Inst_ff_SDE_21_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_21_next_state), .CK(clk), .Q(ciphertext[117]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_21_MUX_inst_U1 ( .A(RoundOutput[21]), .B(
        plaintext[21]), .S(reset), .Z(RoundReg_Inst_ff_SDE_21_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_22_current_state_reg_U1 ( .A(ciphertext[118]), 
        .ZN(RoundReg_Inst_ff_SDE_22_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_22_next_state), .CK(clk), .Q(ciphertext[118]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_22_MUX_inst_U1 ( .A(RoundOutput[22]), .B(
        plaintext[22]), .S(reset), .Z(RoundReg_Inst_ff_SDE_22_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_23_current_state_reg_U1 ( .A(ciphertext[119]), 
        .ZN(RoundReg_Inst_ff_SDE_23_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_23_next_state), .CK(clk), .Q(ciphertext[119]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_23_MUX_inst_U1 ( .A(RoundOutput[23]), .B(
        plaintext[23]), .S(reset), .Z(RoundReg_Inst_ff_SDE_23_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_24_current_state_reg_U1 ( .A(ciphertext[24]), 
        .ZN(RoundReg_Inst_ff_SDE_24_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_24_next_state), .CK(clk), .Q(ciphertext[24]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_24_MUX_inst_U1 ( .A(RoundOutput[24]), .B(
        plaintext[24]), .S(reset), .Z(RoundReg_Inst_ff_SDE_24_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_25_current_state_reg_U1 ( .A(ciphertext[25]), 
        .ZN(RoundReg_Inst_ff_SDE_25_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_25_next_state), .CK(clk), .Q(ciphertext[25]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_25_MUX_inst_U1 ( .A(RoundOutput[25]), .B(
        plaintext[25]), .S(reset), .Z(RoundReg_Inst_ff_SDE_25_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_26_current_state_reg_U1 ( .A(ciphertext[26]), 
        .ZN(RoundReg_Inst_ff_SDE_26_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_26_next_state), .CK(clk), .Q(ciphertext[26]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_26_MUX_inst_U1 ( .A(RoundOutput[26]), .B(
        plaintext[26]), .S(reset), .Z(RoundReg_Inst_ff_SDE_26_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_27_current_state_reg_U1 ( .A(ciphertext[27]), 
        .ZN(RoundReg_Inst_ff_SDE_27_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_27_next_state), .CK(clk), .Q(ciphertext[27]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_27_MUX_inst_U1 ( .A(RoundOutput[27]), .B(
        plaintext[27]), .S(reset), .Z(RoundReg_Inst_ff_SDE_27_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_28_current_state_reg_U1 ( .A(ciphertext[28]), 
        .ZN(RoundReg_Inst_ff_SDE_28_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_28_next_state), .CK(clk), .Q(ciphertext[28]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_28_MUX_inst_U1 ( .A(RoundOutput[28]), .B(
        plaintext[28]), .S(reset), .Z(RoundReg_Inst_ff_SDE_28_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_29_current_state_reg_U1 ( .A(ciphertext[29]), 
        .ZN(RoundReg_Inst_ff_SDE_29_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_29_next_state), .CK(clk), .Q(ciphertext[29]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_29_MUX_inst_U1 ( .A(RoundOutput[29]), .B(
        plaintext[29]), .S(reset), .Z(RoundReg_Inst_ff_SDE_29_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_30_current_state_reg_U1 ( .A(ciphertext[30]), 
        .ZN(RoundReg_Inst_ff_SDE_30_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_30_next_state), .CK(clk), .Q(ciphertext[30]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_30_MUX_inst_U1 ( .A(RoundOutput[30]), .B(
        plaintext[30]), .S(reset), .Z(RoundReg_Inst_ff_SDE_30_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_31_current_state_reg_U1 ( .A(ciphertext[31]), 
        .ZN(RoundReg_Inst_ff_SDE_31_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_31_next_state), .CK(clk), .Q(ciphertext[31]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_31_MUX_inst_U1 ( .A(RoundOutput[31]), .B(
        plaintext[31]), .S(reset), .Z(RoundReg_Inst_ff_SDE_31_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_32_current_state_reg_U1 ( .A(ciphertext[64]), 
        .ZN(RoundReg_Inst_ff_SDE_32_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_32_next_state), .CK(clk), .Q(ciphertext[64]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_32_MUX_inst_U1 ( .A(RoundOutput[32]), .B(
        plaintext[32]), .S(reset), .Z(RoundReg_Inst_ff_SDE_32_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_33_current_state_reg_U1 ( .A(ciphertext[65]), 
        .ZN(RoundReg_Inst_ff_SDE_33_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_33_next_state), .CK(clk), .Q(ciphertext[65]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_33_MUX_inst_U1 ( .A(RoundOutput[33]), .B(
        plaintext[33]), .S(reset), .Z(RoundReg_Inst_ff_SDE_33_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_34_current_state_reg_U1 ( .A(ciphertext[66]), 
        .ZN(RoundReg_Inst_ff_SDE_34_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_34_next_state), .CK(clk), .Q(ciphertext[66]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_34_MUX_inst_U1 ( .A(RoundOutput[34]), .B(
        plaintext[34]), .S(reset), .Z(RoundReg_Inst_ff_SDE_34_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_35_current_state_reg_U1 ( .A(ciphertext[67]), 
        .ZN(RoundReg_Inst_ff_SDE_35_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_35_next_state), .CK(clk), .Q(ciphertext[67]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_35_MUX_inst_U1 ( .A(RoundOutput[35]), .B(
        plaintext[35]), .S(reset), .Z(RoundReg_Inst_ff_SDE_35_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_36_current_state_reg_U1 ( .A(ciphertext[68]), 
        .ZN(RoundReg_Inst_ff_SDE_36_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_36_next_state), .CK(clk), .Q(ciphertext[68]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_36_MUX_inst_U1 ( .A(RoundOutput[36]), .B(
        plaintext[36]), .S(reset), .Z(RoundReg_Inst_ff_SDE_36_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_37_current_state_reg_U1 ( .A(ciphertext[69]), 
        .ZN(RoundReg_Inst_ff_SDE_37_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_37_next_state), .CK(clk), .Q(ciphertext[69]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_37_MUX_inst_U1 ( .A(RoundOutput[37]), .B(
        plaintext[37]), .S(reset), .Z(RoundReg_Inst_ff_SDE_37_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_38_current_state_reg_U1 ( .A(ciphertext[70]), 
        .ZN(RoundReg_Inst_ff_SDE_38_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_38_next_state), .CK(clk), .Q(ciphertext[70]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_38_MUX_inst_U1 ( .A(RoundOutput[38]), .B(
        plaintext[38]), .S(reset), .Z(RoundReg_Inst_ff_SDE_38_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_39_current_state_reg_U1 ( .A(ciphertext[71]), 
        .ZN(RoundReg_Inst_ff_SDE_39_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_39_next_state), .CK(clk), .Q(ciphertext[71]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_39_MUX_inst_U1 ( .A(RoundOutput[39]), .B(
        plaintext[39]), .S(reset), .Z(RoundReg_Inst_ff_SDE_39_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_40_current_state_reg_U1 ( .A(ciphertext[104]), 
        .ZN(RoundReg_Inst_ff_SDE_40_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_40_next_state), .CK(clk), .Q(ciphertext[104]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_40_MUX_inst_U1 ( .A(RoundOutput[40]), .B(
        plaintext[40]), .S(reset), .Z(RoundReg_Inst_ff_SDE_40_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_41_current_state_reg_U1 ( .A(ciphertext[105]), 
        .ZN(RoundReg_Inst_ff_SDE_41_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_41_next_state), .CK(clk), .Q(ciphertext[105]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_41_MUX_inst_U1 ( .A(RoundOutput[41]), .B(
        plaintext[41]), .S(reset), .Z(RoundReg_Inst_ff_SDE_41_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_42_current_state_reg_U1 ( .A(ciphertext[106]), 
        .ZN(RoundReg_Inst_ff_SDE_42_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_42_next_state), .CK(clk), .Q(ciphertext[106]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_42_MUX_inst_U1 ( .A(RoundOutput[42]), .B(
        plaintext[42]), .S(reset), .Z(RoundReg_Inst_ff_SDE_42_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_43_current_state_reg_U1 ( .A(ciphertext[107]), 
        .ZN(RoundReg_Inst_ff_SDE_43_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_43_next_state), .CK(clk), .Q(ciphertext[107]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_43_MUX_inst_U1 ( .A(RoundOutput[43]), .B(
        plaintext[43]), .S(reset), .Z(RoundReg_Inst_ff_SDE_43_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_44_current_state_reg_U1 ( .A(ciphertext[108]), 
        .ZN(RoundReg_Inst_ff_SDE_44_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_44_next_state), .CK(clk), .Q(ciphertext[108]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_44_MUX_inst_U1 ( .A(RoundOutput[44]), .B(
        plaintext[44]), .S(reset), .Z(RoundReg_Inst_ff_SDE_44_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_45_current_state_reg_U1 ( .A(ciphertext[109]), 
        .ZN(RoundReg_Inst_ff_SDE_45_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_45_next_state), .CK(clk), .Q(ciphertext[109]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_45_MUX_inst_U1 ( .A(RoundOutput[45]), .B(
        plaintext[45]), .S(reset), .Z(RoundReg_Inst_ff_SDE_45_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_46_current_state_reg_U1 ( .A(ciphertext[110]), 
        .ZN(RoundReg_Inst_ff_SDE_46_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_46_next_state), .CK(clk), .Q(ciphertext[110]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_46_MUX_inst_U1 ( .A(RoundOutput[46]), .B(
        plaintext[46]), .S(reset), .Z(RoundReg_Inst_ff_SDE_46_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_47_current_state_reg_U1 ( .A(ciphertext[111]), 
        .ZN(RoundReg_Inst_ff_SDE_47_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_47_next_state), .CK(clk), .Q(ciphertext[111]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_47_MUX_inst_U1 ( .A(RoundOutput[47]), .B(
        plaintext[47]), .S(reset), .Z(RoundReg_Inst_ff_SDE_47_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_48_current_state_reg_U1 ( .A(ciphertext[16]), 
        .ZN(RoundReg_Inst_ff_SDE_48_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_48_next_state), .CK(clk), .Q(ciphertext[16]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_48_MUX_inst_U1 ( .A(RoundOutput[48]), .B(
        plaintext[48]), .S(reset), .Z(RoundReg_Inst_ff_SDE_48_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_49_current_state_reg_U1 ( .A(ciphertext[17]), 
        .ZN(RoundReg_Inst_ff_SDE_49_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_49_next_state), .CK(clk), .Q(ciphertext[17]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_49_MUX_inst_U1 ( .A(RoundOutput[49]), .B(
        plaintext[49]), .S(reset), .Z(RoundReg_Inst_ff_SDE_49_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_50_current_state_reg_U1 ( .A(ciphertext[18]), 
        .ZN(RoundReg_Inst_ff_SDE_50_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_50_next_state), .CK(clk), .Q(ciphertext[18]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_50_MUX_inst_U1 ( .A(RoundOutput[50]), .B(
        plaintext[50]), .S(reset), .Z(RoundReg_Inst_ff_SDE_50_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_51_current_state_reg_U1 ( .A(ciphertext[19]), 
        .ZN(RoundReg_Inst_ff_SDE_51_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_51_next_state), .CK(clk), .Q(ciphertext[19]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_51_MUX_inst_U1 ( .A(RoundOutput[51]), .B(
        plaintext[51]), .S(reset), .Z(RoundReg_Inst_ff_SDE_51_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_52_current_state_reg_U1 ( .A(ciphertext[20]), 
        .ZN(RoundReg_Inst_ff_SDE_52_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_52_next_state), .CK(clk), .Q(ciphertext[20]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_52_MUX_inst_U1 ( .A(RoundOutput[52]), .B(
        plaintext[52]), .S(reset), .Z(RoundReg_Inst_ff_SDE_52_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_53_current_state_reg_U1 ( .A(ciphertext[21]), 
        .ZN(RoundReg_Inst_ff_SDE_53_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_53_next_state), .CK(clk), .Q(ciphertext[21]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_53_MUX_inst_U1 ( .A(RoundOutput[53]), .B(
        plaintext[53]), .S(reset), .Z(RoundReg_Inst_ff_SDE_53_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_54_current_state_reg_U1 ( .A(ciphertext[22]), 
        .ZN(RoundReg_Inst_ff_SDE_54_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_54_next_state), .CK(clk), .Q(ciphertext[22]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_54_MUX_inst_U1 ( .A(RoundOutput[54]), .B(
        plaintext[54]), .S(reset), .Z(RoundReg_Inst_ff_SDE_54_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_55_current_state_reg_U1 ( .A(ciphertext[23]), 
        .ZN(RoundReg_Inst_ff_SDE_55_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_55_next_state), .CK(clk), .Q(ciphertext[23]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_55_MUX_inst_U1 ( .A(RoundOutput[55]), .B(
        plaintext[55]), .S(reset), .Z(RoundReg_Inst_ff_SDE_55_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_56_current_state_reg_U1 ( .A(ciphertext[56]), 
        .ZN(RoundReg_Inst_ff_SDE_56_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_56_next_state), .CK(clk), .Q(ciphertext[56]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_56_MUX_inst_U1 ( .A(RoundOutput[56]), .B(
        plaintext[56]), .S(reset), .Z(RoundReg_Inst_ff_SDE_56_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_57_current_state_reg_U1 ( .A(ciphertext[57]), 
        .ZN(RoundReg_Inst_ff_SDE_57_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_57_next_state), .CK(clk), .Q(ciphertext[57]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_57_MUX_inst_U1 ( .A(RoundOutput[57]), .B(
        plaintext[57]), .S(reset), .Z(RoundReg_Inst_ff_SDE_57_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_58_current_state_reg_U1 ( .A(ciphertext[58]), 
        .ZN(RoundReg_Inst_ff_SDE_58_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_58_next_state), .CK(clk), .Q(ciphertext[58]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_58_MUX_inst_U1 ( .A(RoundOutput[58]), .B(
        plaintext[58]), .S(reset), .Z(RoundReg_Inst_ff_SDE_58_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_59_current_state_reg_U1 ( .A(ciphertext[59]), 
        .ZN(RoundReg_Inst_ff_SDE_59_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_59_next_state), .CK(clk), .Q(ciphertext[59]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_59_MUX_inst_U1 ( .A(RoundOutput[59]), .B(
        plaintext[59]), .S(reset), .Z(RoundReg_Inst_ff_SDE_59_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_60_current_state_reg_U1 ( .A(ciphertext[60]), 
        .ZN(RoundReg_Inst_ff_SDE_60_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_60_next_state), .CK(clk), .Q(ciphertext[60]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_60_MUX_inst_U1 ( .A(RoundOutput[60]), .B(
        plaintext[60]), .S(reset), .Z(RoundReg_Inst_ff_SDE_60_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_61_current_state_reg_U1 ( .A(ciphertext[61]), 
        .ZN(RoundReg_Inst_ff_SDE_61_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_61_next_state), .CK(clk), .Q(ciphertext[61]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_61_MUX_inst_U1 ( .A(RoundOutput[61]), .B(
        plaintext[61]), .S(reset), .Z(RoundReg_Inst_ff_SDE_61_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_62_current_state_reg_U1 ( .A(ciphertext[62]), 
        .ZN(RoundReg_Inst_ff_SDE_62_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_62_next_state), .CK(clk), .Q(ciphertext[62]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_62_MUX_inst_U1 ( .A(RoundOutput[62]), .B(
        plaintext[62]), .S(reset), .Z(RoundReg_Inst_ff_SDE_62_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_63_current_state_reg_U1 ( .A(ciphertext[63]), 
        .ZN(RoundReg_Inst_ff_SDE_63_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_63_next_state), .CK(clk), .Q(ciphertext[63]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_63_MUX_inst_U1 ( .A(RoundOutput[63]), .B(
        plaintext[63]), .S(reset), .Z(RoundReg_Inst_ff_SDE_63_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_64_current_state_reg_U1 ( .A(ciphertext[96]), 
        .ZN(RoundReg_Inst_ff_SDE_64_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_64_next_state), .CK(clk), .Q(ciphertext[96]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_64_MUX_inst_U1 ( .A(RoundOutput[64]), .B(
        plaintext[64]), .S(reset), .Z(RoundReg_Inst_ff_SDE_64_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_65_current_state_reg_U1 ( .A(ciphertext[97]), 
        .ZN(RoundReg_Inst_ff_SDE_65_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_65_next_state), .CK(clk), .Q(ciphertext[97]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_65_MUX_inst_U1 ( .A(RoundOutput[65]), .B(
        plaintext[65]), .S(reset), .Z(RoundReg_Inst_ff_SDE_65_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_66_current_state_reg_U1 ( .A(ciphertext[98]), 
        .ZN(RoundReg_Inst_ff_SDE_66_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_66_next_state), .CK(clk), .Q(ciphertext[98]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_66_MUX_inst_U1 ( .A(RoundOutput[66]), .B(
        plaintext[66]), .S(reset), .Z(RoundReg_Inst_ff_SDE_66_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_67_current_state_reg_U1 ( .A(ciphertext[99]), 
        .ZN(RoundReg_Inst_ff_SDE_67_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_67_next_state), .CK(clk), .Q(ciphertext[99]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_67_MUX_inst_U1 ( .A(RoundOutput[67]), .B(
        plaintext[67]), .S(reset), .Z(RoundReg_Inst_ff_SDE_67_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_68_current_state_reg_U1 ( .A(ciphertext[100]), 
        .ZN(RoundReg_Inst_ff_SDE_68_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_68_next_state), .CK(clk), .Q(ciphertext[100]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_68_MUX_inst_U1 ( .A(RoundOutput[68]), .B(
        plaintext[68]), .S(reset), .Z(RoundReg_Inst_ff_SDE_68_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_69_current_state_reg_U1 ( .A(ciphertext[101]), 
        .ZN(RoundReg_Inst_ff_SDE_69_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_69_next_state), .CK(clk), .Q(ciphertext[101]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_69_MUX_inst_U1 ( .A(RoundOutput[69]), .B(
        plaintext[69]), .S(reset), .Z(RoundReg_Inst_ff_SDE_69_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_70_current_state_reg_U1 ( .A(ciphertext[102]), 
        .ZN(RoundReg_Inst_ff_SDE_70_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_70_next_state), .CK(clk), .Q(ciphertext[102]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_70_MUX_inst_U1 ( .A(RoundOutput[70]), .B(
        plaintext[70]), .S(reset), .Z(RoundReg_Inst_ff_SDE_70_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_71_current_state_reg_U1 ( .A(ciphertext[103]), 
        .ZN(RoundReg_Inst_ff_SDE_71_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_71_next_state), .CK(clk), .Q(ciphertext[103]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_71_MUX_inst_U1 ( .A(RoundOutput[71]), .B(
        plaintext[71]), .S(reset), .Z(RoundReg_Inst_ff_SDE_71_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_72_current_state_reg_U1 ( .A(ciphertext[8]), 
        .ZN(RoundReg_Inst_ff_SDE_72_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_72_next_state), .CK(clk), .Q(ciphertext[8]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_72_MUX_inst_U1 ( .A(RoundOutput[72]), .B(
        plaintext[72]), .S(reset), .Z(RoundReg_Inst_ff_SDE_72_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_73_current_state_reg_U1 ( .A(ciphertext[9]), 
        .ZN(RoundReg_Inst_ff_SDE_73_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_73_next_state), .CK(clk), .Q(ciphertext[9]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_73_MUX_inst_U1 ( .A(RoundOutput[73]), .B(
        plaintext[73]), .S(reset), .Z(RoundReg_Inst_ff_SDE_73_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_74_current_state_reg_U1 ( .A(ciphertext[10]), 
        .ZN(RoundReg_Inst_ff_SDE_74_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_74_next_state), .CK(clk), .Q(ciphertext[10]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_74_MUX_inst_U1 ( .A(RoundOutput[74]), .B(
        plaintext[74]), .S(reset), .Z(RoundReg_Inst_ff_SDE_74_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_75_current_state_reg_U1 ( .A(ciphertext[11]), 
        .ZN(RoundReg_Inst_ff_SDE_75_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_75_next_state), .CK(clk), .Q(ciphertext[11]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_75_MUX_inst_U1 ( .A(RoundOutput[75]), .B(
        plaintext[75]), .S(reset), .Z(RoundReg_Inst_ff_SDE_75_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_76_current_state_reg_U1 ( .A(ciphertext[12]), 
        .ZN(RoundReg_Inst_ff_SDE_76_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_76_next_state), .CK(clk), .Q(ciphertext[12]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_76_MUX_inst_U1 ( .A(RoundOutput[76]), .B(
        plaintext[76]), .S(reset), .Z(RoundReg_Inst_ff_SDE_76_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_77_current_state_reg_U1 ( .A(ciphertext[13]), 
        .ZN(RoundReg_Inst_ff_SDE_77_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_77_next_state), .CK(clk), .Q(ciphertext[13]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_77_MUX_inst_U1 ( .A(RoundOutput[77]), .B(
        plaintext[77]), .S(reset), .Z(RoundReg_Inst_ff_SDE_77_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_78_current_state_reg_U1 ( .A(ciphertext[14]), 
        .ZN(RoundReg_Inst_ff_SDE_78_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_78_next_state), .CK(clk), .Q(ciphertext[14]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_78_MUX_inst_U1 ( .A(RoundOutput[78]), .B(
        plaintext[78]), .S(reset), .Z(RoundReg_Inst_ff_SDE_78_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_79_current_state_reg_U1 ( .A(ciphertext[15]), 
        .ZN(RoundReg_Inst_ff_SDE_79_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_79_next_state), .CK(clk), .Q(ciphertext[15]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_79_MUX_inst_U1 ( .A(RoundOutput[79]), .B(
        plaintext[79]), .S(reset), .Z(RoundReg_Inst_ff_SDE_79_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_80_current_state_reg_U1 ( .A(ciphertext[48]), 
        .ZN(RoundReg_Inst_ff_SDE_80_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_80_next_state), .CK(clk), .Q(ciphertext[48]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_80_MUX_inst_U1 ( .A(RoundOutput[80]), .B(
        plaintext[80]), .S(reset), .Z(RoundReg_Inst_ff_SDE_80_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_81_current_state_reg_U1 ( .A(ciphertext[49]), 
        .ZN(RoundReg_Inst_ff_SDE_81_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_81_next_state), .CK(clk), .Q(ciphertext[49]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_81_MUX_inst_U1 ( .A(RoundOutput[81]), .B(
        plaintext[81]), .S(reset), .Z(RoundReg_Inst_ff_SDE_81_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_82_current_state_reg_U1 ( .A(ciphertext[50]), 
        .ZN(RoundReg_Inst_ff_SDE_82_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_82_next_state), .CK(clk), .Q(ciphertext[50]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_82_MUX_inst_U1 ( .A(RoundOutput[82]), .B(
        plaintext[82]), .S(reset), .Z(RoundReg_Inst_ff_SDE_82_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_83_current_state_reg_U1 ( .A(ciphertext[51]), 
        .ZN(RoundReg_Inst_ff_SDE_83_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_83_next_state), .CK(clk), .Q(ciphertext[51]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_83_MUX_inst_U1 ( .A(RoundOutput[83]), .B(
        plaintext[83]), .S(reset), .Z(RoundReg_Inst_ff_SDE_83_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_84_current_state_reg_U1 ( .A(ciphertext[52]), 
        .ZN(RoundReg_Inst_ff_SDE_84_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_84_next_state), .CK(clk), .Q(ciphertext[52]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_84_MUX_inst_U1 ( .A(RoundOutput[84]), .B(
        plaintext[84]), .S(reset), .Z(RoundReg_Inst_ff_SDE_84_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_85_current_state_reg_U1 ( .A(ciphertext[53]), 
        .ZN(RoundReg_Inst_ff_SDE_85_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_85_next_state), .CK(clk), .Q(ciphertext[53]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_85_MUX_inst_U1 ( .A(RoundOutput[85]), .B(
        plaintext[85]), .S(reset), .Z(RoundReg_Inst_ff_SDE_85_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_86_current_state_reg_U1 ( .A(ciphertext[54]), 
        .ZN(RoundReg_Inst_ff_SDE_86_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_86_next_state), .CK(clk), .Q(ciphertext[54]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_86_MUX_inst_U1 ( .A(RoundOutput[86]), .B(
        plaintext[86]), .S(reset), .Z(RoundReg_Inst_ff_SDE_86_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_87_current_state_reg_U1 ( .A(ciphertext[55]), 
        .ZN(RoundReg_Inst_ff_SDE_87_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_87_next_state), .CK(clk), .Q(ciphertext[55]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_87_MUX_inst_U1 ( .A(RoundOutput[87]), .B(
        plaintext[87]), .S(reset), .Z(RoundReg_Inst_ff_SDE_87_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_88_current_state_reg_U1 ( .A(ciphertext[88]), 
        .ZN(RoundReg_Inst_ff_SDE_88_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_88_next_state), .CK(clk), .Q(ciphertext[88]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_88_MUX_inst_U1 ( .A(RoundOutput[88]), .B(
        plaintext[88]), .S(reset), .Z(RoundReg_Inst_ff_SDE_88_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_89_current_state_reg_U1 ( .A(ciphertext[89]), 
        .ZN(RoundReg_Inst_ff_SDE_89_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_89_next_state), .CK(clk), .Q(ciphertext[89]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_89_MUX_inst_U1 ( .A(RoundOutput[89]), .B(
        plaintext[89]), .S(reset), .Z(RoundReg_Inst_ff_SDE_89_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_90_current_state_reg_U1 ( .A(ciphertext[90]), 
        .ZN(RoundReg_Inst_ff_SDE_90_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_90_next_state), .CK(clk), .Q(ciphertext[90]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_90_MUX_inst_U1 ( .A(RoundOutput[90]), .B(
        plaintext[90]), .S(reset), .Z(RoundReg_Inst_ff_SDE_90_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_91_current_state_reg_U1 ( .A(ciphertext[91]), 
        .ZN(RoundReg_Inst_ff_SDE_91_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_91_next_state), .CK(clk), .Q(ciphertext[91]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_91_MUX_inst_U1 ( .A(RoundOutput[91]), .B(
        plaintext[91]), .S(reset), .Z(RoundReg_Inst_ff_SDE_91_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_92_current_state_reg_U1 ( .A(ciphertext[92]), 
        .ZN(RoundReg_Inst_ff_SDE_92_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_92_next_state), .CK(clk), .Q(ciphertext[92]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_92_MUX_inst_U1 ( .A(RoundOutput[92]), .B(
        plaintext[92]), .S(reset), .Z(RoundReg_Inst_ff_SDE_92_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_93_current_state_reg_U1 ( .A(ciphertext[93]), 
        .ZN(RoundReg_Inst_ff_SDE_93_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_93_next_state), .CK(clk), .Q(ciphertext[93]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_93_MUX_inst_U1 ( .A(RoundOutput[93]), .B(
        plaintext[93]), .S(reset), .Z(RoundReg_Inst_ff_SDE_93_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_94_current_state_reg_U1 ( .A(ciphertext[94]), 
        .ZN(RoundReg_Inst_ff_SDE_94_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_94_next_state), .CK(clk), .Q(ciphertext[94]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_94_MUX_inst_U1 ( .A(RoundOutput[94]), .B(
        plaintext[94]), .S(reset), .Z(RoundReg_Inst_ff_SDE_94_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_95_current_state_reg_U1 ( .A(ciphertext[95]), 
        .ZN(RoundReg_Inst_ff_SDE_95_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_95_next_state), .CK(clk), .Q(ciphertext[95]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_95_MUX_inst_U1 ( .A(RoundOutput[95]), .B(
        plaintext[95]), .S(reset), .Z(RoundReg_Inst_ff_SDE_95_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_96_current_state_reg_U1 ( .A(ciphertext[0]), 
        .ZN(RoundReg_Inst_ff_SDE_96_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_96_next_state), .CK(clk), .Q(ciphertext[0]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_96_MUX_inst_U1 ( .A(RoundOutput[96]), .B(
        plaintext[96]), .S(reset), .Z(RoundReg_Inst_ff_SDE_96_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_97_current_state_reg_U1 ( .A(ciphertext[1]), 
        .ZN(RoundReg_Inst_ff_SDE_97_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_97_next_state), .CK(clk), .Q(ciphertext[1]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_97_MUX_inst_U1 ( .A(RoundOutput[97]), .B(
        plaintext[97]), .S(reset), .Z(RoundReg_Inst_ff_SDE_97_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_98_current_state_reg_U1 ( .A(ciphertext[2]), 
        .ZN(RoundReg_Inst_ff_SDE_98_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_98_next_state), .CK(clk), .Q(ciphertext[2]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_98_MUX_inst_U1 ( .A(RoundOutput[98]), .B(
        plaintext[98]), .S(reset), .Z(RoundReg_Inst_ff_SDE_98_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_99_current_state_reg_U1 ( .A(ciphertext[3]), 
        .ZN(RoundReg_Inst_ff_SDE_99_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_99_next_state), .CK(clk), .Q(ciphertext[3]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_99_MUX_inst_U1 ( .A(RoundOutput[99]), .B(
        plaintext[99]), .S(reset), .Z(RoundReg_Inst_ff_SDE_99_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_100_current_state_reg_U1 ( .A(ciphertext[4]), 
        .ZN(RoundReg_Inst_ff_SDE_100_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_100_next_state), .CK(clk), .Q(ciphertext[4]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_100_MUX_inst_U1 ( .A(RoundOutput[100]), .B(
        plaintext[100]), .S(reset), .Z(RoundReg_Inst_ff_SDE_100_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_101_current_state_reg_U1 ( .A(ciphertext[5]), 
        .ZN(RoundReg_Inst_ff_SDE_101_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_101_next_state), .CK(clk), .Q(ciphertext[5]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_101_MUX_inst_U1 ( .A(RoundOutput[101]), .B(
        plaintext[101]), .S(reset), .Z(RoundReg_Inst_ff_SDE_101_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_102_current_state_reg_U1 ( .A(ciphertext[6]), 
        .ZN(RoundReg_Inst_ff_SDE_102_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_102_next_state), .CK(clk), .Q(ciphertext[6]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_102_MUX_inst_U1 ( .A(RoundOutput[102]), .B(
        plaintext[102]), .S(reset), .Z(RoundReg_Inst_ff_SDE_102_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_103_current_state_reg_U1 ( .A(ciphertext[7]), 
        .ZN(RoundReg_Inst_ff_SDE_103_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_103_next_state), .CK(clk), .Q(ciphertext[7]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_103_MUX_inst_U1 ( .A(RoundOutput[103]), .B(
        plaintext[103]), .S(reset), .Z(RoundReg_Inst_ff_SDE_103_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_104_current_state_reg_U1 ( .A(ciphertext[40]), 
        .ZN(RoundReg_Inst_ff_SDE_104_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_104_next_state), .CK(clk), .Q(ciphertext[40]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_104_MUX_inst_U1 ( .A(RoundOutput[104]), .B(
        plaintext[104]), .S(reset), .Z(RoundReg_Inst_ff_SDE_104_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_105_current_state_reg_U1 ( .A(ciphertext[41]), 
        .ZN(RoundReg_Inst_ff_SDE_105_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_105_next_state), .CK(clk), .Q(ciphertext[41]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_105_MUX_inst_U1 ( .A(RoundOutput[105]), .B(
        plaintext[105]), .S(reset), .Z(RoundReg_Inst_ff_SDE_105_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_106_current_state_reg_U1 ( .A(ciphertext[42]), 
        .ZN(RoundReg_Inst_ff_SDE_106_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_106_next_state), .CK(clk), .Q(ciphertext[42]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_106_MUX_inst_U1 ( .A(RoundOutput[106]), .B(
        plaintext[106]), .S(reset), .Z(RoundReg_Inst_ff_SDE_106_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_107_current_state_reg_U1 ( .A(ciphertext[43]), 
        .ZN(RoundReg_Inst_ff_SDE_107_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_107_next_state), .CK(clk), .Q(ciphertext[43]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_107_MUX_inst_U1 ( .A(RoundOutput[107]), .B(
        plaintext[107]), .S(reset), .Z(RoundReg_Inst_ff_SDE_107_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_108_current_state_reg_U1 ( .A(ciphertext[44]), 
        .ZN(RoundReg_Inst_ff_SDE_108_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_108_next_state), .CK(clk), .Q(ciphertext[44]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_108_MUX_inst_U1 ( .A(RoundOutput[108]), .B(
        plaintext[108]), .S(reset), .Z(RoundReg_Inst_ff_SDE_108_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_109_current_state_reg_U1 ( .A(ciphertext[45]), 
        .ZN(RoundReg_Inst_ff_SDE_109_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_109_next_state), .CK(clk), .Q(ciphertext[45]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_109_MUX_inst_U1 ( .A(RoundOutput[109]), .B(
        plaintext[109]), .S(reset), .Z(RoundReg_Inst_ff_SDE_109_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_110_current_state_reg_U1 ( .A(ciphertext[46]), 
        .ZN(RoundReg_Inst_ff_SDE_110_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_110_next_state), .CK(clk), .Q(ciphertext[46]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_110_MUX_inst_U1 ( .A(RoundOutput[110]), .B(
        plaintext[110]), .S(reset), .Z(RoundReg_Inst_ff_SDE_110_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_111_current_state_reg_U1 ( .A(ciphertext[47]), 
        .ZN(RoundReg_Inst_ff_SDE_111_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_111_next_state), .CK(clk), .Q(ciphertext[47]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_111_MUX_inst_U1 ( .A(RoundOutput[111]), .B(
        plaintext[111]), .S(reset), .Z(RoundReg_Inst_ff_SDE_111_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_112_current_state_reg_U1 ( .A(ciphertext[80]), 
        .ZN(RoundReg_Inst_ff_SDE_112_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_112_next_state), .CK(clk), .Q(ciphertext[80]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_112_MUX_inst_U1 ( .A(RoundOutput[112]), .B(
        plaintext[112]), .S(reset), .Z(RoundReg_Inst_ff_SDE_112_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_113_current_state_reg_U1 ( .A(ciphertext[81]), 
        .ZN(RoundReg_Inst_ff_SDE_113_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_113_next_state), .CK(clk), .Q(ciphertext[81]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_113_MUX_inst_U1 ( .A(RoundOutput[113]), .B(
        plaintext[113]), .S(reset), .Z(RoundReg_Inst_ff_SDE_113_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_114_current_state_reg_U1 ( .A(ciphertext[82]), 
        .ZN(RoundReg_Inst_ff_SDE_114_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_114_next_state), .CK(clk), .Q(ciphertext[82]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_114_MUX_inst_U1 ( .A(RoundOutput[114]), .B(
        plaintext[114]), .S(reset), .Z(RoundReg_Inst_ff_SDE_114_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_115_current_state_reg_U1 ( .A(ciphertext[83]), 
        .ZN(RoundReg_Inst_ff_SDE_115_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_115_next_state), .CK(clk), .Q(ciphertext[83]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_115_MUX_inst_U1 ( .A(RoundOutput[115]), .B(
        plaintext[115]), .S(reset), .Z(RoundReg_Inst_ff_SDE_115_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_116_current_state_reg_U1 ( .A(ciphertext[84]), 
        .ZN(RoundReg_Inst_ff_SDE_116_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_116_next_state), .CK(clk), .Q(ciphertext[84]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_116_MUX_inst_U1 ( .A(RoundOutput[116]), .B(
        plaintext[116]), .S(reset), .Z(RoundReg_Inst_ff_SDE_116_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_117_current_state_reg_U1 ( .A(ciphertext[85]), 
        .ZN(RoundReg_Inst_ff_SDE_117_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_117_next_state), .CK(clk), .Q(ciphertext[85]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_117_MUX_inst_U1 ( .A(RoundOutput[117]), .B(
        plaintext[117]), .S(reset), .Z(RoundReg_Inst_ff_SDE_117_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_118_current_state_reg_U1 ( .A(ciphertext[86]), 
        .ZN(RoundReg_Inst_ff_SDE_118_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_118_next_state), .CK(clk), .Q(ciphertext[86]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_118_MUX_inst_U1 ( .A(RoundOutput[118]), .B(
        plaintext[118]), .S(reset), .Z(RoundReg_Inst_ff_SDE_118_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_119_current_state_reg_U1 ( .A(ciphertext[87]), 
        .ZN(RoundReg_Inst_ff_SDE_119_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_119_next_state), .CK(clk), .Q(ciphertext[87]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_119_MUX_inst_U1 ( .A(RoundOutput[119]), .B(
        plaintext[119]), .S(reset), .Z(RoundReg_Inst_ff_SDE_119_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_120_current_state_reg_U1 ( .A(ciphertext[120]), 
        .ZN(RoundReg_Inst_ff_SDE_120_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_120_next_state), .CK(clk), .Q(ciphertext[120]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_120_MUX_inst_U1 ( .A(RoundOutput[120]), .B(
        plaintext[120]), .S(reset), .Z(RoundReg_Inst_ff_SDE_120_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_121_current_state_reg_U1 ( .A(ciphertext[121]), 
        .ZN(RoundReg_Inst_ff_SDE_121_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_121_next_state), .CK(clk), .Q(ciphertext[121]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_121_MUX_inst_U1 ( .A(RoundOutput[121]), .B(
        plaintext[121]), .S(reset), .Z(RoundReg_Inst_ff_SDE_121_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_122_current_state_reg_U1 ( .A(ciphertext[122]), 
        .ZN(RoundReg_Inst_ff_SDE_122_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_122_next_state), .CK(clk), .Q(ciphertext[122]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_122_MUX_inst_U1 ( .A(RoundOutput[122]), .B(
        plaintext[122]), .S(reset), .Z(RoundReg_Inst_ff_SDE_122_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_123_current_state_reg_U1 ( .A(ciphertext[123]), 
        .ZN(RoundReg_Inst_ff_SDE_123_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_123_next_state), .CK(clk), .Q(ciphertext[123]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_123_MUX_inst_U1 ( .A(RoundOutput[123]), .B(
        plaintext[123]), .S(reset), .Z(RoundReg_Inst_ff_SDE_123_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_124_current_state_reg_U1 ( .A(ciphertext[124]), 
        .ZN(RoundReg_Inst_ff_SDE_124_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_124_next_state), .CK(clk), .Q(ciphertext[124]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_124_MUX_inst_U1 ( .A(RoundOutput[124]), .B(
        plaintext[124]), .S(reset), .Z(RoundReg_Inst_ff_SDE_124_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_125_current_state_reg_U1 ( .A(ciphertext[125]), 
        .ZN(RoundReg_Inst_ff_SDE_125_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_125_next_state), .CK(clk), .Q(ciphertext[125]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_125_MUX_inst_U1 ( .A(RoundOutput[125]), .B(
        plaintext[125]), .S(reset), .Z(RoundReg_Inst_ff_SDE_125_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_126_current_state_reg_U1 ( .A(ciphertext[126]), 
        .ZN(RoundReg_Inst_ff_SDE_126_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_126_next_state), .CK(clk), .Q(ciphertext[126]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_126_MUX_inst_U1 ( .A(RoundOutput[126]), .B(
        plaintext[126]), .S(reset), .Z(RoundReg_Inst_ff_SDE_126_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_127_current_state_reg_U1 ( .A(ciphertext[127]), 
        .ZN(RoundReg_Inst_ff_SDE_127_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_127_next_state), .CK(clk), .Q(ciphertext[127]), 
        .QN() );
  MUX2_X1 RoundReg_Inst_ff_SDE_127_MUX_inst_U1 ( .A(RoundOutput[127]), .B(
        plaintext[127]), .S(reset), .Z(RoundReg_Inst_ff_SDE_127_next_state) );
  INV_X1 MuxSboxIn_U3 ( .A(AKSRnotDone), .ZN(MuxSboxIn_n7) );
  INV_X1 MuxSboxIn_U2 ( .A(MuxSboxIn_n7), .ZN(MuxSboxIn_n5) );
  INV_X1 MuxSboxIn_U1 ( .A(MuxSboxIn_n7), .ZN(MuxSboxIn_n6) );
  MUX2_X1 MuxSboxIn_mux_inst_0_U1 ( .A(ciphertext[0]), .B(KSSubBytesInput[0]), 
        .S(MuxSboxIn_n6), .Z(SubBytesInput[0]) );
  MUX2_X1 MuxSboxIn_mux_inst_1_U1 ( .A(ciphertext[1]), .B(KSSubBytesInput[1]), 
        .S(MuxSboxIn_n6), .Z(SubBytesInput[1]) );
  MUX2_X1 MuxSboxIn_mux_inst_2_U1 ( .A(ciphertext[2]), .B(KSSubBytesInput[2]), 
        .S(MuxSboxIn_n6), .Z(SubBytesInput[2]) );
  MUX2_X1 MuxSboxIn_mux_inst_3_U1 ( .A(ciphertext[3]), .B(KSSubBytesInput[3]), 
        .S(MuxSboxIn_n6), .Z(SubBytesInput[3]) );
  MUX2_X1 MuxSboxIn_mux_inst_4_U1 ( .A(ciphertext[4]), .B(KSSubBytesInput[4]), 
        .S(MuxSboxIn_n6), .Z(SubBytesInput[4]) );
  MUX2_X1 MuxSboxIn_mux_inst_5_U1 ( .A(ciphertext[5]), .B(KSSubBytesInput[5]), 
        .S(MuxSboxIn_n6), .Z(SubBytesInput[5]) );
  MUX2_X1 MuxSboxIn_mux_inst_6_U1 ( .A(ciphertext[6]), .B(KSSubBytesInput[6]), 
        .S(MuxSboxIn_n6), .Z(SubBytesInput[6]) );
  MUX2_X1 MuxSboxIn_mux_inst_7_U1 ( .A(ciphertext[7]), .B(KSSubBytesInput[7]), 
        .S(MuxSboxIn_n6), .Z(SubBytesInput[7]) );
  MUX2_X1 MuxSboxIn_mux_inst_8_U1 ( .A(ciphertext[40]), .B(KSSubBytesInput[8]), 
        .S(AKSRnotDone), .Z(SubBytesInput[8]) );
  MUX2_X1 MuxSboxIn_mux_inst_9_U1 ( .A(ciphertext[41]), .B(KSSubBytesInput[9]), 
        .S(MuxSboxIn_n5), .Z(SubBytesInput[9]) );
  MUX2_X1 MuxSboxIn_mux_inst_10_U1 ( .A(ciphertext[42]), .B(
        KSSubBytesInput[10]), .S(MuxSboxIn_n5), .Z(SubBytesInput[10]) );
  MUX2_X1 MuxSboxIn_mux_inst_11_U1 ( .A(ciphertext[43]), .B(
        KSSubBytesInput[11]), .S(MuxSboxIn_n5), .Z(SubBytesInput[11]) );
  MUX2_X1 MuxSboxIn_mux_inst_12_U1 ( .A(ciphertext[44]), .B(
        KSSubBytesInput[12]), .S(MuxSboxIn_n5), .Z(SubBytesInput[12]) );
  MUX2_X1 MuxSboxIn_mux_inst_13_U1 ( .A(ciphertext[45]), .B(
        KSSubBytesInput[13]), .S(MuxSboxIn_n6), .Z(SubBytesInput[13]) );
  MUX2_X1 MuxSboxIn_mux_inst_14_U1 ( .A(ciphertext[46]), .B(
        KSSubBytesInput[14]), .S(MuxSboxIn_n6), .Z(SubBytesInput[14]) );
  MUX2_X1 MuxSboxIn_mux_inst_15_U1 ( .A(ciphertext[47]), .B(
        KSSubBytesInput[15]), .S(MuxSboxIn_n5), .Z(SubBytesInput[15]) );
  MUX2_X1 MuxSboxIn_mux_inst_16_U1 ( .A(ciphertext[80]), .B(
        KSSubBytesInput[16]), .S(MuxSboxIn_n6), .Z(SubBytesInput[16]) );
  MUX2_X1 MuxSboxIn_mux_inst_17_U1 ( .A(ciphertext[81]), .B(
        KSSubBytesInput[17]), .S(MuxSboxIn_n5), .Z(SubBytesInput[17]) );
  MUX2_X1 MuxSboxIn_mux_inst_18_U1 ( .A(ciphertext[82]), .B(
        KSSubBytesInput[18]), .S(MuxSboxIn_n5), .Z(SubBytesInput[18]) );
  MUX2_X1 MuxSboxIn_mux_inst_19_U1 ( .A(ciphertext[83]), .B(
        KSSubBytesInput[19]), .S(MuxSboxIn_n5), .Z(SubBytesInput[19]) );
  MUX2_X1 MuxSboxIn_mux_inst_20_U1 ( .A(ciphertext[84]), .B(
        KSSubBytesInput[20]), .S(MuxSboxIn_n5), .Z(SubBytesInput[20]) );
  MUX2_X1 MuxSboxIn_mux_inst_21_U1 ( .A(ciphertext[85]), .B(
        KSSubBytesInput[21]), .S(MuxSboxIn_n5), .Z(SubBytesInput[21]) );
  MUX2_X1 MuxSboxIn_mux_inst_22_U1 ( .A(ciphertext[86]), .B(
        KSSubBytesInput[22]), .S(MuxSboxIn_n5), .Z(SubBytesInput[22]) );
  MUX2_X1 MuxSboxIn_mux_inst_23_U1 ( .A(ciphertext[87]), .B(
        KSSubBytesInput[23]), .S(MuxSboxIn_n5), .Z(SubBytesInput[23]) );
  MUX2_X1 MuxSboxIn_mux_inst_24_U1 ( .A(ciphertext[120]), .B(
        KSSubBytesInput[24]), .S(MuxSboxIn_n5), .Z(SubBytesInput[24]) );
  MUX2_X1 MuxSboxIn_mux_inst_25_U1 ( .A(ciphertext[121]), .B(
        KSSubBytesInput[25]), .S(MuxSboxIn_n5), .Z(SubBytesInput[25]) );
  MUX2_X1 MuxSboxIn_mux_inst_26_U1 ( .A(ciphertext[122]), .B(
        KSSubBytesInput[26]), .S(MuxSboxIn_n5), .Z(SubBytesInput[26]) );
  MUX2_X1 MuxSboxIn_mux_inst_27_U1 ( .A(ciphertext[123]), .B(
        KSSubBytesInput[27]), .S(MuxSboxIn_n5), .Z(SubBytesInput[27]) );
  MUX2_X1 MuxSboxIn_mux_inst_28_U1 ( .A(ciphertext[124]), .B(
        KSSubBytesInput[28]), .S(MuxSboxIn_n5), .Z(SubBytesInput[28]) );
  MUX2_X1 MuxSboxIn_mux_inst_29_U1 ( .A(ciphertext[125]), .B(
        KSSubBytesInput[29]), .S(MuxSboxIn_n5), .Z(SubBytesInput[29]) );
  MUX2_X1 MuxSboxIn_mux_inst_30_U1 ( .A(ciphertext[126]), .B(
        KSSubBytesInput[30]), .S(MuxSboxIn_n5), .Z(SubBytesInput[30]) );
  MUX2_X1 MuxSboxIn_mux_inst_31_U1 ( .A(ciphertext[127]), .B(
        KSSubBytesInput[31]), .S(MuxSboxIn_n5), .Z(SubBytesInput[31]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T1_U1 ( .A(SubBytesInput[7]), .B(
        SubBytesInput[4]), .Z(SubBytesIns_Inst_Sbox_0_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T2_U1 ( .A(SubBytesInput[7]), .B(
        SubBytesInput[2]), .Z(SubBytesIns_Inst_Sbox_0_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T3_U1 ( .A(SubBytesInput[7]), .B(
        SubBytesInput[1]), .Z(SubBytesIns_Inst_Sbox_0_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T4_U1 ( .A(SubBytesInput[4]), .B(
        SubBytesInput[2]), .Z(SubBytesIns_Inst_Sbox_0_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T5_U1 ( .A(SubBytesInput[3]), .B(
        SubBytesInput[1]), .Z(SubBytesIns_Inst_Sbox_0_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_0_T1), 
        .B(SubBytesIns_Inst_Sbox_0_T5), .Z(SubBytesIns_Inst_Sbox_0_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T7_U1 ( .A(SubBytesInput[6]), .B(
        SubBytesInput[5]), .Z(SubBytesIns_Inst_Sbox_0_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T8_U1 ( .A(SubBytesInput[0]), .B(
        SubBytesIns_Inst_Sbox_0_T6), .Z(SubBytesIns_Inst_Sbox_0_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T9_U1 ( .A(SubBytesInput[0]), .B(
        SubBytesIns_Inst_Sbox_0_T7), .Z(SubBytesIns_Inst_Sbox_0_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_0_T6), 
        .B(SubBytesIns_Inst_Sbox_0_T7), .Z(SubBytesIns_Inst_Sbox_0_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T11_U1 ( .A(SubBytesInput[6]), .B(
        SubBytesInput[2]), .Z(SubBytesIns_Inst_Sbox_0_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T12_U1 ( .A(SubBytesInput[5]), .B(
        SubBytesInput[2]), .Z(SubBytesIns_Inst_Sbox_0_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_0_T3), 
        .B(SubBytesIns_Inst_Sbox_0_T4), .Z(SubBytesIns_Inst_Sbox_0_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_0_T6), 
        .B(SubBytesIns_Inst_Sbox_0_T11), .Z(SubBytesIns_Inst_Sbox_0_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_0_T5), 
        .B(SubBytesIns_Inst_Sbox_0_T11), .Z(SubBytesIns_Inst_Sbox_0_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_0_T5), 
        .B(SubBytesIns_Inst_Sbox_0_T12), .Z(SubBytesIns_Inst_Sbox_0_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_0_T9), 
        .B(SubBytesIns_Inst_Sbox_0_T16), .Z(SubBytesIns_Inst_Sbox_0_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T18_U1 ( .A(SubBytesInput[4]), .B(
        SubBytesInput[0]), .Z(SubBytesIns_Inst_Sbox_0_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_0_T7), 
        .B(SubBytesIns_Inst_Sbox_0_T18), .Z(SubBytesIns_Inst_Sbox_0_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_0_T1), 
        .B(SubBytesIns_Inst_Sbox_0_T19), .Z(SubBytesIns_Inst_Sbox_0_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T21_U1 ( .A(SubBytesInput[1]), .B(
        SubBytesInput[0]), .Z(SubBytesIns_Inst_Sbox_0_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_0_T7), 
        .B(SubBytesIns_Inst_Sbox_0_T21), .Z(SubBytesIns_Inst_Sbox_0_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_0_T2), 
        .B(SubBytesIns_Inst_Sbox_0_T22), .Z(SubBytesIns_Inst_Sbox_0_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_0_T2), 
        .B(SubBytesIns_Inst_Sbox_0_T10), .Z(SubBytesIns_Inst_Sbox_0_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_0_T20), 
        .B(SubBytesIns_Inst_Sbox_0_T17), .Z(SubBytesIns_Inst_Sbox_0_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_0_T3), 
        .B(SubBytesIns_Inst_Sbox_0_T16), .Z(SubBytesIns_Inst_Sbox_0_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_0_T1), 
        .B(SubBytesIns_Inst_Sbox_0_T12), .Z(SubBytesIns_Inst_Sbox_0_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T13), 
        .A2(SubBytesIns_Inst_Sbox_0_T6), .ZN(SubBytesIns_Inst_Sbox_0_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T23), 
        .A2(SubBytesIns_Inst_Sbox_0_T8), .ZN(SubBytesIns_Inst_Sbox_0_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_0_T14), 
        .B(SubBytesIns_Inst_Sbox_0_M1), .Z(SubBytesIns_Inst_Sbox_0_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T19), 
        .A2(SubBytesInput[0]), .ZN(SubBytesIns_Inst_Sbox_0_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_0_M4), 
        .B(SubBytesIns_Inst_Sbox_0_M1), .Z(SubBytesIns_Inst_Sbox_0_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T3), 
        .A2(SubBytesIns_Inst_Sbox_0_T16), .ZN(SubBytesIns_Inst_Sbox_0_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T22), 
        .A2(SubBytesIns_Inst_Sbox_0_T9), .ZN(SubBytesIns_Inst_Sbox_0_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_0_T26), 
        .B(SubBytesIns_Inst_Sbox_0_M6), .Z(SubBytesIns_Inst_Sbox_0_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T20), 
        .A2(SubBytesIns_Inst_Sbox_0_T17), .ZN(SubBytesIns_Inst_Sbox_0_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_0_M9), 
        .B(SubBytesIns_Inst_Sbox_0_M6), .Z(SubBytesIns_Inst_Sbox_0_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T1), 
        .A2(SubBytesIns_Inst_Sbox_0_T15), .ZN(SubBytesIns_Inst_Sbox_0_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T4), 
        .A2(SubBytesIns_Inst_Sbox_0_T27), .ZN(SubBytesIns_Inst_Sbox_0_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_0_M12), 
        .B(SubBytesIns_Inst_Sbox_0_M11), .Z(SubBytesIns_Inst_Sbox_0_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T2), 
        .A2(SubBytesIns_Inst_Sbox_0_T10), .ZN(SubBytesIns_Inst_Sbox_0_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_0_M14), 
        .B(SubBytesIns_Inst_Sbox_0_M11), .Z(SubBytesIns_Inst_Sbox_0_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_0_M3), 
        .B(SubBytesIns_Inst_Sbox_0_M2), .Z(SubBytesIns_Inst_Sbox_0_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_0_M5), 
        .B(SubBytesIns_Inst_Sbox_0_T24), .Z(SubBytesIns_Inst_Sbox_0_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_0_M8), 
        .B(SubBytesIns_Inst_Sbox_0_M7), .Z(SubBytesIns_Inst_Sbox_0_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_0_M10), 
        .B(SubBytesIns_Inst_Sbox_0_M15), .Z(SubBytesIns_Inst_Sbox_0_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_0_M16), 
        .B(SubBytesIns_Inst_Sbox_0_M13), .Z(SubBytesIns_Inst_Sbox_0_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_0_M17), 
        .B(SubBytesIns_Inst_Sbox_0_M15), .Z(SubBytesIns_Inst_Sbox_0_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_0_M18), 
        .B(SubBytesIns_Inst_Sbox_0_M13), .Z(SubBytesIns_Inst_Sbox_0_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_0_M19), 
        .B(SubBytesIns_Inst_Sbox_0_T25), .Z(SubBytesIns_Inst_Sbox_0_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_0_M22), 
        .B(SubBytesIns_Inst_Sbox_0_M23), .Z(SubBytesIns_Inst_Sbox_0_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M22), .A2(SubBytesIns_Inst_Sbox_0_M20), .ZN(SubBytesIns_Inst_Sbox_0_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_0_M21), 
        .B(SubBytesIns_Inst_Sbox_0_M25), .Z(SubBytesIns_Inst_Sbox_0_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_0_M20), 
        .B(SubBytesIns_Inst_Sbox_0_M21), .Z(SubBytesIns_Inst_Sbox_0_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_0_M23), 
        .B(SubBytesIns_Inst_Sbox_0_M25), .Z(SubBytesIns_Inst_Sbox_0_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M28), .A2(SubBytesIns_Inst_Sbox_0_M27), .ZN(SubBytesIns_Inst_Sbox_0_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M26), .A2(SubBytesIns_Inst_Sbox_0_M24), .ZN(SubBytesIns_Inst_Sbox_0_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M20), .A2(SubBytesIns_Inst_Sbox_0_M23), .ZN(SubBytesIns_Inst_Sbox_0_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M27), .A2(SubBytesIns_Inst_Sbox_0_M31), .ZN(SubBytesIns_Inst_Sbox_0_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_0_M27), 
        .B(SubBytesIns_Inst_Sbox_0_M25), .Z(SubBytesIns_Inst_Sbox_0_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M21), .A2(SubBytesIns_Inst_Sbox_0_M22), .ZN(SubBytesIns_Inst_Sbox_0_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M24), .A2(SubBytesIns_Inst_Sbox_0_M34), .ZN(SubBytesIns_Inst_Sbox_0_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_0_M24), 
        .B(SubBytesIns_Inst_Sbox_0_M25), .Z(SubBytesIns_Inst_Sbox_0_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_0_M21), 
        .B(SubBytesIns_Inst_Sbox_0_M29), .Z(SubBytesIns_Inst_Sbox_0_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_0_M32), 
        .B(SubBytesIns_Inst_Sbox_0_M33), .Z(SubBytesIns_Inst_Sbox_0_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_0_M23), 
        .B(SubBytesIns_Inst_Sbox_0_M30), .Z(SubBytesIns_Inst_Sbox_0_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_0_M35), 
        .B(SubBytesIns_Inst_Sbox_0_M36), .Z(SubBytesIns_Inst_Sbox_0_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_0_M38), 
        .B(SubBytesIns_Inst_Sbox_0_M40), .Z(SubBytesIns_Inst_Sbox_0_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_0_M37), 
        .B(SubBytesIns_Inst_Sbox_0_M39), .Z(SubBytesIns_Inst_Sbox_0_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_0_M37), 
        .B(SubBytesIns_Inst_Sbox_0_M38), .Z(SubBytesIns_Inst_Sbox_0_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_0_M39), 
        .B(SubBytesIns_Inst_Sbox_0_M40), .Z(SubBytesIns_Inst_Sbox_0_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_0_M42), 
        .B(SubBytesIns_Inst_Sbox_0_M41), .Z(SubBytesIns_Inst_Sbox_0_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M44), .A2(SubBytesIns_Inst_Sbox_0_T6), .ZN(SubBytesIns_Inst_Sbox_0_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M40), .A2(SubBytesIns_Inst_Sbox_0_T8), .ZN(SubBytesIns_Inst_Sbox_0_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M39), .A2(SubBytesInput[0]), .ZN(SubBytesIns_Inst_Sbox_0_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M43), .A2(SubBytesIns_Inst_Sbox_0_T16), .ZN(SubBytesIns_Inst_Sbox_0_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M38), .A2(SubBytesIns_Inst_Sbox_0_T9), .ZN(SubBytesIns_Inst_Sbox_0_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M37), .A2(SubBytesIns_Inst_Sbox_0_T17), .ZN(SubBytesIns_Inst_Sbox_0_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M42), .A2(SubBytesIns_Inst_Sbox_0_T15), .ZN(SubBytesIns_Inst_Sbox_0_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M45), .A2(SubBytesIns_Inst_Sbox_0_T27), .ZN(SubBytesIns_Inst_Sbox_0_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M41), .A2(SubBytesIns_Inst_Sbox_0_T10), .ZN(SubBytesIns_Inst_Sbox_0_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M44), .A2(SubBytesIns_Inst_Sbox_0_T13), .ZN(SubBytesIns_Inst_Sbox_0_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M40), .A2(SubBytesIns_Inst_Sbox_0_T23), .ZN(SubBytesIns_Inst_Sbox_0_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M39), .A2(SubBytesIns_Inst_Sbox_0_T19), .ZN(SubBytesIns_Inst_Sbox_0_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M43), .A2(SubBytesIns_Inst_Sbox_0_T3), .ZN(SubBytesIns_Inst_Sbox_0_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M38), .A2(SubBytesIns_Inst_Sbox_0_T22), .ZN(SubBytesIns_Inst_Sbox_0_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M37), .A2(SubBytesIns_Inst_Sbox_0_T20), .ZN(SubBytesIns_Inst_Sbox_0_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M42), .A2(SubBytesIns_Inst_Sbox_0_T1), .ZN(SubBytesIns_Inst_Sbox_0_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M45), .A2(SubBytesIns_Inst_Sbox_0_T4), .ZN(SubBytesIns_Inst_Sbox_0_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M41), .A2(SubBytesIns_Inst_Sbox_0_T2), .ZN(SubBytesIns_Inst_Sbox_0_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_0_M61), 
        .B(SubBytesIns_Inst_Sbox_0_M62), .Z(SubBytesIns_Inst_Sbox_0_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_0_M50), 
        .B(SubBytesIns_Inst_Sbox_0_M56), .Z(SubBytesIns_Inst_Sbox_0_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_0_M46), 
        .B(SubBytesIns_Inst_Sbox_0_M48), .Z(SubBytesIns_Inst_Sbox_0_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_0_M47), 
        .B(SubBytesIns_Inst_Sbox_0_M55), .Z(SubBytesIns_Inst_Sbox_0_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_0_M54), 
        .B(SubBytesIns_Inst_Sbox_0_M58), .Z(SubBytesIns_Inst_Sbox_0_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_0_M49), 
        .B(SubBytesIns_Inst_Sbox_0_M61), .Z(SubBytesIns_Inst_Sbox_0_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_0_M62), 
        .B(SubBytesIns_Inst_Sbox_0_L5), .Z(SubBytesIns_Inst_Sbox_0_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_0_M46), 
        .B(SubBytesIns_Inst_Sbox_0_L3), .Z(SubBytesIns_Inst_Sbox_0_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_0_M51), 
        .B(SubBytesIns_Inst_Sbox_0_M59), .Z(SubBytesIns_Inst_Sbox_0_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_0_M52), 
        .B(SubBytesIns_Inst_Sbox_0_M53), .Z(SubBytesIns_Inst_Sbox_0_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_0_M53), 
        .B(SubBytesIns_Inst_Sbox_0_L4), .Z(SubBytesIns_Inst_Sbox_0_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_0_M60), 
        .B(SubBytesIns_Inst_Sbox_0_L2), .Z(SubBytesIns_Inst_Sbox_0_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_0_M48), 
        .B(SubBytesIns_Inst_Sbox_0_M51), .Z(SubBytesIns_Inst_Sbox_0_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_0_M50), 
        .B(SubBytesIns_Inst_Sbox_0_L0), .Z(SubBytesIns_Inst_Sbox_0_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_0_M52), 
        .B(SubBytesIns_Inst_Sbox_0_M61), .Z(SubBytesIns_Inst_Sbox_0_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_0_M55), 
        .B(SubBytesIns_Inst_Sbox_0_L1), .Z(SubBytesIns_Inst_Sbox_0_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_0_M56), 
        .B(SubBytesIns_Inst_Sbox_0_L0), .Z(SubBytesIns_Inst_Sbox_0_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_0_M57), 
        .B(SubBytesIns_Inst_Sbox_0_L1), .Z(SubBytesIns_Inst_Sbox_0_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_0_M58), 
        .B(SubBytesIns_Inst_Sbox_0_L8), .Z(SubBytesIns_Inst_Sbox_0_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_0_M63), 
        .B(SubBytesIns_Inst_Sbox_0_L4), .Z(SubBytesIns_Inst_Sbox_0_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_0_L0), 
        .B(SubBytesIns_Inst_Sbox_0_L1), .Z(SubBytesIns_Inst_Sbox_0_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_0_L1), 
        .B(SubBytesIns_Inst_Sbox_0_L7), .Z(SubBytesIns_Inst_Sbox_0_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_0_L3), 
        .B(SubBytesIns_Inst_Sbox_0_L12), .Z(SubBytesIns_Inst_Sbox_0_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_0_L18), 
        .B(SubBytesIns_Inst_Sbox_0_L2), .Z(SubBytesIns_Inst_Sbox_0_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_0_L15), 
        .B(SubBytesIns_Inst_Sbox_0_L9), .Z(SubBytesIns_Inst_Sbox_0_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_0_L6), 
        .B(SubBytesIns_Inst_Sbox_0_L10), .Z(SubBytesIns_Inst_Sbox_0_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_0_L7), 
        .B(SubBytesIns_Inst_Sbox_0_L9), .Z(SubBytesIns_Inst_Sbox_0_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_0_L8), 
        .B(SubBytesIns_Inst_Sbox_0_L10), .Z(SubBytesIns_Inst_Sbox_0_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_0_L11), 
        .B(SubBytesIns_Inst_Sbox_0_L14), .Z(SubBytesIns_Inst_Sbox_0_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_0_L11), 
        .B(SubBytesIns_Inst_Sbox_0_L17), .Z(SubBytesIns_Inst_Sbox_0_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_0_L6), 
        .B(SubBytesIns_Inst_Sbox_0_L24), .Z(MixColumnsIns_DoubleBytes[0]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_0_L16), 
        .B(SubBytesIns_Inst_Sbox_0_L26), .ZN(MixColumnsIns_DoubleBytes[7]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_0_L19), 
        .B(SubBytesIns_Inst_Sbox_0_L28), .ZN(MixColumnsIns_DoubleBytes[6]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_0_L6), 
        .B(SubBytesIns_Inst_Sbox_0_L21), .Z(MixColumnsIns_DoubleBytes[5]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_0_L20), 
        .B(SubBytesIns_Inst_Sbox_0_L22), .Z(SubBytesOutput[3]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_0_L25), 
        .B(SubBytesIns_Inst_Sbox_0_L29), .Z(SubBytesOutput[2]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_0_L13), 
        .B(SubBytesIns_Inst_Sbox_0_L27), .ZN(MixColumnsIns_DoubleBytes[2]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_0_L6), 
        .B(SubBytesIns_Inst_Sbox_0_L23), .ZN(SubBytesOutput[0]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T1_U1 ( .A(SubBytesInput[15]), .B(
        SubBytesInput[12]), .Z(SubBytesIns_Inst_Sbox_1_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T2_U1 ( .A(SubBytesInput[15]), .B(
        SubBytesInput[10]), .Z(SubBytesIns_Inst_Sbox_1_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T3_U1 ( .A(SubBytesInput[15]), .B(
        SubBytesInput[9]), .Z(SubBytesIns_Inst_Sbox_1_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T4_U1 ( .A(SubBytesInput[12]), .B(
        SubBytesInput[10]), .Z(SubBytesIns_Inst_Sbox_1_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T5_U1 ( .A(SubBytesInput[11]), .B(
        SubBytesInput[9]), .Z(SubBytesIns_Inst_Sbox_1_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_1_T1), 
        .B(SubBytesIns_Inst_Sbox_1_T5), .Z(SubBytesIns_Inst_Sbox_1_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T7_U1 ( .A(SubBytesInput[14]), .B(
        SubBytesInput[13]), .Z(SubBytesIns_Inst_Sbox_1_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T8_U1 ( .A(SubBytesInput[8]), .B(
        SubBytesIns_Inst_Sbox_1_T6), .Z(SubBytesIns_Inst_Sbox_1_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T9_U1 ( .A(SubBytesInput[8]), .B(
        SubBytesIns_Inst_Sbox_1_T7), .Z(SubBytesIns_Inst_Sbox_1_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_1_T6), 
        .B(SubBytesIns_Inst_Sbox_1_T7), .Z(SubBytesIns_Inst_Sbox_1_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T11_U1 ( .A(SubBytesInput[14]), .B(
        SubBytesInput[10]), .Z(SubBytesIns_Inst_Sbox_1_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T12_U1 ( .A(SubBytesInput[13]), .B(
        SubBytesInput[10]), .Z(SubBytesIns_Inst_Sbox_1_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_1_T3), 
        .B(SubBytesIns_Inst_Sbox_1_T4), .Z(SubBytesIns_Inst_Sbox_1_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_1_T6), 
        .B(SubBytesIns_Inst_Sbox_1_T11), .Z(SubBytesIns_Inst_Sbox_1_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_1_T5), 
        .B(SubBytesIns_Inst_Sbox_1_T11), .Z(SubBytesIns_Inst_Sbox_1_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_1_T5), 
        .B(SubBytesIns_Inst_Sbox_1_T12), .Z(SubBytesIns_Inst_Sbox_1_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_1_T9), 
        .B(SubBytesIns_Inst_Sbox_1_T16), .Z(SubBytesIns_Inst_Sbox_1_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T18_U1 ( .A(SubBytesInput[12]), .B(
        SubBytesInput[8]), .Z(SubBytesIns_Inst_Sbox_1_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_1_T7), 
        .B(SubBytesIns_Inst_Sbox_1_T18), .Z(SubBytesIns_Inst_Sbox_1_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_1_T1), 
        .B(SubBytesIns_Inst_Sbox_1_T19), .Z(SubBytesIns_Inst_Sbox_1_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T21_U1 ( .A(SubBytesInput[9]), .B(
        SubBytesInput[8]), .Z(SubBytesIns_Inst_Sbox_1_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_1_T7), 
        .B(SubBytesIns_Inst_Sbox_1_T21), .Z(SubBytesIns_Inst_Sbox_1_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_1_T2), 
        .B(SubBytesIns_Inst_Sbox_1_T22), .Z(SubBytesIns_Inst_Sbox_1_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_1_T2), 
        .B(SubBytesIns_Inst_Sbox_1_T10), .Z(SubBytesIns_Inst_Sbox_1_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_1_T20), 
        .B(SubBytesIns_Inst_Sbox_1_T17), .Z(SubBytesIns_Inst_Sbox_1_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_1_T3), 
        .B(SubBytesIns_Inst_Sbox_1_T16), .Z(SubBytesIns_Inst_Sbox_1_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_1_T1), 
        .B(SubBytesIns_Inst_Sbox_1_T12), .Z(SubBytesIns_Inst_Sbox_1_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T13), 
        .A2(SubBytesIns_Inst_Sbox_1_T6), .ZN(SubBytesIns_Inst_Sbox_1_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T23), 
        .A2(SubBytesIns_Inst_Sbox_1_T8), .ZN(SubBytesIns_Inst_Sbox_1_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_1_T14), 
        .B(SubBytesIns_Inst_Sbox_1_M1), .Z(SubBytesIns_Inst_Sbox_1_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T19), 
        .A2(SubBytesInput[8]), .ZN(SubBytesIns_Inst_Sbox_1_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_1_M4), 
        .B(SubBytesIns_Inst_Sbox_1_M1), .Z(SubBytesIns_Inst_Sbox_1_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T3), 
        .A2(SubBytesIns_Inst_Sbox_1_T16), .ZN(SubBytesIns_Inst_Sbox_1_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T22), 
        .A2(SubBytesIns_Inst_Sbox_1_T9), .ZN(SubBytesIns_Inst_Sbox_1_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_1_T26), 
        .B(SubBytesIns_Inst_Sbox_1_M6), .Z(SubBytesIns_Inst_Sbox_1_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T20), 
        .A2(SubBytesIns_Inst_Sbox_1_T17), .ZN(SubBytesIns_Inst_Sbox_1_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_1_M9), 
        .B(SubBytesIns_Inst_Sbox_1_M6), .Z(SubBytesIns_Inst_Sbox_1_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T1), 
        .A2(SubBytesIns_Inst_Sbox_1_T15), .ZN(SubBytesIns_Inst_Sbox_1_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T4), 
        .A2(SubBytesIns_Inst_Sbox_1_T27), .ZN(SubBytesIns_Inst_Sbox_1_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_1_M12), 
        .B(SubBytesIns_Inst_Sbox_1_M11), .Z(SubBytesIns_Inst_Sbox_1_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T2), 
        .A2(SubBytesIns_Inst_Sbox_1_T10), .ZN(SubBytesIns_Inst_Sbox_1_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_1_M14), 
        .B(SubBytesIns_Inst_Sbox_1_M11), .Z(SubBytesIns_Inst_Sbox_1_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_1_M3), 
        .B(SubBytesIns_Inst_Sbox_1_M2), .Z(SubBytesIns_Inst_Sbox_1_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_1_M5), 
        .B(SubBytesIns_Inst_Sbox_1_T24), .Z(SubBytesIns_Inst_Sbox_1_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_1_M8), 
        .B(SubBytesIns_Inst_Sbox_1_M7), .Z(SubBytesIns_Inst_Sbox_1_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_1_M10), 
        .B(SubBytesIns_Inst_Sbox_1_M15), .Z(SubBytesIns_Inst_Sbox_1_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_1_M16), 
        .B(SubBytesIns_Inst_Sbox_1_M13), .Z(SubBytesIns_Inst_Sbox_1_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_1_M17), 
        .B(SubBytesIns_Inst_Sbox_1_M15), .Z(SubBytesIns_Inst_Sbox_1_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_1_M18), 
        .B(SubBytesIns_Inst_Sbox_1_M13), .Z(SubBytesIns_Inst_Sbox_1_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_1_M19), 
        .B(SubBytesIns_Inst_Sbox_1_T25), .Z(SubBytesIns_Inst_Sbox_1_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_1_M22), 
        .B(SubBytesIns_Inst_Sbox_1_M23), .Z(SubBytesIns_Inst_Sbox_1_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M22), .A2(SubBytesIns_Inst_Sbox_1_M20), .ZN(SubBytesIns_Inst_Sbox_1_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_1_M21), 
        .B(SubBytesIns_Inst_Sbox_1_M25), .Z(SubBytesIns_Inst_Sbox_1_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_1_M20), 
        .B(SubBytesIns_Inst_Sbox_1_M21), .Z(SubBytesIns_Inst_Sbox_1_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_1_M23), 
        .B(SubBytesIns_Inst_Sbox_1_M25), .Z(SubBytesIns_Inst_Sbox_1_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M28), .A2(SubBytesIns_Inst_Sbox_1_M27), .ZN(SubBytesIns_Inst_Sbox_1_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M26), .A2(SubBytesIns_Inst_Sbox_1_M24), .ZN(SubBytesIns_Inst_Sbox_1_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M20), .A2(SubBytesIns_Inst_Sbox_1_M23), .ZN(SubBytesIns_Inst_Sbox_1_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M27), .A2(SubBytesIns_Inst_Sbox_1_M31), .ZN(SubBytesIns_Inst_Sbox_1_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_1_M27), 
        .B(SubBytesIns_Inst_Sbox_1_M25), .Z(SubBytesIns_Inst_Sbox_1_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M21), .A2(SubBytesIns_Inst_Sbox_1_M22), .ZN(SubBytesIns_Inst_Sbox_1_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M24), .A2(SubBytesIns_Inst_Sbox_1_M34), .ZN(SubBytesIns_Inst_Sbox_1_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_1_M24), 
        .B(SubBytesIns_Inst_Sbox_1_M25), .Z(SubBytesIns_Inst_Sbox_1_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_1_M21), 
        .B(SubBytesIns_Inst_Sbox_1_M29), .Z(SubBytesIns_Inst_Sbox_1_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_1_M32), 
        .B(SubBytesIns_Inst_Sbox_1_M33), .Z(SubBytesIns_Inst_Sbox_1_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_1_M23), 
        .B(SubBytesIns_Inst_Sbox_1_M30), .Z(SubBytesIns_Inst_Sbox_1_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_1_M35), 
        .B(SubBytesIns_Inst_Sbox_1_M36), .Z(SubBytesIns_Inst_Sbox_1_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_1_M38), 
        .B(SubBytesIns_Inst_Sbox_1_M40), .Z(SubBytesIns_Inst_Sbox_1_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_1_M37), 
        .B(SubBytesIns_Inst_Sbox_1_M39), .Z(SubBytesIns_Inst_Sbox_1_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_1_M37), 
        .B(SubBytesIns_Inst_Sbox_1_M38), .Z(SubBytesIns_Inst_Sbox_1_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_1_M39), 
        .B(SubBytesIns_Inst_Sbox_1_M40), .Z(SubBytesIns_Inst_Sbox_1_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_1_M42), 
        .B(SubBytesIns_Inst_Sbox_1_M41), .Z(SubBytesIns_Inst_Sbox_1_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M44), .A2(SubBytesIns_Inst_Sbox_1_T6), .ZN(SubBytesIns_Inst_Sbox_1_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M40), .A2(SubBytesIns_Inst_Sbox_1_T8), .ZN(SubBytesIns_Inst_Sbox_1_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M39), .A2(SubBytesInput[8]), .ZN(SubBytesIns_Inst_Sbox_1_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M43), .A2(SubBytesIns_Inst_Sbox_1_T16), .ZN(SubBytesIns_Inst_Sbox_1_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M38), .A2(SubBytesIns_Inst_Sbox_1_T9), .ZN(SubBytesIns_Inst_Sbox_1_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M37), .A2(SubBytesIns_Inst_Sbox_1_T17), .ZN(SubBytesIns_Inst_Sbox_1_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M42), .A2(SubBytesIns_Inst_Sbox_1_T15), .ZN(SubBytesIns_Inst_Sbox_1_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M45), .A2(SubBytesIns_Inst_Sbox_1_T27), .ZN(SubBytesIns_Inst_Sbox_1_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M41), .A2(SubBytesIns_Inst_Sbox_1_T10), .ZN(SubBytesIns_Inst_Sbox_1_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M44), .A2(SubBytesIns_Inst_Sbox_1_T13), .ZN(SubBytesIns_Inst_Sbox_1_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M40), .A2(SubBytesIns_Inst_Sbox_1_T23), .ZN(SubBytesIns_Inst_Sbox_1_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M39), .A2(SubBytesIns_Inst_Sbox_1_T19), .ZN(SubBytesIns_Inst_Sbox_1_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M43), .A2(SubBytesIns_Inst_Sbox_1_T3), .ZN(SubBytesIns_Inst_Sbox_1_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M38), .A2(SubBytesIns_Inst_Sbox_1_T22), .ZN(SubBytesIns_Inst_Sbox_1_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M37), .A2(SubBytesIns_Inst_Sbox_1_T20), .ZN(SubBytesIns_Inst_Sbox_1_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M42), .A2(SubBytesIns_Inst_Sbox_1_T1), .ZN(SubBytesIns_Inst_Sbox_1_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M45), .A2(SubBytesIns_Inst_Sbox_1_T4), .ZN(SubBytesIns_Inst_Sbox_1_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M41), .A2(SubBytesIns_Inst_Sbox_1_T2), .ZN(SubBytesIns_Inst_Sbox_1_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_1_M61), 
        .B(SubBytesIns_Inst_Sbox_1_M62), .Z(SubBytesIns_Inst_Sbox_1_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_1_M50), 
        .B(SubBytesIns_Inst_Sbox_1_M56), .Z(SubBytesIns_Inst_Sbox_1_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_1_M46), 
        .B(SubBytesIns_Inst_Sbox_1_M48), .Z(SubBytesIns_Inst_Sbox_1_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_1_M47), 
        .B(SubBytesIns_Inst_Sbox_1_M55), .Z(SubBytesIns_Inst_Sbox_1_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_1_M54), 
        .B(SubBytesIns_Inst_Sbox_1_M58), .Z(SubBytesIns_Inst_Sbox_1_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_1_M49), 
        .B(SubBytesIns_Inst_Sbox_1_M61), .Z(SubBytesIns_Inst_Sbox_1_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_1_M62), 
        .B(SubBytesIns_Inst_Sbox_1_L5), .Z(SubBytesIns_Inst_Sbox_1_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_1_M46), 
        .B(SubBytesIns_Inst_Sbox_1_L3), .Z(SubBytesIns_Inst_Sbox_1_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_1_M51), 
        .B(SubBytesIns_Inst_Sbox_1_M59), .Z(SubBytesIns_Inst_Sbox_1_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_1_M52), 
        .B(SubBytesIns_Inst_Sbox_1_M53), .Z(SubBytesIns_Inst_Sbox_1_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_1_M53), 
        .B(SubBytesIns_Inst_Sbox_1_L4), .Z(SubBytesIns_Inst_Sbox_1_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_1_M60), 
        .B(SubBytesIns_Inst_Sbox_1_L2), .Z(SubBytesIns_Inst_Sbox_1_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_1_M48), 
        .B(SubBytesIns_Inst_Sbox_1_M51), .Z(SubBytesIns_Inst_Sbox_1_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_1_M50), 
        .B(SubBytesIns_Inst_Sbox_1_L0), .Z(SubBytesIns_Inst_Sbox_1_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_1_M52), 
        .B(SubBytesIns_Inst_Sbox_1_M61), .Z(SubBytesIns_Inst_Sbox_1_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_1_M55), 
        .B(SubBytesIns_Inst_Sbox_1_L1), .Z(SubBytesIns_Inst_Sbox_1_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_1_M56), 
        .B(SubBytesIns_Inst_Sbox_1_L0), .Z(SubBytesIns_Inst_Sbox_1_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_1_M57), 
        .B(SubBytesIns_Inst_Sbox_1_L1), .Z(SubBytesIns_Inst_Sbox_1_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_1_M58), 
        .B(SubBytesIns_Inst_Sbox_1_L8), .Z(SubBytesIns_Inst_Sbox_1_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_1_M63), 
        .B(SubBytesIns_Inst_Sbox_1_L4), .Z(SubBytesIns_Inst_Sbox_1_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_1_L0), 
        .B(SubBytesIns_Inst_Sbox_1_L1), .Z(SubBytesIns_Inst_Sbox_1_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_1_L1), 
        .B(SubBytesIns_Inst_Sbox_1_L7), .Z(SubBytesIns_Inst_Sbox_1_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_1_L3), 
        .B(SubBytesIns_Inst_Sbox_1_L12), .Z(SubBytesIns_Inst_Sbox_1_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_1_L18), 
        .B(SubBytesIns_Inst_Sbox_1_L2), .Z(SubBytesIns_Inst_Sbox_1_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_1_L15), 
        .B(SubBytesIns_Inst_Sbox_1_L9), .Z(SubBytesIns_Inst_Sbox_1_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_1_L6), 
        .B(SubBytesIns_Inst_Sbox_1_L10), .Z(SubBytesIns_Inst_Sbox_1_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_1_L7), 
        .B(SubBytesIns_Inst_Sbox_1_L9), .Z(SubBytesIns_Inst_Sbox_1_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_1_L8), 
        .B(SubBytesIns_Inst_Sbox_1_L10), .Z(SubBytesIns_Inst_Sbox_1_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_1_L11), 
        .B(SubBytesIns_Inst_Sbox_1_L14), .Z(SubBytesIns_Inst_Sbox_1_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_1_L11), 
        .B(SubBytesIns_Inst_Sbox_1_L17), .Z(SubBytesIns_Inst_Sbox_1_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_1_L6), 
        .B(SubBytesIns_Inst_Sbox_1_L24), .Z(KeyExpansionIns_tmp[23]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_1_L16), 
        .B(SubBytesIns_Inst_Sbox_1_L26), .ZN(KeyExpansionIns_tmp[22]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_1_L19), 
        .B(SubBytesIns_Inst_Sbox_1_L28), .ZN(KeyExpansionIns_tmp[21]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_1_L6), 
        .B(SubBytesIns_Inst_Sbox_1_L21), .Z(KeyExpansionIns_tmp[20]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_1_L20), 
        .B(SubBytesIns_Inst_Sbox_1_L22), .Z(KeyExpansionIns_tmp[19]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_1_L25), 
        .B(SubBytesIns_Inst_Sbox_1_L29), .Z(KeyExpansionIns_tmp[18]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_1_L13), 
        .B(SubBytesIns_Inst_Sbox_1_L27), .ZN(KeyExpansionIns_tmp[17]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_1_L6), 
        .B(SubBytesIns_Inst_Sbox_1_L23), .ZN(KeyExpansionIns_tmp[16]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T1_U1 ( .A(SubBytesInput[23]), .B(
        SubBytesInput[20]), .Z(SubBytesIns_Inst_Sbox_2_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T2_U1 ( .A(SubBytesInput[23]), .B(
        SubBytesInput[18]), .Z(SubBytesIns_Inst_Sbox_2_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T3_U1 ( .A(SubBytesInput[23]), .B(
        SubBytesInput[17]), .Z(SubBytesIns_Inst_Sbox_2_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T4_U1 ( .A(SubBytesInput[20]), .B(
        SubBytesInput[18]), .Z(SubBytesIns_Inst_Sbox_2_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T5_U1 ( .A(SubBytesInput[19]), .B(
        SubBytesInput[17]), .Z(SubBytesIns_Inst_Sbox_2_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_2_T1), 
        .B(SubBytesIns_Inst_Sbox_2_T5), .Z(SubBytesIns_Inst_Sbox_2_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T7_U1 ( .A(SubBytesInput[22]), .B(
        SubBytesInput[21]), .Z(SubBytesIns_Inst_Sbox_2_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T8_U1 ( .A(SubBytesInput[16]), .B(
        SubBytesIns_Inst_Sbox_2_T6), .Z(SubBytesIns_Inst_Sbox_2_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T9_U1 ( .A(SubBytesInput[16]), .B(
        SubBytesIns_Inst_Sbox_2_T7), .Z(SubBytesIns_Inst_Sbox_2_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_2_T6), 
        .B(SubBytesIns_Inst_Sbox_2_T7), .Z(SubBytesIns_Inst_Sbox_2_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T11_U1 ( .A(SubBytesInput[22]), .B(
        SubBytesInput[18]), .Z(SubBytesIns_Inst_Sbox_2_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T12_U1 ( .A(SubBytesInput[21]), .B(
        SubBytesInput[18]), .Z(SubBytesIns_Inst_Sbox_2_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_2_T3), 
        .B(SubBytesIns_Inst_Sbox_2_T4), .Z(SubBytesIns_Inst_Sbox_2_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_2_T6), 
        .B(SubBytesIns_Inst_Sbox_2_T11), .Z(SubBytesIns_Inst_Sbox_2_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_2_T5), 
        .B(SubBytesIns_Inst_Sbox_2_T11), .Z(SubBytesIns_Inst_Sbox_2_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_2_T5), 
        .B(SubBytesIns_Inst_Sbox_2_T12), .Z(SubBytesIns_Inst_Sbox_2_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_2_T9), 
        .B(SubBytesIns_Inst_Sbox_2_T16), .Z(SubBytesIns_Inst_Sbox_2_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T18_U1 ( .A(SubBytesInput[20]), .B(
        SubBytesInput[16]), .Z(SubBytesIns_Inst_Sbox_2_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_2_T7), 
        .B(SubBytesIns_Inst_Sbox_2_T18), .Z(SubBytesIns_Inst_Sbox_2_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_2_T1), 
        .B(SubBytesIns_Inst_Sbox_2_T19), .Z(SubBytesIns_Inst_Sbox_2_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T21_U1 ( .A(SubBytesInput[17]), .B(
        SubBytesInput[16]), .Z(SubBytesIns_Inst_Sbox_2_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_2_T7), 
        .B(SubBytesIns_Inst_Sbox_2_T21), .Z(SubBytesIns_Inst_Sbox_2_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_2_T2), 
        .B(SubBytesIns_Inst_Sbox_2_T22), .Z(SubBytesIns_Inst_Sbox_2_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_2_T2), 
        .B(SubBytesIns_Inst_Sbox_2_T10), .Z(SubBytesIns_Inst_Sbox_2_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_2_T20), 
        .B(SubBytesIns_Inst_Sbox_2_T17), .Z(SubBytesIns_Inst_Sbox_2_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_2_T3), 
        .B(SubBytesIns_Inst_Sbox_2_T16), .Z(SubBytesIns_Inst_Sbox_2_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_2_T1), 
        .B(SubBytesIns_Inst_Sbox_2_T12), .Z(SubBytesIns_Inst_Sbox_2_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T13), 
        .A2(SubBytesIns_Inst_Sbox_2_T6), .ZN(SubBytesIns_Inst_Sbox_2_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T23), 
        .A2(SubBytesIns_Inst_Sbox_2_T8), .ZN(SubBytesIns_Inst_Sbox_2_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_2_T14), 
        .B(SubBytesIns_Inst_Sbox_2_M1), .Z(SubBytesIns_Inst_Sbox_2_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T19), 
        .A2(SubBytesInput[16]), .ZN(SubBytesIns_Inst_Sbox_2_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_2_M4), 
        .B(SubBytesIns_Inst_Sbox_2_M1), .Z(SubBytesIns_Inst_Sbox_2_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T3), 
        .A2(SubBytesIns_Inst_Sbox_2_T16), .ZN(SubBytesIns_Inst_Sbox_2_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T22), 
        .A2(SubBytesIns_Inst_Sbox_2_T9), .ZN(SubBytesIns_Inst_Sbox_2_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_2_T26), 
        .B(SubBytesIns_Inst_Sbox_2_M6), .Z(SubBytesIns_Inst_Sbox_2_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T20), 
        .A2(SubBytesIns_Inst_Sbox_2_T17), .ZN(SubBytesIns_Inst_Sbox_2_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_2_M9), 
        .B(SubBytesIns_Inst_Sbox_2_M6), .Z(SubBytesIns_Inst_Sbox_2_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T1), 
        .A2(SubBytesIns_Inst_Sbox_2_T15), .ZN(SubBytesIns_Inst_Sbox_2_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T4), 
        .A2(SubBytesIns_Inst_Sbox_2_T27), .ZN(SubBytesIns_Inst_Sbox_2_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_2_M12), 
        .B(SubBytesIns_Inst_Sbox_2_M11), .Z(SubBytesIns_Inst_Sbox_2_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T2), 
        .A2(SubBytesIns_Inst_Sbox_2_T10), .ZN(SubBytesIns_Inst_Sbox_2_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_2_M14), 
        .B(SubBytesIns_Inst_Sbox_2_M11), .Z(SubBytesIns_Inst_Sbox_2_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_2_M3), 
        .B(SubBytesIns_Inst_Sbox_2_M2), .Z(SubBytesIns_Inst_Sbox_2_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_2_M5), 
        .B(SubBytesIns_Inst_Sbox_2_T24), .Z(SubBytesIns_Inst_Sbox_2_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_2_M8), 
        .B(SubBytesIns_Inst_Sbox_2_M7), .Z(SubBytesIns_Inst_Sbox_2_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_2_M10), 
        .B(SubBytesIns_Inst_Sbox_2_M15), .Z(SubBytesIns_Inst_Sbox_2_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_2_M16), 
        .B(SubBytesIns_Inst_Sbox_2_M13), .Z(SubBytesIns_Inst_Sbox_2_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_2_M17), 
        .B(SubBytesIns_Inst_Sbox_2_M15), .Z(SubBytesIns_Inst_Sbox_2_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_2_M18), 
        .B(SubBytesIns_Inst_Sbox_2_M13), .Z(SubBytesIns_Inst_Sbox_2_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_2_M19), 
        .B(SubBytesIns_Inst_Sbox_2_T25), .Z(SubBytesIns_Inst_Sbox_2_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_2_M22), 
        .B(SubBytesIns_Inst_Sbox_2_M23), .Z(SubBytesIns_Inst_Sbox_2_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M22), .A2(SubBytesIns_Inst_Sbox_2_M20), .ZN(SubBytesIns_Inst_Sbox_2_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_2_M21), 
        .B(SubBytesIns_Inst_Sbox_2_M25), .Z(SubBytesIns_Inst_Sbox_2_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_2_M20), 
        .B(SubBytesIns_Inst_Sbox_2_M21), .Z(SubBytesIns_Inst_Sbox_2_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_2_M23), 
        .B(SubBytesIns_Inst_Sbox_2_M25), .Z(SubBytesIns_Inst_Sbox_2_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M28), .A2(SubBytesIns_Inst_Sbox_2_M27), .ZN(SubBytesIns_Inst_Sbox_2_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M26), .A2(SubBytesIns_Inst_Sbox_2_M24), .ZN(SubBytesIns_Inst_Sbox_2_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M20), .A2(SubBytesIns_Inst_Sbox_2_M23), .ZN(SubBytesIns_Inst_Sbox_2_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M27), .A2(SubBytesIns_Inst_Sbox_2_M31), .ZN(SubBytesIns_Inst_Sbox_2_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_2_M27), 
        .B(SubBytesIns_Inst_Sbox_2_M25), .Z(SubBytesIns_Inst_Sbox_2_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M21), .A2(SubBytesIns_Inst_Sbox_2_M22), .ZN(SubBytesIns_Inst_Sbox_2_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M24), .A2(SubBytesIns_Inst_Sbox_2_M34), .ZN(SubBytesIns_Inst_Sbox_2_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_2_M24), 
        .B(SubBytesIns_Inst_Sbox_2_M25), .Z(SubBytesIns_Inst_Sbox_2_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_2_M21), 
        .B(SubBytesIns_Inst_Sbox_2_M29), .Z(SubBytesIns_Inst_Sbox_2_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_2_M32), 
        .B(SubBytesIns_Inst_Sbox_2_M33), .Z(SubBytesIns_Inst_Sbox_2_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_2_M23), 
        .B(SubBytesIns_Inst_Sbox_2_M30), .Z(SubBytesIns_Inst_Sbox_2_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_2_M35), 
        .B(SubBytesIns_Inst_Sbox_2_M36), .Z(SubBytesIns_Inst_Sbox_2_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_2_M38), 
        .B(SubBytesIns_Inst_Sbox_2_M40), .Z(SubBytesIns_Inst_Sbox_2_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_2_M37), 
        .B(SubBytesIns_Inst_Sbox_2_M39), .Z(SubBytesIns_Inst_Sbox_2_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_2_M37), 
        .B(SubBytesIns_Inst_Sbox_2_M38), .Z(SubBytesIns_Inst_Sbox_2_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_2_M39), 
        .B(SubBytesIns_Inst_Sbox_2_M40), .Z(SubBytesIns_Inst_Sbox_2_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_2_M42), 
        .B(SubBytesIns_Inst_Sbox_2_M41), .Z(SubBytesIns_Inst_Sbox_2_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M44), .A2(SubBytesIns_Inst_Sbox_2_T6), .ZN(SubBytesIns_Inst_Sbox_2_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M40), .A2(SubBytesIns_Inst_Sbox_2_T8), .ZN(SubBytesIns_Inst_Sbox_2_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M39), .A2(SubBytesInput[16]), .ZN(SubBytesIns_Inst_Sbox_2_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M43), .A2(SubBytesIns_Inst_Sbox_2_T16), .ZN(SubBytesIns_Inst_Sbox_2_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M38), .A2(SubBytesIns_Inst_Sbox_2_T9), .ZN(SubBytesIns_Inst_Sbox_2_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M37), .A2(SubBytesIns_Inst_Sbox_2_T17), .ZN(SubBytesIns_Inst_Sbox_2_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M42), .A2(SubBytesIns_Inst_Sbox_2_T15), .ZN(SubBytesIns_Inst_Sbox_2_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M45), .A2(SubBytesIns_Inst_Sbox_2_T27), .ZN(SubBytesIns_Inst_Sbox_2_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M41), .A2(SubBytesIns_Inst_Sbox_2_T10), .ZN(SubBytesIns_Inst_Sbox_2_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M44), .A2(SubBytesIns_Inst_Sbox_2_T13), .ZN(SubBytesIns_Inst_Sbox_2_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M40), .A2(SubBytesIns_Inst_Sbox_2_T23), .ZN(SubBytesIns_Inst_Sbox_2_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M39), .A2(SubBytesIns_Inst_Sbox_2_T19), .ZN(SubBytesIns_Inst_Sbox_2_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M43), .A2(SubBytesIns_Inst_Sbox_2_T3), .ZN(SubBytesIns_Inst_Sbox_2_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M38), .A2(SubBytesIns_Inst_Sbox_2_T22), .ZN(SubBytesIns_Inst_Sbox_2_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M37), .A2(SubBytesIns_Inst_Sbox_2_T20), .ZN(SubBytesIns_Inst_Sbox_2_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M42), .A2(SubBytesIns_Inst_Sbox_2_T1), .ZN(SubBytesIns_Inst_Sbox_2_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M45), .A2(SubBytesIns_Inst_Sbox_2_T4), .ZN(SubBytesIns_Inst_Sbox_2_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M41), .A2(SubBytesIns_Inst_Sbox_2_T2), .ZN(SubBytesIns_Inst_Sbox_2_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_2_M61), 
        .B(SubBytesIns_Inst_Sbox_2_M62), .Z(SubBytesIns_Inst_Sbox_2_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_2_M50), 
        .B(SubBytesIns_Inst_Sbox_2_M56), .Z(SubBytesIns_Inst_Sbox_2_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_2_M46), 
        .B(SubBytesIns_Inst_Sbox_2_M48), .Z(SubBytesIns_Inst_Sbox_2_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_2_M47), 
        .B(SubBytesIns_Inst_Sbox_2_M55), .Z(SubBytesIns_Inst_Sbox_2_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_2_M54), 
        .B(SubBytesIns_Inst_Sbox_2_M58), .Z(SubBytesIns_Inst_Sbox_2_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_2_M49), 
        .B(SubBytesIns_Inst_Sbox_2_M61), .Z(SubBytesIns_Inst_Sbox_2_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_2_M62), 
        .B(SubBytesIns_Inst_Sbox_2_L5), .Z(SubBytesIns_Inst_Sbox_2_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_2_M46), 
        .B(SubBytesIns_Inst_Sbox_2_L3), .Z(SubBytesIns_Inst_Sbox_2_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_2_M51), 
        .B(SubBytesIns_Inst_Sbox_2_M59), .Z(SubBytesIns_Inst_Sbox_2_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_2_M52), 
        .B(SubBytesIns_Inst_Sbox_2_M53), .Z(SubBytesIns_Inst_Sbox_2_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_2_M53), 
        .B(SubBytesIns_Inst_Sbox_2_L4), .Z(SubBytesIns_Inst_Sbox_2_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_2_M60), 
        .B(SubBytesIns_Inst_Sbox_2_L2), .Z(SubBytesIns_Inst_Sbox_2_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_2_M48), 
        .B(SubBytesIns_Inst_Sbox_2_M51), .Z(SubBytesIns_Inst_Sbox_2_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_2_M50), 
        .B(SubBytesIns_Inst_Sbox_2_L0), .Z(SubBytesIns_Inst_Sbox_2_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_2_M52), 
        .B(SubBytesIns_Inst_Sbox_2_M61), .Z(SubBytesIns_Inst_Sbox_2_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_2_M55), 
        .B(SubBytesIns_Inst_Sbox_2_L1), .Z(SubBytesIns_Inst_Sbox_2_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_2_M56), 
        .B(SubBytesIns_Inst_Sbox_2_L0), .Z(SubBytesIns_Inst_Sbox_2_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_2_M57), 
        .B(SubBytesIns_Inst_Sbox_2_L1), .Z(SubBytesIns_Inst_Sbox_2_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_2_M58), 
        .B(SubBytesIns_Inst_Sbox_2_L8), .Z(SubBytesIns_Inst_Sbox_2_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_2_M63), 
        .B(SubBytesIns_Inst_Sbox_2_L4), .Z(SubBytesIns_Inst_Sbox_2_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_2_L0), 
        .B(SubBytesIns_Inst_Sbox_2_L1), .Z(SubBytesIns_Inst_Sbox_2_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_2_L1), 
        .B(SubBytesIns_Inst_Sbox_2_L7), .Z(SubBytesIns_Inst_Sbox_2_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_2_L3), 
        .B(SubBytesIns_Inst_Sbox_2_L12), .Z(SubBytesIns_Inst_Sbox_2_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_2_L18), 
        .B(SubBytesIns_Inst_Sbox_2_L2), .Z(SubBytesIns_Inst_Sbox_2_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_2_L15), 
        .B(SubBytesIns_Inst_Sbox_2_L9), .Z(SubBytesIns_Inst_Sbox_2_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_2_L6), 
        .B(SubBytesIns_Inst_Sbox_2_L10), .Z(SubBytesIns_Inst_Sbox_2_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_2_L7), 
        .B(SubBytesIns_Inst_Sbox_2_L9), .Z(SubBytesIns_Inst_Sbox_2_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_2_L8), 
        .B(SubBytesIns_Inst_Sbox_2_L10), .Z(SubBytesIns_Inst_Sbox_2_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_2_L11), 
        .B(SubBytesIns_Inst_Sbox_2_L14), .Z(SubBytesIns_Inst_Sbox_2_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_2_L11), 
        .B(SubBytesIns_Inst_Sbox_2_L17), .Z(SubBytesIns_Inst_Sbox_2_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_2_L6), 
        .B(SubBytesIns_Inst_Sbox_2_L24), .Z(KeyExpansionIns_tmp[15]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_2_L16), 
        .B(SubBytesIns_Inst_Sbox_2_L26), .ZN(KeyExpansionIns_tmp[14]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_2_L19), 
        .B(SubBytesIns_Inst_Sbox_2_L28), .ZN(KeyExpansionIns_tmp[13]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_2_L6), 
        .B(SubBytesIns_Inst_Sbox_2_L21), .Z(KeyExpansionIns_tmp[12]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_2_L20), 
        .B(SubBytesIns_Inst_Sbox_2_L22), .Z(KeyExpansionIns_tmp[11]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_2_L25), 
        .B(SubBytesIns_Inst_Sbox_2_L29), .Z(KeyExpansionIns_tmp[10]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_2_L13), 
        .B(SubBytesIns_Inst_Sbox_2_L27), .ZN(KeyExpansionIns_tmp[9]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_2_L6), 
        .B(SubBytesIns_Inst_Sbox_2_L23), .ZN(KeyExpansionIns_tmp[8]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T1_U1 ( .A(SubBytesInput[31]), .B(
        SubBytesInput[28]), .Z(SubBytesIns_Inst_Sbox_3_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T2_U1 ( .A(SubBytesInput[31]), .B(
        SubBytesInput[26]), .Z(SubBytesIns_Inst_Sbox_3_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T3_U1 ( .A(SubBytesInput[31]), .B(
        SubBytesInput[25]), .Z(SubBytesIns_Inst_Sbox_3_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T4_U1 ( .A(SubBytesInput[28]), .B(
        SubBytesInput[26]), .Z(SubBytesIns_Inst_Sbox_3_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T5_U1 ( .A(SubBytesInput[27]), .B(
        SubBytesInput[25]), .Z(SubBytesIns_Inst_Sbox_3_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_3_T1), 
        .B(SubBytesIns_Inst_Sbox_3_T5), .Z(SubBytesIns_Inst_Sbox_3_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T7_U1 ( .A(SubBytesInput[30]), .B(
        SubBytesInput[29]), .Z(SubBytesIns_Inst_Sbox_3_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T8_U1 ( .A(SubBytesInput[24]), .B(
        SubBytesIns_Inst_Sbox_3_T6), .Z(SubBytesIns_Inst_Sbox_3_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T9_U1 ( .A(SubBytesInput[24]), .B(
        SubBytesIns_Inst_Sbox_3_T7), .Z(SubBytesIns_Inst_Sbox_3_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_3_T6), 
        .B(SubBytesIns_Inst_Sbox_3_T7), .Z(SubBytesIns_Inst_Sbox_3_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T11_U1 ( .A(SubBytesInput[30]), .B(
        SubBytesInput[26]), .Z(SubBytesIns_Inst_Sbox_3_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T12_U1 ( .A(SubBytesInput[29]), .B(
        SubBytesInput[26]), .Z(SubBytesIns_Inst_Sbox_3_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_3_T3), 
        .B(SubBytesIns_Inst_Sbox_3_T4), .Z(SubBytesIns_Inst_Sbox_3_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_3_T6), 
        .B(SubBytesIns_Inst_Sbox_3_T11), .Z(SubBytesIns_Inst_Sbox_3_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_3_T5), 
        .B(SubBytesIns_Inst_Sbox_3_T11), .Z(SubBytesIns_Inst_Sbox_3_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_3_T5), 
        .B(SubBytesIns_Inst_Sbox_3_T12), .Z(SubBytesIns_Inst_Sbox_3_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_3_T9), 
        .B(SubBytesIns_Inst_Sbox_3_T16), .Z(SubBytesIns_Inst_Sbox_3_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T18_U1 ( .A(SubBytesInput[28]), .B(
        SubBytesInput[24]), .Z(SubBytesIns_Inst_Sbox_3_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_3_T7), 
        .B(SubBytesIns_Inst_Sbox_3_T18), .Z(SubBytesIns_Inst_Sbox_3_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_3_T1), 
        .B(SubBytesIns_Inst_Sbox_3_T19), .Z(SubBytesIns_Inst_Sbox_3_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T21_U1 ( .A(SubBytesInput[25]), .B(
        SubBytesInput[24]), .Z(SubBytesIns_Inst_Sbox_3_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_3_T7), 
        .B(SubBytesIns_Inst_Sbox_3_T21), .Z(SubBytesIns_Inst_Sbox_3_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_3_T2), 
        .B(SubBytesIns_Inst_Sbox_3_T22), .Z(SubBytesIns_Inst_Sbox_3_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_3_T2), 
        .B(SubBytesIns_Inst_Sbox_3_T10), .Z(SubBytesIns_Inst_Sbox_3_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_3_T20), 
        .B(SubBytesIns_Inst_Sbox_3_T17), .Z(SubBytesIns_Inst_Sbox_3_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_3_T3), 
        .B(SubBytesIns_Inst_Sbox_3_T16), .Z(SubBytesIns_Inst_Sbox_3_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_3_T1), 
        .B(SubBytesIns_Inst_Sbox_3_T12), .Z(SubBytesIns_Inst_Sbox_3_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T13), 
        .A2(SubBytesIns_Inst_Sbox_3_T6), .ZN(SubBytesIns_Inst_Sbox_3_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T23), 
        .A2(SubBytesIns_Inst_Sbox_3_T8), .ZN(SubBytesIns_Inst_Sbox_3_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_3_T14), 
        .B(SubBytesIns_Inst_Sbox_3_M1), .Z(SubBytesIns_Inst_Sbox_3_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T19), 
        .A2(SubBytesInput[24]), .ZN(SubBytesIns_Inst_Sbox_3_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_3_M4), 
        .B(SubBytesIns_Inst_Sbox_3_M1), .Z(SubBytesIns_Inst_Sbox_3_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T3), 
        .A2(SubBytesIns_Inst_Sbox_3_T16), .ZN(SubBytesIns_Inst_Sbox_3_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T22), 
        .A2(SubBytesIns_Inst_Sbox_3_T9), .ZN(SubBytesIns_Inst_Sbox_3_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_3_T26), 
        .B(SubBytesIns_Inst_Sbox_3_M6), .Z(SubBytesIns_Inst_Sbox_3_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T20), 
        .A2(SubBytesIns_Inst_Sbox_3_T17), .ZN(SubBytesIns_Inst_Sbox_3_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_3_M9), 
        .B(SubBytesIns_Inst_Sbox_3_M6), .Z(SubBytesIns_Inst_Sbox_3_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T1), 
        .A2(SubBytesIns_Inst_Sbox_3_T15), .ZN(SubBytesIns_Inst_Sbox_3_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T4), 
        .A2(SubBytesIns_Inst_Sbox_3_T27), .ZN(SubBytesIns_Inst_Sbox_3_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_3_M12), 
        .B(SubBytesIns_Inst_Sbox_3_M11), .Z(SubBytesIns_Inst_Sbox_3_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T2), 
        .A2(SubBytesIns_Inst_Sbox_3_T10), .ZN(SubBytesIns_Inst_Sbox_3_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_3_M14), 
        .B(SubBytesIns_Inst_Sbox_3_M11), .Z(SubBytesIns_Inst_Sbox_3_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_3_M3), 
        .B(SubBytesIns_Inst_Sbox_3_M2), .Z(SubBytesIns_Inst_Sbox_3_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_3_M5), 
        .B(SubBytesIns_Inst_Sbox_3_T24), .Z(SubBytesIns_Inst_Sbox_3_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_3_M8), 
        .B(SubBytesIns_Inst_Sbox_3_M7), .Z(SubBytesIns_Inst_Sbox_3_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_3_M10), 
        .B(SubBytesIns_Inst_Sbox_3_M15), .Z(SubBytesIns_Inst_Sbox_3_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_3_M16), 
        .B(SubBytesIns_Inst_Sbox_3_M13), .Z(SubBytesIns_Inst_Sbox_3_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_3_M17), 
        .B(SubBytesIns_Inst_Sbox_3_M15), .Z(SubBytesIns_Inst_Sbox_3_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_3_M18), 
        .B(SubBytesIns_Inst_Sbox_3_M13), .Z(SubBytesIns_Inst_Sbox_3_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_3_M19), 
        .B(SubBytesIns_Inst_Sbox_3_T25), .Z(SubBytesIns_Inst_Sbox_3_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_3_M22), 
        .B(SubBytesIns_Inst_Sbox_3_M23), .Z(SubBytesIns_Inst_Sbox_3_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M22), .A2(SubBytesIns_Inst_Sbox_3_M20), .ZN(SubBytesIns_Inst_Sbox_3_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_3_M21), 
        .B(SubBytesIns_Inst_Sbox_3_M25), .Z(SubBytesIns_Inst_Sbox_3_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_3_M20), 
        .B(SubBytesIns_Inst_Sbox_3_M21), .Z(SubBytesIns_Inst_Sbox_3_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_3_M23), 
        .B(SubBytesIns_Inst_Sbox_3_M25), .Z(SubBytesIns_Inst_Sbox_3_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M28), .A2(SubBytesIns_Inst_Sbox_3_M27), .ZN(SubBytesIns_Inst_Sbox_3_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M26), .A2(SubBytesIns_Inst_Sbox_3_M24), .ZN(SubBytesIns_Inst_Sbox_3_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M20), .A2(SubBytesIns_Inst_Sbox_3_M23), .ZN(SubBytesIns_Inst_Sbox_3_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M27), .A2(SubBytesIns_Inst_Sbox_3_M31), .ZN(SubBytesIns_Inst_Sbox_3_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_3_M27), 
        .B(SubBytesIns_Inst_Sbox_3_M25), .Z(SubBytesIns_Inst_Sbox_3_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M21), .A2(SubBytesIns_Inst_Sbox_3_M22), .ZN(SubBytesIns_Inst_Sbox_3_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M24), .A2(SubBytesIns_Inst_Sbox_3_M34), .ZN(SubBytesIns_Inst_Sbox_3_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_3_M24), 
        .B(SubBytesIns_Inst_Sbox_3_M25), .Z(SubBytesIns_Inst_Sbox_3_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_3_M21), 
        .B(SubBytesIns_Inst_Sbox_3_M29), .Z(SubBytesIns_Inst_Sbox_3_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_3_M32), 
        .B(SubBytesIns_Inst_Sbox_3_M33), .Z(SubBytesIns_Inst_Sbox_3_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_3_M23), 
        .B(SubBytesIns_Inst_Sbox_3_M30), .Z(SubBytesIns_Inst_Sbox_3_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_3_M35), 
        .B(SubBytesIns_Inst_Sbox_3_M36), .Z(SubBytesIns_Inst_Sbox_3_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_3_M38), 
        .B(SubBytesIns_Inst_Sbox_3_M40), .Z(SubBytesIns_Inst_Sbox_3_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_3_M37), 
        .B(SubBytesIns_Inst_Sbox_3_M39), .Z(SubBytesIns_Inst_Sbox_3_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_3_M37), 
        .B(SubBytesIns_Inst_Sbox_3_M38), .Z(SubBytesIns_Inst_Sbox_3_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_3_M39), 
        .B(SubBytesIns_Inst_Sbox_3_M40), .Z(SubBytesIns_Inst_Sbox_3_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_3_M42), 
        .B(SubBytesIns_Inst_Sbox_3_M41), .Z(SubBytesIns_Inst_Sbox_3_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M44), .A2(SubBytesIns_Inst_Sbox_3_T6), .ZN(SubBytesIns_Inst_Sbox_3_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M40), .A2(SubBytesIns_Inst_Sbox_3_T8), .ZN(SubBytesIns_Inst_Sbox_3_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M39), .A2(SubBytesInput[24]), .ZN(SubBytesIns_Inst_Sbox_3_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M43), .A2(SubBytesIns_Inst_Sbox_3_T16), .ZN(SubBytesIns_Inst_Sbox_3_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M38), .A2(SubBytesIns_Inst_Sbox_3_T9), .ZN(SubBytesIns_Inst_Sbox_3_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M37), .A2(SubBytesIns_Inst_Sbox_3_T17), .ZN(SubBytesIns_Inst_Sbox_3_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M42), .A2(SubBytesIns_Inst_Sbox_3_T15), .ZN(SubBytesIns_Inst_Sbox_3_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M45), .A2(SubBytesIns_Inst_Sbox_3_T27), .ZN(SubBytesIns_Inst_Sbox_3_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M41), .A2(SubBytesIns_Inst_Sbox_3_T10), .ZN(SubBytesIns_Inst_Sbox_3_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M44), .A2(SubBytesIns_Inst_Sbox_3_T13), .ZN(SubBytesIns_Inst_Sbox_3_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M40), .A2(SubBytesIns_Inst_Sbox_3_T23), .ZN(SubBytesIns_Inst_Sbox_3_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M39), .A2(SubBytesIns_Inst_Sbox_3_T19), .ZN(SubBytesIns_Inst_Sbox_3_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M43), .A2(SubBytesIns_Inst_Sbox_3_T3), .ZN(SubBytesIns_Inst_Sbox_3_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M38), .A2(SubBytesIns_Inst_Sbox_3_T22), .ZN(SubBytesIns_Inst_Sbox_3_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M37), .A2(SubBytesIns_Inst_Sbox_3_T20), .ZN(SubBytesIns_Inst_Sbox_3_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M42), .A2(SubBytesIns_Inst_Sbox_3_T1), .ZN(SubBytesIns_Inst_Sbox_3_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M45), .A2(SubBytesIns_Inst_Sbox_3_T4), .ZN(SubBytesIns_Inst_Sbox_3_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M41), .A2(SubBytesIns_Inst_Sbox_3_T2), .ZN(SubBytesIns_Inst_Sbox_3_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_3_M61), 
        .B(SubBytesIns_Inst_Sbox_3_M62), .Z(SubBytesIns_Inst_Sbox_3_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_3_M50), 
        .B(SubBytesIns_Inst_Sbox_3_M56), .Z(SubBytesIns_Inst_Sbox_3_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_3_M46), 
        .B(SubBytesIns_Inst_Sbox_3_M48), .Z(SubBytesIns_Inst_Sbox_3_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_3_M47), 
        .B(SubBytesIns_Inst_Sbox_3_M55), .Z(SubBytesIns_Inst_Sbox_3_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_3_M54), 
        .B(SubBytesIns_Inst_Sbox_3_M58), .Z(SubBytesIns_Inst_Sbox_3_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_3_M49), 
        .B(SubBytesIns_Inst_Sbox_3_M61), .Z(SubBytesIns_Inst_Sbox_3_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_3_M62), 
        .B(SubBytesIns_Inst_Sbox_3_L5), .Z(SubBytesIns_Inst_Sbox_3_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_3_M46), 
        .B(SubBytesIns_Inst_Sbox_3_L3), .Z(SubBytesIns_Inst_Sbox_3_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_3_M51), 
        .B(SubBytesIns_Inst_Sbox_3_M59), .Z(SubBytesIns_Inst_Sbox_3_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_3_M52), 
        .B(SubBytesIns_Inst_Sbox_3_M53), .Z(SubBytesIns_Inst_Sbox_3_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_3_M53), 
        .B(SubBytesIns_Inst_Sbox_3_L4), .Z(SubBytesIns_Inst_Sbox_3_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_3_M60), 
        .B(SubBytesIns_Inst_Sbox_3_L2), .Z(SubBytesIns_Inst_Sbox_3_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_3_M48), 
        .B(SubBytesIns_Inst_Sbox_3_M51), .Z(SubBytesIns_Inst_Sbox_3_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_3_M50), 
        .B(SubBytesIns_Inst_Sbox_3_L0), .Z(SubBytesIns_Inst_Sbox_3_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_3_M52), 
        .B(SubBytesIns_Inst_Sbox_3_M61), .Z(SubBytesIns_Inst_Sbox_3_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_3_M55), 
        .B(SubBytesIns_Inst_Sbox_3_L1), .Z(SubBytesIns_Inst_Sbox_3_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_3_M56), 
        .B(SubBytesIns_Inst_Sbox_3_L0), .Z(SubBytesIns_Inst_Sbox_3_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_3_M57), 
        .B(SubBytesIns_Inst_Sbox_3_L1), .Z(SubBytesIns_Inst_Sbox_3_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_3_M58), 
        .B(SubBytesIns_Inst_Sbox_3_L8), .Z(SubBytesIns_Inst_Sbox_3_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_3_M63), 
        .B(SubBytesIns_Inst_Sbox_3_L4), .Z(SubBytesIns_Inst_Sbox_3_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_3_L0), 
        .B(SubBytesIns_Inst_Sbox_3_L1), .Z(SubBytesIns_Inst_Sbox_3_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_3_L1), 
        .B(SubBytesIns_Inst_Sbox_3_L7), .Z(SubBytesIns_Inst_Sbox_3_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_3_L3), 
        .B(SubBytesIns_Inst_Sbox_3_L12), .Z(SubBytesIns_Inst_Sbox_3_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_3_L18), 
        .B(SubBytesIns_Inst_Sbox_3_L2), .Z(SubBytesIns_Inst_Sbox_3_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_3_L15), 
        .B(SubBytesIns_Inst_Sbox_3_L9), .Z(SubBytesIns_Inst_Sbox_3_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_3_L6), 
        .B(SubBytesIns_Inst_Sbox_3_L10), .Z(SubBytesIns_Inst_Sbox_3_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_3_L7), 
        .B(SubBytesIns_Inst_Sbox_3_L9), .Z(SubBytesIns_Inst_Sbox_3_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_3_L8), 
        .B(SubBytesIns_Inst_Sbox_3_L10), .Z(SubBytesIns_Inst_Sbox_3_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_3_L11), 
        .B(SubBytesIns_Inst_Sbox_3_L14), .Z(SubBytesIns_Inst_Sbox_3_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_3_L11), 
        .B(SubBytesIns_Inst_Sbox_3_L17), .Z(SubBytesIns_Inst_Sbox_3_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_3_L6), 
        .B(SubBytesIns_Inst_Sbox_3_L24), .Z(KeyExpansionIns_tmp[7]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_3_L16), 
        .B(SubBytesIns_Inst_Sbox_3_L26), .ZN(KeyExpansionIns_tmp[6]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_3_L19), 
        .B(SubBytesIns_Inst_Sbox_3_L28), .ZN(KeyExpansionIns_tmp[5]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_3_L6), 
        .B(SubBytesIns_Inst_Sbox_3_L21), .Z(KeyExpansionIns_tmp[4]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_3_L20), 
        .B(SubBytesIns_Inst_Sbox_3_L22), .Z(KeyExpansionIns_tmp[3]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_3_L25), 
        .B(SubBytesIns_Inst_Sbox_3_L29), .Z(KeyExpansionIns_tmp[2]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_3_L13), 
        .B(SubBytesIns_Inst_Sbox_3_L27), .ZN(KeyExpansionIns_tmp[1]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_3_L6), 
        .B(SubBytesIns_Inst_Sbox_3_L23), .ZN(KeyExpansionIns_tmp[0]) );
  XNOR2_X1 MixColumnsIns_U96 ( .A(MixColumnsIns_n64), .B(
        KeyExpansionIns_tmp[9]), .ZN(MixColumnsOutput[9]) );
  XNOR2_X1 MixColumnsIns_U95 ( .A(MixColumnsIns_n63), .B(MixColumnsIns_n62), 
        .ZN(MixColumnsIns_n64) );
  XNOR2_X1 MixColumnsIns_U94 ( .A(MixColumnsIns_n61), .B(MixColumnsIns_n60), 
        .ZN(MixColumnsOutput[8]) );
  XNOR2_X1 MixColumnsIns_U93 ( .A(MixColumnsIns_n59), .B(
        KeyExpansionIns_tmp[8]), .ZN(MixColumnsIns_n61) );
  XNOR2_X1 MixColumnsIns_U92 ( .A(MixColumnsIns_n58), .B(MixColumnsIns_n57), 
        .ZN(MixColumnsOutput[7]) );
  XNOR2_X1 MixColumnsIns_U91 ( .A(MixColumnsIns_n56), .B(
        KeyExpansionIns_tmp[23]), .ZN(MixColumnsIns_n58) );
  XNOR2_X1 MixColumnsIns_U90 ( .A(MixColumnsIns_n55), .B(MixColumnsIns_n54), 
        .ZN(MixColumnsOutput[6]) );
  XNOR2_X1 MixColumnsIns_U89 ( .A(MixColumnsIns_n53), .B(
        KeyExpansionIns_tmp[22]), .ZN(MixColumnsIns_n55) );
  XNOR2_X1 MixColumnsIns_U88 ( .A(MixColumnsIns_n52), .B(MixColumnsIns_n51), 
        .ZN(MixColumnsOutput[5]) );
  XNOR2_X1 MixColumnsIns_U87 ( .A(MixColumnsIns_n50), .B(
        KeyExpansionIns_tmp[21]), .ZN(MixColumnsIns_n52) );
  XNOR2_X1 MixColumnsIns_U86 ( .A(MixColumnsIns_n49), .B(MixColumnsIns_n48), 
        .ZN(MixColumnsOutput[4]) );
  XNOR2_X1 MixColumnsIns_U85 ( .A(MixColumnsIns_n47), .B(
        KeyExpansionIns_tmp[20]), .ZN(MixColumnsIns_n49) );
  XNOR2_X1 MixColumnsIns_U84 ( .A(MixColumnsIns_n46), .B(MixColumnsIns_n45), 
        .ZN(MixColumnsOutput[3]) );
  XNOR2_X1 MixColumnsIns_U83 ( .A(MixColumnsIns_n44), .B(
        KeyExpansionIns_tmp[19]), .ZN(MixColumnsIns_n46) );
  XNOR2_X1 MixColumnsIns_U82 ( .A(MixColumnsIns_n43), .B(MixColumnsIns_n57), 
        .ZN(MixColumnsOutput[31]) );
  XOR2_X1 MixColumnsIns_U81 ( .A(KeyExpansionIns_tmp[15]), .B(
        KeyExpansionIns_tmp[6]), .Z(MixColumnsIns_n57) );
  XNOR2_X1 MixColumnsIns_U80 ( .A(MixColumnsIns_DoubleBytes[0]), .B(
        MixColumnsIns_n42), .ZN(MixColumnsIns_n43) );
  XNOR2_X1 MixColumnsIns_U79 ( .A(MixColumnsIns_n41), .B(MixColumnsIns_n54), 
        .ZN(MixColumnsOutput[30]) );
  XOR2_X1 MixColumnsIns_U78 ( .A(KeyExpansionIns_tmp[14]), .B(
        KeyExpansionIns_tmp[5]), .Z(MixColumnsIns_n54) );
  XNOR2_X1 MixColumnsIns_U77 ( .A(MixColumnsIns_DoubleBytes[7]), .B(
        MixColumnsIns_n40), .ZN(MixColumnsIns_n41) );
  XNOR2_X1 MixColumnsIns_U76 ( .A(MixColumnsIns_n39), .B(MixColumnsIns_n38), 
        .ZN(MixColumnsOutput[2]) );
  XNOR2_X1 MixColumnsIns_U75 ( .A(MixColumnsIns_n37), .B(
        KeyExpansionIns_tmp[18]), .ZN(MixColumnsIns_n39) );
  XNOR2_X1 MixColumnsIns_U74 ( .A(MixColumnsIns_n36), .B(MixColumnsIns_n51), 
        .ZN(MixColumnsOutput[29]) );
  XOR2_X1 MixColumnsIns_U73 ( .A(KeyExpansionIns_tmp[13]), .B(
        KeyExpansionIns_tmp[4]), .Z(MixColumnsIns_n51) );
  XNOR2_X1 MixColumnsIns_U72 ( .A(MixColumnsIns_DoubleBytes[6]), .B(
        MixColumnsIns_n35), .ZN(MixColumnsIns_n36) );
  XNOR2_X1 MixColumnsIns_U71 ( .A(MixColumnsIns_n34), .B(MixColumnsIns_n48), 
        .ZN(MixColumnsOutput[28]) );
  XOR2_X1 MixColumnsIns_U70 ( .A(KeyExpansionIns_tmp[12]), .B(
        MixColumnsIns_DoubleBytes[28]), .Z(MixColumnsIns_n48) );
  XNOR2_X1 MixColumnsIns_U69 ( .A(MixColumnsIns_DoubleBytes[5]), .B(
        MixColumnsIns_n33), .ZN(MixColumnsIns_n34) );
  XNOR2_X1 MixColumnsIns_U68 ( .A(MixColumnsIns_n32), .B(MixColumnsIns_n45), 
        .ZN(MixColumnsOutput[27]) );
  XOR2_X1 MixColumnsIns_U67 ( .A(KeyExpansionIns_tmp[11]), .B(
        MixColumnsIns_DoubleBytes[27]), .Z(MixColumnsIns_n45) );
  XNOR2_X1 MixColumnsIns_U66 ( .A(SubBytesOutput[3]), .B(MixColumnsIns_n31), 
        .ZN(MixColumnsIns_n32) );
  XNOR2_X1 MixColumnsIns_U65 ( .A(MixColumnsIns_n30), .B(MixColumnsIns_n38), 
        .ZN(MixColumnsOutput[26]) );
  XOR2_X1 MixColumnsIns_U64 ( .A(KeyExpansionIns_tmp[10]), .B(
        KeyExpansionIns_tmp[1]), .Z(MixColumnsIns_n38) );
  XNOR2_X1 MixColumnsIns_U63 ( .A(SubBytesOutput[2]), .B(MixColumnsIns_n29), 
        .ZN(MixColumnsIns_n30) );
  XNOR2_X1 MixColumnsIns_U62 ( .A(MixColumnsIns_n28), .B(MixColumnsIns_n27), 
        .ZN(MixColumnsOutput[25]) );
  XNOR2_X1 MixColumnsIns_U61 ( .A(MixColumnsIns_DoubleBytes[2]), .B(
        MixColumnsIns_n26), .ZN(MixColumnsIns_n28) );
  XNOR2_X1 MixColumnsIns_U60 ( .A(MixColumnsIns_n25), .B(MixColumnsIns_n24), 
        .ZN(MixColumnsOutput[24]) );
  XNOR2_X1 MixColumnsIns_U59 ( .A(MixColumnsIns_n23), .B(SubBytesOutput[0]), 
        .ZN(MixColumnsIns_n25) );
  XNOR2_X1 MixColumnsIns_U58 ( .A(MixColumnsIns_n22), .B(MixColumnsIns_n42), 
        .ZN(MixColumnsOutput[23]) );
  XOR2_X1 MixColumnsIns_U57 ( .A(KeyExpansionIns_tmp[23]), .B(
        KeyExpansionIns_tmp[14]), .Z(MixColumnsIns_n42) );
  XNOR2_X1 MixColumnsIns_U56 ( .A(KeyExpansionIns_tmp[7]), .B(
        MixColumnsIns_n21), .ZN(MixColumnsIns_n22) );
  XNOR2_X1 MixColumnsIns_U55 ( .A(MixColumnsIns_n20), .B(MixColumnsIns_n40), 
        .ZN(MixColumnsOutput[22]) );
  XOR2_X1 MixColumnsIns_U54 ( .A(KeyExpansionIns_tmp[22]), .B(
        KeyExpansionIns_tmp[13]), .Z(MixColumnsIns_n40) );
  XNOR2_X1 MixColumnsIns_U53 ( .A(KeyExpansionIns_tmp[6]), .B(
        MixColumnsIns_n19), .ZN(MixColumnsIns_n20) );
  XNOR2_X1 MixColumnsIns_U52 ( .A(MixColumnsIns_n18), .B(MixColumnsIns_n35), 
        .ZN(MixColumnsOutput[21]) );
  XOR2_X1 MixColumnsIns_U51 ( .A(KeyExpansionIns_tmp[21]), .B(
        KeyExpansionIns_tmp[12]), .Z(MixColumnsIns_n35) );
  XNOR2_X1 MixColumnsIns_U50 ( .A(KeyExpansionIns_tmp[5]), .B(
        MixColumnsIns_n17), .ZN(MixColumnsIns_n18) );
  XNOR2_X1 MixColumnsIns_U49 ( .A(MixColumnsIns_n16), .B(MixColumnsIns_n33), 
        .ZN(MixColumnsOutput[20]) );
  XOR2_X1 MixColumnsIns_U48 ( .A(KeyExpansionIns_tmp[20]), .B(
        MixColumnsIns_DoubleBytes[20]), .Z(MixColumnsIns_n33) );
  XNOR2_X1 MixColumnsIns_U47 ( .A(KeyExpansionIns_tmp[4]), .B(
        MixColumnsIns_n15), .ZN(MixColumnsIns_n16) );
  XNOR2_X1 MixColumnsIns_U46 ( .A(MixColumnsIns_n14), .B(MixColumnsIns_n27), 
        .ZN(MixColumnsOutput[1]) );
  XOR2_X1 MixColumnsIns_U45 ( .A(KeyExpansionIns_tmp[9]), .B(
        MixColumnsIns_DoubleBytes[25]), .Z(MixColumnsIns_n27) );
  XNOR2_X1 MixColumnsIns_U44 ( .A(KeyExpansionIns_tmp[17]), .B(
        MixColumnsIns_n62), .ZN(MixColumnsIns_n14) );
  XOR2_X1 MixColumnsIns_U43 ( .A(KeyExpansionIns_tmp[1]), .B(
        MixColumnsIns_DoubleBytes[1]), .Z(MixColumnsIns_n62) );
  XNOR2_X1 MixColumnsIns_U42 ( .A(MixColumnsIns_n13), .B(MixColumnsIns_n31), 
        .ZN(MixColumnsOutput[19]) );
  XOR2_X1 MixColumnsIns_U41 ( .A(KeyExpansionIns_tmp[19]), .B(
        MixColumnsIns_DoubleBytes[19]), .Z(MixColumnsIns_n31) );
  XNOR2_X1 MixColumnsIns_U40 ( .A(KeyExpansionIns_tmp[3]), .B(
        MixColumnsIns_n12), .ZN(MixColumnsIns_n13) );
  XNOR2_X1 MixColumnsIns_U39 ( .A(MixColumnsIns_n11), .B(MixColumnsIns_n29), 
        .ZN(MixColumnsOutput[18]) );
  XOR2_X1 MixColumnsIns_U38 ( .A(KeyExpansionIns_tmp[18]), .B(
        KeyExpansionIns_tmp[9]), .Z(MixColumnsIns_n29) );
  XNOR2_X1 MixColumnsIns_U37 ( .A(KeyExpansionIns_tmp[2]), .B(
        MixColumnsIns_n10), .ZN(MixColumnsIns_n11) );
  XNOR2_X1 MixColumnsIns_U36 ( .A(MixColumnsIns_n9), .B(MixColumnsIns_n26), 
        .ZN(MixColumnsOutput[17]) );
  XOR2_X1 MixColumnsIns_U35 ( .A(MixColumnsIns_DoubleBytes[17]), .B(
        KeyExpansionIns_tmp[17]), .Z(MixColumnsIns_n26) );
  XNOR2_X1 MixColumnsIns_U34 ( .A(MixColumnsIns_n63), .B(
        KeyExpansionIns_tmp[1]), .ZN(MixColumnsIns_n9) );
  XOR2_X1 MixColumnsIns_U33 ( .A(MixColumnsIns_DoubleBytes[9]), .B(
        MixColumnsIns_DoubleBytes[2]), .Z(MixColumnsIns_n63) );
  XNOR2_X1 MixColumnsIns_U32 ( .A(MixColumnsIns_n8), .B(MixColumnsIns_n24), 
        .ZN(MixColumnsOutput[16]) );
  XOR2_X1 MixColumnsIns_U31 ( .A(KeyExpansionIns_tmp[16]), .B(
        KeyExpansionIns_tmp[15]), .Z(MixColumnsIns_n24) );
  XNOR2_X1 MixColumnsIns_U30 ( .A(KeyExpansionIns_tmp[0]), .B(
        MixColumnsIns_n60), .ZN(MixColumnsIns_n8) );
  XOR2_X1 MixColumnsIns_U29 ( .A(KeyExpansionIns_tmp[23]), .B(
        SubBytesOutput[0]), .Z(MixColumnsIns_n60) );
  XNOR2_X1 MixColumnsIns_U28 ( .A(MixColumnsIns_n7), .B(MixColumnsIns_n21), 
        .ZN(MixColumnsOutput[15]) );
  XOR2_X1 MixColumnsIns_U27 ( .A(MixColumnsIns_DoubleBytes[0]), .B(
        KeyExpansionIns_tmp[22]), .Z(MixColumnsIns_n21) );
  XNOR2_X1 MixColumnsIns_U26 ( .A(MixColumnsIns_n56), .B(
        KeyExpansionIns_tmp[15]), .ZN(MixColumnsIns_n7) );
  XOR2_X1 MixColumnsIns_U25 ( .A(MixColumnsIns_DoubleBytes[7]), .B(
        KeyExpansionIns_tmp[7]), .Z(MixColumnsIns_n56) );
  XNOR2_X1 MixColumnsIns_U24 ( .A(MixColumnsIns_n6), .B(MixColumnsIns_n19), 
        .ZN(MixColumnsOutput[14]) );
  XOR2_X1 MixColumnsIns_U23 ( .A(MixColumnsIns_DoubleBytes[7]), .B(
        KeyExpansionIns_tmp[21]), .Z(MixColumnsIns_n19) );
  XNOR2_X1 MixColumnsIns_U22 ( .A(MixColumnsIns_n53), .B(
        KeyExpansionIns_tmp[14]), .ZN(MixColumnsIns_n6) );
  XOR2_X1 MixColumnsIns_U21 ( .A(MixColumnsIns_DoubleBytes[6]), .B(
        KeyExpansionIns_tmp[6]), .Z(MixColumnsIns_n53) );
  XNOR2_X1 MixColumnsIns_U20 ( .A(MixColumnsIns_n5), .B(MixColumnsIns_n17), 
        .ZN(MixColumnsOutput[13]) );
  XOR2_X1 MixColumnsIns_U19 ( .A(MixColumnsIns_DoubleBytes[6]), .B(
        KeyExpansionIns_tmp[20]), .Z(MixColumnsIns_n17) );
  XNOR2_X1 MixColumnsIns_U18 ( .A(MixColumnsIns_n50), .B(
        KeyExpansionIns_tmp[13]), .ZN(MixColumnsIns_n5) );
  XOR2_X1 MixColumnsIns_U17 ( .A(MixColumnsIns_DoubleBytes[5]), .B(
        KeyExpansionIns_tmp[5]), .Z(MixColumnsIns_n50) );
  XNOR2_X1 MixColumnsIns_U16 ( .A(MixColumnsIns_n4), .B(MixColumnsIns_n15), 
        .ZN(MixColumnsOutput[12]) );
  XOR2_X1 MixColumnsIns_U15 ( .A(MixColumnsIns_DoubleBytes[5]), .B(
        MixColumnsIns_DoubleBytes[12]), .Z(MixColumnsIns_n15) );
  XNOR2_X1 MixColumnsIns_U14 ( .A(MixColumnsIns_n47), .B(
        KeyExpansionIns_tmp[12]), .ZN(MixColumnsIns_n4) );
  XOR2_X1 MixColumnsIns_U13 ( .A(MixColumnsIns_DoubleBytes[4]), .B(
        KeyExpansionIns_tmp[4]), .Z(MixColumnsIns_n47) );
  XNOR2_X1 MixColumnsIns_U12 ( .A(MixColumnsIns_n3), .B(MixColumnsIns_n12), 
        .ZN(MixColumnsOutput[11]) );
  XOR2_X1 MixColumnsIns_U11 ( .A(SubBytesOutput[3]), .B(
        MixColumnsIns_DoubleBytes[11]), .Z(MixColumnsIns_n12) );
  XNOR2_X1 MixColumnsIns_U10 ( .A(MixColumnsIns_n44), .B(
        KeyExpansionIns_tmp[11]), .ZN(MixColumnsIns_n3) );
  XOR2_X1 MixColumnsIns_U9 ( .A(MixColumnsIns_DoubleBytes[3]), .B(
        KeyExpansionIns_tmp[3]), .Z(MixColumnsIns_n44) );
  XNOR2_X1 MixColumnsIns_U8 ( .A(MixColumnsIns_n2), .B(MixColumnsIns_n10), 
        .ZN(MixColumnsOutput[10]) );
  XOR2_X1 MixColumnsIns_U7 ( .A(SubBytesOutput[2]), .B(KeyExpansionIns_tmp[17]), .Z(MixColumnsIns_n10) );
  XNOR2_X1 MixColumnsIns_U6 ( .A(MixColumnsIns_n37), .B(
        KeyExpansionIns_tmp[10]), .ZN(MixColumnsIns_n2) );
  XOR2_X1 MixColumnsIns_U5 ( .A(MixColumnsIns_DoubleBytes[2]), .B(
        KeyExpansionIns_tmp[2]), .Z(MixColumnsIns_n37) );
  XNOR2_X1 MixColumnsIns_U4 ( .A(MixColumnsIns_n1), .B(KeyExpansionIns_tmp[16]), .ZN(MixColumnsOutput[0]) );
  XNOR2_X1 MixColumnsIns_U3 ( .A(MixColumnsIns_n59), .B(MixColumnsIns_n23), 
        .ZN(MixColumnsIns_n1) );
  XOR2_X1 MixColumnsIns_U2 ( .A(KeyExpansionIns_tmp[8]), .B(
        KeyExpansionIns_tmp[7]), .Z(MixColumnsIns_n23) );
  XOR2_X1 MixColumnsIns_U1 ( .A(MixColumnsIns_DoubleBytes[0]), .B(
        KeyExpansionIns_tmp[0]), .Z(MixColumnsIns_n59) );
  XOR2_X1 MixColumnsIns_Mul2Inst_0_U3 ( .A(KeyExpansionIns_tmp[7]), .B(
        KeyExpansionIns_tmp[3]), .Z(MixColumnsIns_DoubleBytes[28]) );
  XOR2_X1 MixColumnsIns_Mul2Inst_0_U2 ( .A(KeyExpansionIns_tmp[7]), .B(
        KeyExpansionIns_tmp[2]), .Z(MixColumnsIns_DoubleBytes[27]) );
  XOR2_X1 MixColumnsIns_Mul2Inst_0_U1 ( .A(KeyExpansionIns_tmp[7]), .B(
        KeyExpansionIns_tmp[0]), .Z(MixColumnsIns_DoubleBytes[25]) );
  XOR2_X1 MixColumnsIns_Mul2Inst_1_U3 ( .A(KeyExpansionIns_tmp[15]), .B(
        KeyExpansionIns_tmp[11]), .Z(MixColumnsIns_DoubleBytes[20]) );
  XOR2_X1 MixColumnsIns_Mul2Inst_1_U2 ( .A(KeyExpansionIns_tmp[15]), .B(
        KeyExpansionIns_tmp[10]), .Z(MixColumnsIns_DoubleBytes[19]) );
  XOR2_X1 MixColumnsIns_Mul2Inst_1_U1 ( .A(KeyExpansionIns_tmp[15]), .B(
        KeyExpansionIns_tmp[8]), .Z(MixColumnsIns_DoubleBytes[17]) );
  XOR2_X1 MixColumnsIns_Mul2Inst_2_U3 ( .A(KeyExpansionIns_tmp[23]), .B(
        KeyExpansionIns_tmp[19]), .Z(MixColumnsIns_DoubleBytes[12]) );
  XOR2_X1 MixColumnsIns_Mul2Inst_2_U2 ( .A(KeyExpansionIns_tmp[23]), .B(
        KeyExpansionIns_tmp[18]), .Z(MixColumnsIns_DoubleBytes[11]) );
  XOR2_X1 MixColumnsIns_Mul2Inst_2_U1 ( .A(KeyExpansionIns_tmp[23]), .B(
        KeyExpansionIns_tmp[16]), .Z(MixColumnsIns_DoubleBytes[9]) );
  XOR2_X1 MixColumnsIns_Mul2Inst_3_U3 ( .A(MixColumnsIns_DoubleBytes[0]), .B(
        SubBytesOutput[3]), .Z(MixColumnsIns_DoubleBytes[4]) );
  XOR2_X1 MixColumnsIns_Mul2Inst_3_U2 ( .A(MixColumnsIns_DoubleBytes[0]), .B(
        SubBytesOutput[2]), .Z(MixColumnsIns_DoubleBytes[3]) );
  XOR2_X1 MixColumnsIns_Mul2Inst_3_U1 ( .A(MixColumnsIns_DoubleBytes[0]), .B(
        SubBytesOutput[0]), .Z(MixColumnsIns_DoubleBytes[1]) );
  INV_X1 MuxMCOut_U3 ( .A(LastRoundorDone), .ZN(MuxMCOut_n6) );
  INV_X1 MuxMCOut_U2 ( .A(MuxMCOut_n6), .ZN(MuxMCOut_n5) );
  INV_X1 MuxMCOut_U1 ( .A(MuxMCOut_n6), .ZN(MuxMCOut_n4) );
  MUX2_X1 MuxMCOut_mux_inst_0_U1 ( .A(MixColumnsOutput[0]), .B(
        SubBytesOutput[0]), .S(MuxMCOut_n5), .Z(ColumnOutput[0]) );
  MUX2_X1 MuxMCOut_mux_inst_1_U1 ( .A(MixColumnsOutput[1]), .B(
        MixColumnsIns_DoubleBytes[2]), .S(LastRoundorDone), .Z(ColumnOutput[1]) );
  MUX2_X1 MuxMCOut_mux_inst_2_U1 ( .A(MixColumnsOutput[2]), .B(
        SubBytesOutput[2]), .S(LastRoundorDone), .Z(ColumnOutput[2]) );
  MUX2_X1 MuxMCOut_mux_inst_3_U1 ( .A(MixColumnsOutput[3]), .B(
        SubBytesOutput[3]), .S(LastRoundorDone), .Z(ColumnOutput[3]) );
  MUX2_X1 MuxMCOut_mux_inst_4_U1 ( .A(MixColumnsOutput[4]), .B(
        MixColumnsIns_DoubleBytes[5]), .S(LastRoundorDone), .Z(ColumnOutput[4]) );
  MUX2_X1 MuxMCOut_mux_inst_5_U1 ( .A(MixColumnsOutput[5]), .B(
        MixColumnsIns_DoubleBytes[6]), .S(LastRoundorDone), .Z(ColumnOutput[5]) );
  MUX2_X1 MuxMCOut_mux_inst_6_U1 ( .A(MixColumnsOutput[6]), .B(
        MixColumnsIns_DoubleBytes[7]), .S(LastRoundorDone), .Z(ColumnOutput[6]) );
  MUX2_X1 MuxMCOut_mux_inst_7_U1 ( .A(MixColumnsOutput[7]), .B(
        MixColumnsIns_DoubleBytes[0]), .S(MuxMCOut_n4), .Z(ColumnOutput[7]) );
  MUX2_X1 MuxMCOut_mux_inst_8_U1 ( .A(MixColumnsOutput[8]), .B(
        KeyExpansionIns_tmp[16]), .S(MuxMCOut_n5), .Z(ColumnOutput[8]) );
  MUX2_X1 MuxMCOut_mux_inst_9_U1 ( .A(MixColumnsOutput[9]), .B(
        KeyExpansionIns_tmp[17]), .S(MuxMCOut_n5), .Z(ColumnOutput[9]) );
  MUX2_X1 MuxMCOut_mux_inst_10_U1 ( .A(MixColumnsOutput[10]), .B(
        KeyExpansionIns_tmp[18]), .S(MuxMCOut_n5), .Z(ColumnOutput[10]) );
  MUX2_X1 MuxMCOut_mux_inst_11_U1 ( .A(MixColumnsOutput[11]), .B(
        KeyExpansionIns_tmp[19]), .S(MuxMCOut_n5), .Z(ColumnOutput[11]) );
  MUX2_X1 MuxMCOut_mux_inst_12_U1 ( .A(MixColumnsOutput[12]), .B(
        KeyExpansionIns_tmp[20]), .S(MuxMCOut_n5), .Z(ColumnOutput[12]) );
  MUX2_X1 MuxMCOut_mux_inst_13_U1 ( .A(MixColumnsOutput[13]), .B(
        KeyExpansionIns_tmp[21]), .S(MuxMCOut_n5), .Z(ColumnOutput[13]) );
  MUX2_X1 MuxMCOut_mux_inst_14_U1 ( .A(MixColumnsOutput[14]), .B(
        KeyExpansionIns_tmp[22]), .S(MuxMCOut_n5), .Z(ColumnOutput[14]) );
  MUX2_X1 MuxMCOut_mux_inst_15_U1 ( .A(MixColumnsOutput[15]), .B(
        KeyExpansionIns_tmp[23]), .S(MuxMCOut_n5), .Z(ColumnOutput[15]) );
  MUX2_X1 MuxMCOut_mux_inst_16_U1 ( .A(MixColumnsOutput[16]), .B(
        KeyExpansionIns_tmp[8]), .S(MuxMCOut_n5), .Z(ColumnOutput[16]) );
  MUX2_X1 MuxMCOut_mux_inst_17_U1 ( .A(MixColumnsOutput[17]), .B(
        KeyExpansionIns_tmp[9]), .S(MuxMCOut_n5), .Z(ColumnOutput[17]) );
  MUX2_X1 MuxMCOut_mux_inst_18_U1 ( .A(MixColumnsOutput[18]), .B(
        KeyExpansionIns_tmp[10]), .S(MuxMCOut_n5), .Z(ColumnOutput[18]) );
  MUX2_X1 MuxMCOut_mux_inst_19_U1 ( .A(MixColumnsOutput[19]), .B(
        KeyExpansionIns_tmp[11]), .S(MuxMCOut_n5), .Z(ColumnOutput[19]) );
  MUX2_X1 MuxMCOut_mux_inst_20_U1 ( .A(MixColumnsOutput[20]), .B(
        KeyExpansionIns_tmp[12]), .S(MuxMCOut_n4), .Z(ColumnOutput[20]) );
  MUX2_X1 MuxMCOut_mux_inst_21_U1 ( .A(MixColumnsOutput[21]), .B(
        KeyExpansionIns_tmp[13]), .S(MuxMCOut_n4), .Z(ColumnOutput[21]) );
  MUX2_X1 MuxMCOut_mux_inst_22_U1 ( .A(MixColumnsOutput[22]), .B(
        KeyExpansionIns_tmp[14]), .S(MuxMCOut_n4), .Z(ColumnOutput[22]) );
  MUX2_X1 MuxMCOut_mux_inst_23_U1 ( .A(MixColumnsOutput[23]), .B(
        KeyExpansionIns_tmp[15]), .S(MuxMCOut_n4), .Z(ColumnOutput[23]) );
  MUX2_X1 MuxMCOut_mux_inst_24_U1 ( .A(MixColumnsOutput[24]), .B(
        KeyExpansionIns_tmp[0]), .S(MuxMCOut_n4), .Z(ColumnOutput[24]) );
  MUX2_X1 MuxMCOut_mux_inst_25_U1 ( .A(MixColumnsOutput[25]), .B(
        KeyExpansionIns_tmp[1]), .S(MuxMCOut_n4), .Z(ColumnOutput[25]) );
  MUX2_X1 MuxMCOut_mux_inst_26_U1 ( .A(MixColumnsOutput[26]), .B(
        KeyExpansionIns_tmp[2]), .S(MuxMCOut_n4), .Z(ColumnOutput[26]) );
  MUX2_X1 MuxMCOut_mux_inst_27_U1 ( .A(MixColumnsOutput[27]), .B(
        KeyExpansionIns_tmp[3]), .S(MuxMCOut_n4), .Z(ColumnOutput[27]) );
  MUX2_X1 MuxMCOut_mux_inst_28_U1 ( .A(MixColumnsOutput[28]), .B(
        KeyExpansionIns_tmp[4]), .S(MuxMCOut_n4), .Z(ColumnOutput[28]) );
  MUX2_X1 MuxMCOut_mux_inst_29_U1 ( .A(MixColumnsOutput[29]), .B(
        KeyExpansionIns_tmp[5]), .S(MuxMCOut_n4), .Z(ColumnOutput[29]) );
  MUX2_X1 MuxMCOut_mux_inst_30_U1 ( .A(MixColumnsOutput[30]), .B(
        KeyExpansionIns_tmp[6]), .S(MuxMCOut_n4), .Z(ColumnOutput[30]) );
  MUX2_X1 MuxMCOut_mux_inst_31_U1 ( .A(MixColumnsOutput[31]), .B(
        KeyExpansionIns_tmp[7]), .S(MuxMCOut_n4), .Z(ColumnOutput[31]) );
  INV_X1 MuxRound_U7 ( .A(AKSRnotDone), .ZN(MuxRound_n19) );
  INV_X1 MuxRound_U6 ( .A(MuxRound_n19), .ZN(MuxRound_n16) );
  INV_X1 MuxRound_U5 ( .A(MuxRound_n19), .ZN(MuxRound_n14) );
  INV_X1 MuxRound_U4 ( .A(MuxRound_n19), .ZN(MuxRound_n13) );
  INV_X1 MuxRound_U3 ( .A(MuxRound_n19), .ZN(MuxRound_n15) );
  INV_X1 MuxRound_U2 ( .A(MuxRound_n19), .ZN(MuxRound_n18) );
  INV_X1 MuxRound_U1 ( .A(MuxRound_n19), .ZN(MuxRound_n17) );
  MUX2_X1 MuxRound_mux_inst_0_U1 ( .A(ColumnOutput[0]), .B(ShiftRowsOutput[0]), 
        .S(AKSRnotDone), .Z(RoundOutput[0]) );
  MUX2_X1 MuxRound_mux_inst_1_U1 ( .A(ColumnOutput[1]), .B(ShiftRowsOutput[1]), 
        .S(MuxRound_n13), .Z(RoundOutput[1]) );
  MUX2_X1 MuxRound_mux_inst_2_U1 ( .A(ColumnOutput[2]), .B(ShiftRowsOutput[2]), 
        .S(MuxRound_n14), .Z(RoundOutput[2]) );
  MUX2_X1 MuxRound_mux_inst_3_U1 ( .A(ColumnOutput[3]), .B(ShiftRowsOutput[3]), 
        .S(MuxRound_n15), .Z(RoundOutput[3]) );
  MUX2_X1 MuxRound_mux_inst_4_U1 ( .A(ColumnOutput[4]), .B(ShiftRowsOutput[4]), 
        .S(MuxRound_n16), .Z(RoundOutput[4]) );
  MUX2_X1 MuxRound_mux_inst_5_U1 ( .A(ColumnOutput[5]), .B(ShiftRowsOutput[5]), 
        .S(MuxRound_n17), .Z(RoundOutput[5]) );
  MUX2_X1 MuxRound_mux_inst_6_U1 ( .A(ColumnOutput[6]), .B(ShiftRowsOutput[6]), 
        .S(MuxRound_n18), .Z(RoundOutput[6]) );
  MUX2_X1 MuxRound_mux_inst_7_U1 ( .A(ColumnOutput[7]), .B(ShiftRowsOutput[7]), 
        .S(MuxRound_n13), .Z(RoundOutput[7]) );
  MUX2_X1 MuxRound_mux_inst_8_U1 ( .A(ColumnOutput[8]), .B(ShiftRowsOutput[8]), 
        .S(MuxRound_n16), .Z(RoundOutput[8]) );
  MUX2_X1 MuxRound_mux_inst_9_U1 ( .A(ColumnOutput[9]), .B(ShiftRowsOutput[9]), 
        .S(MuxRound_n13), .Z(RoundOutput[9]) );
  MUX2_X1 MuxRound_mux_inst_10_U1 ( .A(ColumnOutput[10]), .B(
        ShiftRowsOutput[10]), .S(AKSRnotDone), .Z(RoundOutput[10]) );
  MUX2_X1 MuxRound_mux_inst_11_U1 ( .A(ColumnOutput[11]), .B(
        ShiftRowsOutput[11]), .S(AKSRnotDone), .Z(RoundOutput[11]) );
  MUX2_X1 MuxRound_mux_inst_12_U1 ( .A(ColumnOutput[12]), .B(
        ShiftRowsOutput[12]), .S(AKSRnotDone), .Z(RoundOutput[12]) );
  MUX2_X1 MuxRound_mux_inst_13_U1 ( .A(ColumnOutput[13]), .B(
        ShiftRowsOutput[13]), .S(AKSRnotDone), .Z(RoundOutput[13]) );
  MUX2_X1 MuxRound_mux_inst_14_U1 ( .A(ColumnOutput[14]), .B(
        ShiftRowsOutput[14]), .S(AKSRnotDone), .Z(RoundOutput[14]) );
  MUX2_X1 MuxRound_mux_inst_15_U1 ( .A(ColumnOutput[15]), .B(
        ShiftRowsOutput[15]), .S(AKSRnotDone), .Z(RoundOutput[15]) );
  MUX2_X1 MuxRound_mux_inst_16_U1 ( .A(ColumnOutput[16]), .B(
        ShiftRowsOutput[16]), .S(AKSRnotDone), .Z(RoundOutput[16]) );
  MUX2_X1 MuxRound_mux_inst_17_U1 ( .A(ColumnOutput[17]), .B(
        ShiftRowsOutput[17]), .S(AKSRnotDone), .Z(RoundOutput[17]) );
  MUX2_X1 MuxRound_mux_inst_18_U1 ( .A(ColumnOutput[18]), .B(
        ShiftRowsOutput[18]), .S(AKSRnotDone), .Z(RoundOutput[18]) );
  MUX2_X1 MuxRound_mux_inst_19_U1 ( .A(ColumnOutput[19]), .B(
        ShiftRowsOutput[19]), .S(AKSRnotDone), .Z(RoundOutput[19]) );
  MUX2_X1 MuxRound_mux_inst_20_U1 ( .A(ColumnOutput[20]), .B(
        ShiftRowsOutput[20]), .S(MuxRound_n14), .Z(RoundOutput[20]) );
  MUX2_X1 MuxRound_mux_inst_21_U1 ( .A(ColumnOutput[21]), .B(
        ShiftRowsOutput[21]), .S(MuxRound_n15), .Z(RoundOutput[21]) );
  MUX2_X1 MuxRound_mux_inst_22_U1 ( .A(ColumnOutput[22]), .B(
        ShiftRowsOutput[22]), .S(MuxRound_n16), .Z(RoundOutput[22]) );
  MUX2_X1 MuxRound_mux_inst_23_U1 ( .A(ColumnOutput[23]), .B(
        ShiftRowsOutput[23]), .S(MuxRound_n17), .Z(RoundOutput[23]) );
  MUX2_X1 MuxRound_mux_inst_24_U1 ( .A(ColumnOutput[24]), .B(
        ShiftRowsOutput[24]), .S(MuxRound_n18), .Z(RoundOutput[24]) );
  MUX2_X1 MuxRound_mux_inst_25_U1 ( .A(ColumnOutput[25]), .B(
        ShiftRowsOutput[25]), .S(MuxRound_n16), .Z(RoundOutput[25]) );
  MUX2_X1 MuxRound_mux_inst_26_U1 ( .A(ColumnOutput[26]), .B(
        ShiftRowsOutput[26]), .S(MuxRound_n17), .Z(RoundOutput[26]) );
  MUX2_X1 MuxRound_mux_inst_27_U1 ( .A(ColumnOutput[27]), .B(
        ShiftRowsOutput[27]), .S(AKSRnotDone), .Z(RoundOutput[27]) );
  MUX2_X1 MuxRound_mux_inst_28_U1 ( .A(ColumnOutput[28]), .B(
        ShiftRowsOutput[28]), .S(AKSRnotDone), .Z(RoundOutput[28]) );
  MUX2_X1 MuxRound_mux_inst_29_U1 ( .A(ColumnOutput[29]), .B(
        ShiftRowsOutput[29]), .S(MuxRound_n13), .Z(RoundOutput[29]) );
  MUX2_X1 MuxRound_mux_inst_30_U1 ( .A(ColumnOutput[30]), .B(
        ShiftRowsOutput[30]), .S(MuxRound_n14), .Z(RoundOutput[30]) );
  MUX2_X1 MuxRound_mux_inst_31_U1 ( .A(ColumnOutput[31]), .B(
        ShiftRowsOutput[31]), .S(MuxRound_n15), .Z(RoundOutput[31]) );
  MUX2_X1 MuxRound_mux_inst_32_U1 ( .A(ciphertext[32]), .B(ShiftRowsOutput[32]), .S(MuxRound_n18), .Z(RoundOutput[32]) );
  MUX2_X1 MuxRound_mux_inst_33_U1 ( .A(ciphertext[33]), .B(ShiftRowsOutput[33]), .S(MuxRound_n17), .Z(RoundOutput[33]) );
  MUX2_X1 MuxRound_mux_inst_34_U1 ( .A(ciphertext[34]), .B(ShiftRowsOutput[34]), .S(MuxRound_n13), .Z(RoundOutput[34]) );
  MUX2_X1 MuxRound_mux_inst_35_U1 ( .A(ciphertext[35]), .B(ShiftRowsOutput[35]), .S(MuxRound_n14), .Z(RoundOutput[35]) );
  MUX2_X1 MuxRound_mux_inst_36_U1 ( .A(ciphertext[36]), .B(ShiftRowsOutput[36]), .S(MuxRound_n15), .Z(RoundOutput[36]) );
  MUX2_X1 MuxRound_mux_inst_37_U1 ( .A(ciphertext[37]), .B(ShiftRowsOutput[37]), .S(MuxRound_n16), .Z(RoundOutput[37]) );
  MUX2_X1 MuxRound_mux_inst_38_U1 ( .A(ciphertext[38]), .B(ShiftRowsOutput[38]), .S(MuxRound_n17), .Z(RoundOutput[38]) );
  MUX2_X1 MuxRound_mux_inst_39_U1 ( .A(ciphertext[39]), .B(ShiftRowsOutput[39]), .S(MuxRound_n18), .Z(RoundOutput[39]) );
  MUX2_X1 MuxRound_mux_inst_40_U1 ( .A(ciphertext[72]), .B(ShiftRowsOutput[40]), .S(MuxRound_n18), .Z(RoundOutput[40]) );
  MUX2_X1 MuxRound_mux_inst_41_U1 ( .A(ciphertext[73]), .B(ShiftRowsOutput[41]), .S(MuxRound_n13), .Z(RoundOutput[41]) );
  MUX2_X1 MuxRound_mux_inst_42_U1 ( .A(ciphertext[74]), .B(ShiftRowsOutput[42]), .S(MuxRound_n14), .Z(RoundOutput[42]) );
  MUX2_X1 MuxRound_mux_inst_43_U1 ( .A(ciphertext[75]), .B(ShiftRowsOutput[43]), .S(MuxRound_n15), .Z(RoundOutput[43]) );
  MUX2_X1 MuxRound_mux_inst_44_U1 ( .A(ciphertext[76]), .B(ShiftRowsOutput[44]), .S(MuxRound_n13), .Z(RoundOutput[44]) );
  MUX2_X1 MuxRound_mux_inst_45_U1 ( .A(ciphertext[77]), .B(ShiftRowsOutput[45]), .S(MuxRound_n14), .Z(RoundOutput[45]) );
  MUX2_X1 MuxRound_mux_inst_46_U1 ( .A(ciphertext[78]), .B(ShiftRowsOutput[46]), .S(MuxRound_n15), .Z(RoundOutput[46]) );
  MUX2_X1 MuxRound_mux_inst_47_U1 ( .A(ciphertext[79]), .B(ShiftRowsOutput[47]), .S(MuxRound_n16), .Z(RoundOutput[47]) );
  MUX2_X1 MuxRound_mux_inst_48_U1 ( .A(ciphertext[112]), .B(
        ShiftRowsOutput[48]), .S(MuxRound_n17), .Z(RoundOutput[48]) );
  MUX2_X1 MuxRound_mux_inst_49_U1 ( .A(ciphertext[113]), .B(
        ShiftRowsOutput[49]), .S(MuxRound_n18), .Z(RoundOutput[49]) );
  MUX2_X1 MuxRound_mux_inst_50_U1 ( .A(ciphertext[114]), .B(
        ShiftRowsOutput[50]), .S(MuxRound_n13), .Z(RoundOutput[50]) );
  MUX2_X1 MuxRound_mux_inst_51_U1 ( .A(ciphertext[115]), .B(
        ShiftRowsOutput[51]), .S(MuxRound_n14), .Z(RoundOutput[51]) );
  MUX2_X1 MuxRound_mux_inst_52_U1 ( .A(ciphertext[116]), .B(
        ShiftRowsOutput[52]), .S(MuxRound_n15), .Z(RoundOutput[52]) );
  MUX2_X1 MuxRound_mux_inst_53_U1 ( .A(ciphertext[117]), .B(
        ShiftRowsOutput[53]), .S(MuxRound_n16), .Z(RoundOutput[53]) );
  MUX2_X1 MuxRound_mux_inst_54_U1 ( .A(ciphertext[118]), .B(
        ShiftRowsOutput[54]), .S(MuxRound_n17), .Z(RoundOutput[54]) );
  MUX2_X1 MuxRound_mux_inst_55_U1 ( .A(ciphertext[119]), .B(
        ShiftRowsOutput[55]), .S(MuxRound_n18), .Z(RoundOutput[55]) );
  MUX2_X1 MuxRound_mux_inst_56_U1 ( .A(ciphertext[24]), .B(ShiftRowsOutput[56]), .S(MuxRound_n18), .Z(RoundOutput[56]) );
  MUX2_X1 MuxRound_mux_inst_57_U1 ( .A(ciphertext[25]), .B(ShiftRowsOutput[57]), .S(MuxRound_n18), .Z(RoundOutput[57]) );
  MUX2_X1 MuxRound_mux_inst_58_U1 ( .A(ciphertext[26]), .B(ShiftRowsOutput[58]), .S(MuxRound_n18), .Z(RoundOutput[58]) );
  MUX2_X1 MuxRound_mux_inst_59_U1 ( .A(ciphertext[27]), .B(ShiftRowsOutput[59]), .S(MuxRound_n18), .Z(RoundOutput[59]) );
  MUX2_X1 MuxRound_mux_inst_60_U1 ( .A(ciphertext[28]), .B(ShiftRowsOutput[60]), .S(MuxRound_n18), .Z(RoundOutput[60]) );
  MUX2_X1 MuxRound_mux_inst_61_U1 ( .A(ciphertext[29]), .B(ShiftRowsOutput[61]), .S(MuxRound_n18), .Z(RoundOutput[61]) );
  MUX2_X1 MuxRound_mux_inst_62_U1 ( .A(ciphertext[30]), .B(ShiftRowsOutput[62]), .S(MuxRound_n18), .Z(RoundOutput[62]) );
  MUX2_X1 MuxRound_mux_inst_63_U1 ( .A(ciphertext[31]), .B(ShiftRowsOutput[63]), .S(MuxRound_n18), .Z(RoundOutput[63]) );
  MUX2_X1 MuxRound_mux_inst_64_U1 ( .A(ciphertext[64]), .B(ShiftRowsOutput[64]), .S(MuxRound_n18), .Z(RoundOutput[64]) );
  MUX2_X1 MuxRound_mux_inst_65_U1 ( .A(ciphertext[65]), .B(ShiftRowsOutput[65]), .S(MuxRound_n18), .Z(RoundOutput[65]) );
  MUX2_X1 MuxRound_mux_inst_66_U1 ( .A(ciphertext[66]), .B(ShiftRowsOutput[66]), .S(MuxRound_n18), .Z(RoundOutput[66]) );
  MUX2_X1 MuxRound_mux_inst_67_U1 ( .A(ciphertext[67]), .B(ShiftRowsOutput[67]), .S(MuxRound_n18), .Z(RoundOutput[67]) );
  MUX2_X1 MuxRound_mux_inst_68_U1 ( .A(ciphertext[68]), .B(ShiftRowsOutput[68]), .S(MuxRound_n17), .Z(RoundOutput[68]) );
  MUX2_X1 MuxRound_mux_inst_69_U1 ( .A(ciphertext[69]), .B(ShiftRowsOutput[69]), .S(MuxRound_n17), .Z(RoundOutput[69]) );
  MUX2_X1 MuxRound_mux_inst_70_U1 ( .A(ciphertext[70]), .B(ShiftRowsOutput[70]), .S(MuxRound_n17), .Z(RoundOutput[70]) );
  MUX2_X1 MuxRound_mux_inst_71_U1 ( .A(ciphertext[71]), .B(ShiftRowsOutput[71]), .S(MuxRound_n17), .Z(RoundOutput[71]) );
  MUX2_X1 MuxRound_mux_inst_72_U1 ( .A(ciphertext[104]), .B(
        ShiftRowsOutput[72]), .S(MuxRound_n17), .Z(RoundOutput[72]) );
  MUX2_X1 MuxRound_mux_inst_73_U1 ( .A(ciphertext[105]), .B(
        ShiftRowsOutput[73]), .S(MuxRound_n17), .Z(RoundOutput[73]) );
  MUX2_X1 MuxRound_mux_inst_74_U1 ( .A(ciphertext[106]), .B(
        ShiftRowsOutput[74]), .S(MuxRound_n17), .Z(RoundOutput[74]) );
  MUX2_X1 MuxRound_mux_inst_75_U1 ( .A(ciphertext[107]), .B(
        ShiftRowsOutput[75]), .S(MuxRound_n17), .Z(RoundOutput[75]) );
  MUX2_X1 MuxRound_mux_inst_76_U1 ( .A(ciphertext[108]), .B(
        ShiftRowsOutput[76]), .S(MuxRound_n17), .Z(RoundOutput[76]) );
  MUX2_X1 MuxRound_mux_inst_77_U1 ( .A(ciphertext[109]), .B(
        ShiftRowsOutput[77]), .S(MuxRound_n17), .Z(RoundOutput[77]) );
  MUX2_X1 MuxRound_mux_inst_78_U1 ( .A(ciphertext[110]), .B(
        ShiftRowsOutput[78]), .S(MuxRound_n17), .Z(RoundOutput[78]) );
  MUX2_X1 MuxRound_mux_inst_79_U1 ( .A(ciphertext[111]), .B(
        ShiftRowsOutput[79]), .S(MuxRound_n17), .Z(RoundOutput[79]) );
  MUX2_X1 MuxRound_mux_inst_80_U1 ( .A(ciphertext[16]), .B(ShiftRowsOutput[80]), .S(MuxRound_n16), .Z(RoundOutput[80]) );
  MUX2_X1 MuxRound_mux_inst_81_U1 ( .A(ciphertext[17]), .B(ShiftRowsOutput[81]), .S(MuxRound_n16), .Z(RoundOutput[81]) );
  MUX2_X1 MuxRound_mux_inst_82_U1 ( .A(ciphertext[18]), .B(ShiftRowsOutput[82]), .S(MuxRound_n16), .Z(RoundOutput[82]) );
  MUX2_X1 MuxRound_mux_inst_83_U1 ( .A(ciphertext[19]), .B(ShiftRowsOutput[83]), .S(MuxRound_n16), .Z(RoundOutput[83]) );
  MUX2_X1 MuxRound_mux_inst_84_U1 ( .A(ciphertext[20]), .B(ShiftRowsOutput[84]), .S(MuxRound_n16), .Z(RoundOutput[84]) );
  MUX2_X1 MuxRound_mux_inst_85_U1 ( .A(ciphertext[21]), .B(ShiftRowsOutput[85]), .S(MuxRound_n16), .Z(RoundOutput[85]) );
  MUX2_X1 MuxRound_mux_inst_86_U1 ( .A(ciphertext[22]), .B(ShiftRowsOutput[86]), .S(MuxRound_n16), .Z(RoundOutput[86]) );
  MUX2_X1 MuxRound_mux_inst_87_U1 ( .A(ciphertext[23]), .B(ShiftRowsOutput[87]), .S(MuxRound_n16), .Z(RoundOutput[87]) );
  MUX2_X1 MuxRound_mux_inst_88_U1 ( .A(ciphertext[56]), .B(ShiftRowsOutput[88]), .S(MuxRound_n16), .Z(RoundOutput[88]) );
  MUX2_X1 MuxRound_mux_inst_89_U1 ( .A(ciphertext[57]), .B(ShiftRowsOutput[89]), .S(MuxRound_n16), .Z(RoundOutput[89]) );
  MUX2_X1 MuxRound_mux_inst_90_U1 ( .A(ciphertext[58]), .B(ShiftRowsOutput[90]), .S(MuxRound_n16), .Z(RoundOutput[90]) );
  MUX2_X1 MuxRound_mux_inst_91_U1 ( .A(ciphertext[59]), .B(ShiftRowsOutput[91]), .S(MuxRound_n16), .Z(RoundOutput[91]) );
  MUX2_X1 MuxRound_mux_inst_92_U1 ( .A(ciphertext[60]), .B(ShiftRowsOutput[92]), .S(MuxRound_n15), .Z(RoundOutput[92]) );
  MUX2_X1 MuxRound_mux_inst_93_U1 ( .A(ciphertext[61]), .B(ShiftRowsOutput[93]), .S(MuxRound_n15), .Z(RoundOutput[93]) );
  MUX2_X1 MuxRound_mux_inst_94_U1 ( .A(ciphertext[62]), .B(ShiftRowsOutput[94]), .S(MuxRound_n15), .Z(RoundOutput[94]) );
  MUX2_X1 MuxRound_mux_inst_95_U1 ( .A(ciphertext[63]), .B(ShiftRowsOutput[95]), .S(MuxRound_n15), .Z(RoundOutput[95]) );
  MUX2_X1 MuxRound_mux_inst_96_U1 ( .A(ciphertext[96]), .B(ShiftRowsOutput[96]), .S(MuxRound_n15), .Z(RoundOutput[96]) );
  MUX2_X1 MuxRound_mux_inst_97_U1 ( .A(ciphertext[97]), .B(ShiftRowsOutput[97]), .S(MuxRound_n15), .Z(RoundOutput[97]) );
  MUX2_X1 MuxRound_mux_inst_98_U1 ( .A(ciphertext[98]), .B(ShiftRowsOutput[98]), .S(MuxRound_n15), .Z(RoundOutput[98]) );
  MUX2_X1 MuxRound_mux_inst_99_U1 ( .A(ciphertext[99]), .B(ShiftRowsOutput[99]), .S(MuxRound_n15), .Z(RoundOutput[99]) );
  MUX2_X1 MuxRound_mux_inst_100_U1 ( .A(ciphertext[100]), .B(
        ShiftRowsOutput[100]), .S(MuxRound_n15), .Z(RoundOutput[100]) );
  MUX2_X1 MuxRound_mux_inst_101_U1 ( .A(ciphertext[101]), .B(
        ShiftRowsOutput[101]), .S(MuxRound_n15), .Z(RoundOutput[101]) );
  MUX2_X1 MuxRound_mux_inst_102_U1 ( .A(ciphertext[102]), .B(
        ShiftRowsOutput[102]), .S(MuxRound_n15), .Z(RoundOutput[102]) );
  MUX2_X1 MuxRound_mux_inst_103_U1 ( .A(ciphertext[103]), .B(
        ShiftRowsOutput[103]), .S(MuxRound_n15), .Z(RoundOutput[103]) );
  MUX2_X1 MuxRound_mux_inst_104_U1 ( .A(ciphertext[8]), .B(
        ShiftRowsOutput[104]), .S(MuxRound_n14), .Z(RoundOutput[104]) );
  MUX2_X1 MuxRound_mux_inst_105_U1 ( .A(ciphertext[9]), .B(
        ShiftRowsOutput[105]), .S(MuxRound_n14), .Z(RoundOutput[105]) );
  MUX2_X1 MuxRound_mux_inst_106_U1 ( .A(ciphertext[10]), .B(
        ShiftRowsOutput[106]), .S(MuxRound_n14), .Z(RoundOutput[106]) );
  MUX2_X1 MuxRound_mux_inst_107_U1 ( .A(ciphertext[11]), .B(
        ShiftRowsOutput[107]), .S(MuxRound_n14), .Z(RoundOutput[107]) );
  MUX2_X1 MuxRound_mux_inst_108_U1 ( .A(ciphertext[12]), .B(
        ShiftRowsOutput[108]), .S(MuxRound_n14), .Z(RoundOutput[108]) );
  MUX2_X1 MuxRound_mux_inst_109_U1 ( .A(ciphertext[13]), .B(
        ShiftRowsOutput[109]), .S(MuxRound_n14), .Z(RoundOutput[109]) );
  MUX2_X1 MuxRound_mux_inst_110_U1 ( .A(ciphertext[14]), .B(
        ShiftRowsOutput[110]), .S(MuxRound_n14), .Z(RoundOutput[110]) );
  MUX2_X1 MuxRound_mux_inst_111_U1 ( .A(ciphertext[15]), .B(
        ShiftRowsOutput[111]), .S(MuxRound_n14), .Z(RoundOutput[111]) );
  MUX2_X1 MuxRound_mux_inst_112_U1 ( .A(ciphertext[48]), .B(
        ShiftRowsOutput[112]), .S(MuxRound_n14), .Z(RoundOutput[112]) );
  MUX2_X1 MuxRound_mux_inst_113_U1 ( .A(ciphertext[49]), .B(
        ShiftRowsOutput[113]), .S(MuxRound_n14), .Z(RoundOutput[113]) );
  MUX2_X1 MuxRound_mux_inst_114_U1 ( .A(ciphertext[50]), .B(
        ShiftRowsOutput[114]), .S(MuxRound_n14), .Z(RoundOutput[114]) );
  MUX2_X1 MuxRound_mux_inst_115_U1 ( .A(ciphertext[51]), .B(
        ShiftRowsOutput[115]), .S(MuxRound_n14), .Z(RoundOutput[115]) );
  MUX2_X1 MuxRound_mux_inst_116_U1 ( .A(ciphertext[52]), .B(
        ShiftRowsOutput[116]), .S(MuxRound_n13), .Z(RoundOutput[116]) );
  MUX2_X1 MuxRound_mux_inst_117_U1 ( .A(ciphertext[53]), .B(
        ShiftRowsOutput[117]), .S(MuxRound_n13), .Z(RoundOutput[117]) );
  MUX2_X1 MuxRound_mux_inst_118_U1 ( .A(ciphertext[54]), .B(
        ShiftRowsOutput[118]), .S(MuxRound_n13), .Z(RoundOutput[118]) );
  MUX2_X1 MuxRound_mux_inst_119_U1 ( .A(ciphertext[55]), .B(
        ShiftRowsOutput[119]), .S(MuxRound_n13), .Z(RoundOutput[119]) );
  MUX2_X1 MuxRound_mux_inst_120_U1 ( .A(ciphertext[88]), .B(
        ShiftRowsOutput[120]), .S(MuxRound_n13), .Z(RoundOutput[120]) );
  MUX2_X1 MuxRound_mux_inst_121_U1 ( .A(ciphertext[89]), .B(
        ShiftRowsOutput[121]), .S(MuxRound_n13), .Z(RoundOutput[121]) );
  MUX2_X1 MuxRound_mux_inst_122_U1 ( .A(ciphertext[90]), .B(
        ShiftRowsOutput[122]), .S(MuxRound_n13), .Z(RoundOutput[122]) );
  MUX2_X1 MuxRound_mux_inst_123_U1 ( .A(ciphertext[91]), .B(
        ShiftRowsOutput[123]), .S(MuxRound_n13), .Z(RoundOutput[123]) );
  MUX2_X1 MuxRound_mux_inst_124_U1 ( .A(ciphertext[92]), .B(
        ShiftRowsOutput[124]), .S(MuxRound_n13), .Z(RoundOutput[124]) );
  MUX2_X1 MuxRound_mux_inst_125_U1 ( .A(ciphertext[93]), .B(
        ShiftRowsOutput[125]), .S(MuxRound_n13), .Z(RoundOutput[125]) );
  MUX2_X1 MuxRound_mux_inst_126_U1 ( .A(ciphertext[94]), .B(
        ShiftRowsOutput[126]), .S(MuxRound_n13), .Z(RoundOutput[126]) );
  MUX2_X1 MuxRound_mux_inst_127_U1 ( .A(ciphertext[95]), .B(
        ShiftRowsOutput[127]), .S(MuxRound_n13), .Z(RoundOutput[127]) );
  INV_X1 KeyReg_Inst_ff_SDE_0_current_state_reg_U1 ( .A(KSSubBytesInput[16]), 
        .ZN(KeyReg_Inst_ff_SDE_0_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_0_next_state), .CK(clk), .Q(KSSubBytesInput[16]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_0_MUX_inst_U1 ( .A(RoundKeyOutput[0]), .B(key[0]), 
        .S(reset), .Z(KeyReg_Inst_ff_SDE_0_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_1_current_state_reg_U1 ( .A(KSSubBytesInput[17]), 
        .ZN(KeyReg_Inst_ff_SDE_1_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_1_next_state), .CK(clk), .Q(KSSubBytesInput[17]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_1_MUX_inst_U1 ( .A(RoundKeyOutput[1]), .B(key[1]), 
        .S(reset), .Z(KeyReg_Inst_ff_SDE_1_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_2_current_state_reg_U1 ( .A(KSSubBytesInput[18]), 
        .ZN(KeyReg_Inst_ff_SDE_2_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_2_next_state), .CK(clk), .Q(KSSubBytesInput[18]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_2_MUX_inst_U1 ( .A(RoundKeyOutput[2]), .B(key[2]), 
        .S(reset), .Z(KeyReg_Inst_ff_SDE_2_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_3_current_state_reg_U1 ( .A(KSSubBytesInput[19]), 
        .ZN(KeyReg_Inst_ff_SDE_3_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_3_next_state), .CK(clk), .Q(KSSubBytesInput[19]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_3_MUX_inst_U1 ( .A(RoundKeyOutput[3]), .B(key[3]), 
        .S(reset), .Z(KeyReg_Inst_ff_SDE_3_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_4_current_state_reg_U1 ( .A(KSSubBytesInput[20]), 
        .ZN(KeyReg_Inst_ff_SDE_4_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_4_next_state), .CK(clk), .Q(KSSubBytesInput[20]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_4_MUX_inst_U1 ( .A(RoundKeyOutput[4]), .B(key[4]), 
        .S(reset), .Z(KeyReg_Inst_ff_SDE_4_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_5_current_state_reg_U1 ( .A(KSSubBytesInput[21]), 
        .ZN(KeyReg_Inst_ff_SDE_5_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_5_next_state), .CK(clk), .Q(KSSubBytesInput[21]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_5_MUX_inst_U1 ( .A(RoundKeyOutput[5]), .B(key[5]), 
        .S(reset), .Z(KeyReg_Inst_ff_SDE_5_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_6_current_state_reg_U1 ( .A(KSSubBytesInput[22]), 
        .ZN(KeyReg_Inst_ff_SDE_6_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_6_next_state), .CK(clk), .Q(KSSubBytesInput[22]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_6_MUX_inst_U1 ( .A(RoundKeyOutput[6]), .B(key[6]), 
        .S(reset), .Z(KeyReg_Inst_ff_SDE_6_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_7_current_state_reg_U1 ( .A(KSSubBytesInput[23]), 
        .ZN(KeyReg_Inst_ff_SDE_7_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_7_next_state), .CK(clk), .Q(KSSubBytesInput[23]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_7_MUX_inst_U1 ( .A(RoundKeyOutput[7]), .B(key[7]), 
        .S(reset), .Z(KeyReg_Inst_ff_SDE_7_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_8_current_state_reg_U1 ( .A(KSSubBytesInput[8]), 
        .ZN(KeyReg_Inst_ff_SDE_8_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_8_next_state), .CK(clk), .Q(KSSubBytesInput[8]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_8_MUX_inst_U1 ( .A(RoundKeyOutput[8]), .B(key[8]), 
        .S(reset), .Z(KeyReg_Inst_ff_SDE_8_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_9_current_state_reg_U1 ( .A(KSSubBytesInput[9]), 
        .ZN(KeyReg_Inst_ff_SDE_9_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_9_next_state), .CK(clk), .Q(KSSubBytesInput[9]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_9_MUX_inst_U1 ( .A(RoundKeyOutput[9]), .B(key[9]), 
        .S(reset), .Z(KeyReg_Inst_ff_SDE_9_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_10_current_state_reg_U1 ( .A(KSSubBytesInput[10]), 
        .ZN(KeyReg_Inst_ff_SDE_10_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_10_next_state), .CK(clk), .Q(KSSubBytesInput[10]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_10_MUX_inst_U1 ( .A(RoundKeyOutput[10]), .B(
        key[10]), .S(reset), .Z(KeyReg_Inst_ff_SDE_10_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_11_current_state_reg_U1 ( .A(KSSubBytesInput[11]), 
        .ZN(KeyReg_Inst_ff_SDE_11_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_11_next_state), .CK(clk), .Q(KSSubBytesInput[11]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_11_MUX_inst_U1 ( .A(RoundKeyOutput[11]), .B(
        key[11]), .S(reset), .Z(KeyReg_Inst_ff_SDE_11_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_12_current_state_reg_U1 ( .A(KSSubBytesInput[12]), 
        .ZN(KeyReg_Inst_ff_SDE_12_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_12_next_state), .CK(clk), .Q(KSSubBytesInput[12]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_12_MUX_inst_U1 ( .A(RoundKeyOutput[12]), .B(
        key[12]), .S(reset), .Z(KeyReg_Inst_ff_SDE_12_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_13_current_state_reg_U1 ( .A(KSSubBytesInput[13]), 
        .ZN(KeyReg_Inst_ff_SDE_13_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_13_next_state), .CK(clk), .Q(KSSubBytesInput[13]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_13_MUX_inst_U1 ( .A(RoundKeyOutput[13]), .B(
        key[13]), .S(reset), .Z(KeyReg_Inst_ff_SDE_13_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_14_current_state_reg_U1 ( .A(KSSubBytesInput[14]), 
        .ZN(KeyReg_Inst_ff_SDE_14_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_14_next_state), .CK(clk), .Q(KSSubBytesInput[14]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_14_MUX_inst_U1 ( .A(RoundKeyOutput[14]), .B(
        key[14]), .S(reset), .Z(KeyReg_Inst_ff_SDE_14_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_15_current_state_reg_U1 ( .A(KSSubBytesInput[15]), 
        .ZN(KeyReg_Inst_ff_SDE_15_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_15_next_state), .CK(clk), .Q(KSSubBytesInput[15]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_15_MUX_inst_U1 ( .A(RoundKeyOutput[15]), .B(
        key[15]), .S(reset), .Z(KeyReg_Inst_ff_SDE_15_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_16_current_state_reg_U1 ( .A(KSSubBytesInput[0]), 
        .ZN(KeyReg_Inst_ff_SDE_16_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_16_next_state), .CK(clk), .Q(KSSubBytesInput[0]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_16_MUX_inst_U1 ( .A(RoundKeyOutput[16]), .B(
        key[16]), .S(reset), .Z(KeyReg_Inst_ff_SDE_16_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_17_current_state_reg_U1 ( .A(KSSubBytesInput[1]), 
        .ZN(KeyReg_Inst_ff_SDE_17_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_17_next_state), .CK(clk), .Q(KSSubBytesInput[1]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_17_MUX_inst_U1 ( .A(RoundKeyOutput[17]), .B(
        key[17]), .S(reset), .Z(KeyReg_Inst_ff_SDE_17_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_18_current_state_reg_U1 ( .A(KSSubBytesInput[2]), 
        .ZN(KeyReg_Inst_ff_SDE_18_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_18_next_state), .CK(clk), .Q(KSSubBytesInput[2]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_18_MUX_inst_U1 ( .A(RoundKeyOutput[18]), .B(
        key[18]), .S(reset), .Z(KeyReg_Inst_ff_SDE_18_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_19_current_state_reg_U1 ( .A(KSSubBytesInput[3]), 
        .ZN(KeyReg_Inst_ff_SDE_19_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_19_next_state), .CK(clk), .Q(KSSubBytesInput[3]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_19_MUX_inst_U1 ( .A(RoundKeyOutput[19]), .B(
        key[19]), .S(reset), .Z(KeyReg_Inst_ff_SDE_19_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_20_current_state_reg_U1 ( .A(KSSubBytesInput[4]), 
        .ZN(KeyReg_Inst_ff_SDE_20_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_20_next_state), .CK(clk), .Q(KSSubBytesInput[4]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_20_MUX_inst_U1 ( .A(RoundKeyOutput[20]), .B(
        key[20]), .S(reset), .Z(KeyReg_Inst_ff_SDE_20_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_21_current_state_reg_U1 ( .A(KSSubBytesInput[5]), 
        .ZN(KeyReg_Inst_ff_SDE_21_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_21_next_state), .CK(clk), .Q(KSSubBytesInput[5]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_21_MUX_inst_U1 ( .A(RoundKeyOutput[21]), .B(
        key[21]), .S(reset), .Z(KeyReg_Inst_ff_SDE_21_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_22_current_state_reg_U1 ( .A(KSSubBytesInput[6]), 
        .ZN(KeyReg_Inst_ff_SDE_22_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_22_next_state), .CK(clk), .Q(KSSubBytesInput[6]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_22_MUX_inst_U1 ( .A(RoundKeyOutput[22]), .B(
        key[22]), .S(reset), .Z(KeyReg_Inst_ff_SDE_22_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_23_current_state_reg_U1 ( .A(KSSubBytesInput[7]), 
        .ZN(KeyReg_Inst_ff_SDE_23_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_23_next_state), .CK(clk), .Q(KSSubBytesInput[7]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_23_MUX_inst_U1 ( .A(RoundKeyOutput[23]), .B(
        key[23]), .S(reset), .Z(KeyReg_Inst_ff_SDE_23_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_24_current_state_reg_U1 ( .A(KSSubBytesInput[24]), 
        .ZN(KeyReg_Inst_ff_SDE_24_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_24_next_state), .CK(clk), .Q(KSSubBytesInput[24]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_24_MUX_inst_U1 ( .A(RoundKeyOutput[24]), .B(
        key[24]), .S(reset), .Z(KeyReg_Inst_ff_SDE_24_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_25_current_state_reg_U1 ( .A(KSSubBytesInput[25]), 
        .ZN(KeyReg_Inst_ff_SDE_25_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_25_next_state), .CK(clk), .Q(KSSubBytesInput[25]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_25_MUX_inst_U1 ( .A(RoundKeyOutput[25]), .B(
        key[25]), .S(reset), .Z(KeyReg_Inst_ff_SDE_25_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_26_current_state_reg_U1 ( .A(KSSubBytesInput[26]), 
        .ZN(KeyReg_Inst_ff_SDE_26_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_26_next_state), .CK(clk), .Q(KSSubBytesInput[26]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_26_MUX_inst_U1 ( .A(RoundKeyOutput[26]), .B(
        key[26]), .S(reset), .Z(KeyReg_Inst_ff_SDE_26_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_27_current_state_reg_U1 ( .A(KSSubBytesInput[27]), 
        .ZN(KeyReg_Inst_ff_SDE_27_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_27_next_state), .CK(clk), .Q(KSSubBytesInput[27]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_27_MUX_inst_U1 ( .A(RoundKeyOutput[27]), .B(
        key[27]), .S(reset), .Z(KeyReg_Inst_ff_SDE_27_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_28_current_state_reg_U1 ( .A(KSSubBytesInput[28]), 
        .ZN(KeyReg_Inst_ff_SDE_28_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_28_next_state), .CK(clk), .Q(KSSubBytesInput[28]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_28_MUX_inst_U1 ( .A(RoundKeyOutput[28]), .B(
        key[28]), .S(reset), .Z(KeyReg_Inst_ff_SDE_28_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_29_current_state_reg_U1 ( .A(KSSubBytesInput[29]), 
        .ZN(KeyReg_Inst_ff_SDE_29_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_29_next_state), .CK(clk), .Q(KSSubBytesInput[29]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_29_MUX_inst_U1 ( .A(RoundKeyOutput[29]), .B(
        key[29]), .S(reset), .Z(KeyReg_Inst_ff_SDE_29_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_30_current_state_reg_U1 ( .A(KSSubBytesInput[30]), 
        .ZN(KeyReg_Inst_ff_SDE_30_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_30_next_state), .CK(clk), .Q(KSSubBytesInput[30]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_30_MUX_inst_U1 ( .A(RoundKeyOutput[30]), .B(
        key[30]), .S(reset), .Z(KeyReg_Inst_ff_SDE_30_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_31_current_state_reg_U1 ( .A(KSSubBytesInput[31]), 
        .ZN(KeyReg_Inst_ff_SDE_31_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_31_next_state), .CK(clk), .Q(KSSubBytesInput[31]), 
        .QN() );
  MUX2_X1 KeyReg_Inst_ff_SDE_31_MUX_inst_U1 ( .A(RoundKeyOutput[31]), .B(
        key[31]), .S(reset), .Z(KeyReg_Inst_ff_SDE_31_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_32_current_state_reg_U1 ( .A(RoundKey[32]), .ZN(
        KeyReg_Inst_ff_SDE_32_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_32_next_state), .CK(clk), .Q(RoundKey[32]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_32_MUX_inst_U1 ( .A(RoundKeyOutput[32]), .B(
        key[32]), .S(reset), .Z(KeyReg_Inst_ff_SDE_32_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_33_current_state_reg_U1 ( .A(RoundKey[33]), .ZN(
        KeyReg_Inst_ff_SDE_33_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_33_next_state), .CK(clk), .Q(RoundKey[33]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_33_MUX_inst_U1 ( .A(RoundKeyOutput[33]), .B(
        key[33]), .S(reset), .Z(KeyReg_Inst_ff_SDE_33_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_34_current_state_reg_U1 ( .A(RoundKey[34]), .ZN(
        KeyReg_Inst_ff_SDE_34_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_34_next_state), .CK(clk), .Q(RoundKey[34]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_34_MUX_inst_U1 ( .A(RoundKeyOutput[34]), .B(
        key[34]), .S(reset), .Z(KeyReg_Inst_ff_SDE_34_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_35_current_state_reg_U1 ( .A(RoundKey[35]), .ZN(
        KeyReg_Inst_ff_SDE_35_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_35_next_state), .CK(clk), .Q(RoundKey[35]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_35_MUX_inst_U1 ( .A(RoundKeyOutput[35]), .B(
        key[35]), .S(reset), .Z(KeyReg_Inst_ff_SDE_35_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_36_current_state_reg_U1 ( .A(RoundKey[36]), .ZN(
        KeyReg_Inst_ff_SDE_36_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_36_next_state), .CK(clk), .Q(RoundKey[36]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_36_MUX_inst_U1 ( .A(RoundKeyOutput[36]), .B(
        key[36]), .S(reset), .Z(KeyReg_Inst_ff_SDE_36_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_37_current_state_reg_U1 ( .A(RoundKey[37]), .ZN(
        KeyReg_Inst_ff_SDE_37_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_37_next_state), .CK(clk), .Q(RoundKey[37]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_37_MUX_inst_U1 ( .A(RoundKeyOutput[37]), .B(
        key[37]), .S(reset), .Z(KeyReg_Inst_ff_SDE_37_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_38_current_state_reg_U1 ( .A(RoundKey[38]), .ZN(
        KeyReg_Inst_ff_SDE_38_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_38_next_state), .CK(clk), .Q(RoundKey[38]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_38_MUX_inst_U1 ( .A(RoundKeyOutput[38]), .B(
        key[38]), .S(reset), .Z(KeyReg_Inst_ff_SDE_38_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_39_current_state_reg_U1 ( .A(RoundKey[39]), .ZN(
        KeyReg_Inst_ff_SDE_39_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_39_next_state), .CK(clk), .Q(RoundKey[39]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_39_MUX_inst_U1 ( .A(RoundKeyOutput[39]), .B(
        key[39]), .S(reset), .Z(KeyReg_Inst_ff_SDE_39_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_40_current_state_reg_U1 ( .A(RoundKey[40]), .ZN(
        KeyReg_Inst_ff_SDE_40_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_40_next_state), .CK(clk), .Q(RoundKey[40]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_40_MUX_inst_U1 ( .A(RoundKeyOutput[40]), .B(
        key[40]), .S(reset), .Z(KeyReg_Inst_ff_SDE_40_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_41_current_state_reg_U1 ( .A(RoundKey[41]), .ZN(
        KeyReg_Inst_ff_SDE_41_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_41_next_state), .CK(clk), .Q(RoundKey[41]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_41_MUX_inst_U1 ( .A(RoundKeyOutput[41]), .B(
        key[41]), .S(reset), .Z(KeyReg_Inst_ff_SDE_41_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_42_current_state_reg_U1 ( .A(RoundKey[42]), .ZN(
        KeyReg_Inst_ff_SDE_42_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_42_next_state), .CK(clk), .Q(RoundKey[42]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_42_MUX_inst_U1 ( .A(RoundKeyOutput[42]), .B(
        key[42]), .S(reset), .Z(KeyReg_Inst_ff_SDE_42_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_43_current_state_reg_U1 ( .A(RoundKey[43]), .ZN(
        KeyReg_Inst_ff_SDE_43_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_43_next_state), .CK(clk), .Q(RoundKey[43]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_43_MUX_inst_U1 ( .A(RoundKeyOutput[43]), .B(
        key[43]), .S(reset), .Z(KeyReg_Inst_ff_SDE_43_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_44_current_state_reg_U1 ( .A(RoundKey[44]), .ZN(
        KeyReg_Inst_ff_SDE_44_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_44_next_state), .CK(clk), .Q(RoundKey[44]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_44_MUX_inst_U1 ( .A(RoundKeyOutput[44]), .B(
        key[44]), .S(reset), .Z(KeyReg_Inst_ff_SDE_44_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_45_current_state_reg_U1 ( .A(RoundKey[45]), .ZN(
        KeyReg_Inst_ff_SDE_45_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_45_next_state), .CK(clk), .Q(RoundKey[45]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_45_MUX_inst_U1 ( .A(RoundKeyOutput[45]), .B(
        key[45]), .S(reset), .Z(KeyReg_Inst_ff_SDE_45_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_46_current_state_reg_U1 ( .A(RoundKey[46]), .ZN(
        KeyReg_Inst_ff_SDE_46_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_46_next_state), .CK(clk), .Q(RoundKey[46]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_46_MUX_inst_U1 ( .A(RoundKeyOutput[46]), .B(
        key[46]), .S(reset), .Z(KeyReg_Inst_ff_SDE_46_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_47_current_state_reg_U1 ( .A(RoundKey[47]), .ZN(
        KeyReg_Inst_ff_SDE_47_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_47_next_state), .CK(clk), .Q(RoundKey[47]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_47_MUX_inst_U1 ( .A(RoundKeyOutput[47]), .B(
        key[47]), .S(reset), .Z(KeyReg_Inst_ff_SDE_47_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_48_current_state_reg_U1 ( .A(RoundKey[48]), .ZN(
        KeyReg_Inst_ff_SDE_48_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_48_next_state), .CK(clk), .Q(RoundKey[48]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_48_MUX_inst_U1 ( .A(RoundKeyOutput[48]), .B(
        key[48]), .S(reset), .Z(KeyReg_Inst_ff_SDE_48_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_49_current_state_reg_U1 ( .A(RoundKey[49]), .ZN(
        KeyReg_Inst_ff_SDE_49_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_49_next_state), .CK(clk), .Q(RoundKey[49]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_49_MUX_inst_U1 ( .A(RoundKeyOutput[49]), .B(
        key[49]), .S(reset), .Z(KeyReg_Inst_ff_SDE_49_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_50_current_state_reg_U1 ( .A(RoundKey[50]), .ZN(
        KeyReg_Inst_ff_SDE_50_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_50_next_state), .CK(clk), .Q(RoundKey[50]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_50_MUX_inst_U1 ( .A(RoundKeyOutput[50]), .B(
        key[50]), .S(reset), .Z(KeyReg_Inst_ff_SDE_50_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_51_current_state_reg_U1 ( .A(RoundKey[51]), .ZN(
        KeyReg_Inst_ff_SDE_51_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_51_next_state), .CK(clk), .Q(RoundKey[51]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_51_MUX_inst_U1 ( .A(RoundKeyOutput[51]), .B(
        key[51]), .S(reset), .Z(KeyReg_Inst_ff_SDE_51_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_52_current_state_reg_U1 ( .A(RoundKey[52]), .ZN(
        KeyReg_Inst_ff_SDE_52_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_52_next_state), .CK(clk), .Q(RoundKey[52]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_52_MUX_inst_U1 ( .A(RoundKeyOutput[52]), .B(
        key[52]), .S(reset), .Z(KeyReg_Inst_ff_SDE_52_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_53_current_state_reg_U1 ( .A(RoundKey[53]), .ZN(
        KeyReg_Inst_ff_SDE_53_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_53_next_state), .CK(clk), .Q(RoundKey[53]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_53_MUX_inst_U1 ( .A(RoundKeyOutput[53]), .B(
        key[53]), .S(reset), .Z(KeyReg_Inst_ff_SDE_53_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_54_current_state_reg_U1 ( .A(RoundKey[54]), .ZN(
        KeyReg_Inst_ff_SDE_54_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_54_next_state), .CK(clk), .Q(RoundKey[54]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_54_MUX_inst_U1 ( .A(RoundKeyOutput[54]), .B(
        key[54]), .S(reset), .Z(KeyReg_Inst_ff_SDE_54_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_55_current_state_reg_U1 ( .A(RoundKey[55]), .ZN(
        KeyReg_Inst_ff_SDE_55_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_55_next_state), .CK(clk), .Q(RoundKey[55]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_55_MUX_inst_U1 ( .A(RoundKeyOutput[55]), .B(
        key[55]), .S(reset), .Z(KeyReg_Inst_ff_SDE_55_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_56_current_state_reg_U1 ( .A(RoundKey[56]), .ZN(
        KeyReg_Inst_ff_SDE_56_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_56_next_state), .CK(clk), .Q(RoundKey[56]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_56_MUX_inst_U1 ( .A(RoundKeyOutput[56]), .B(
        key[56]), .S(reset), .Z(KeyReg_Inst_ff_SDE_56_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_57_current_state_reg_U1 ( .A(RoundKey[57]), .ZN(
        KeyReg_Inst_ff_SDE_57_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_57_next_state), .CK(clk), .Q(RoundKey[57]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_57_MUX_inst_U1 ( .A(RoundKeyOutput[57]), .B(
        key[57]), .S(reset), .Z(KeyReg_Inst_ff_SDE_57_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_58_current_state_reg_U1 ( .A(RoundKey[58]), .ZN(
        KeyReg_Inst_ff_SDE_58_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_58_next_state), .CK(clk), .Q(RoundKey[58]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_58_MUX_inst_U1 ( .A(RoundKeyOutput[58]), .B(
        key[58]), .S(reset), .Z(KeyReg_Inst_ff_SDE_58_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_59_current_state_reg_U1 ( .A(RoundKey[59]), .ZN(
        KeyReg_Inst_ff_SDE_59_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_59_next_state), .CK(clk), .Q(RoundKey[59]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_59_MUX_inst_U1 ( .A(RoundKeyOutput[59]), .B(
        key[59]), .S(reset), .Z(KeyReg_Inst_ff_SDE_59_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_60_current_state_reg_U1 ( .A(RoundKey[60]), .ZN(
        KeyReg_Inst_ff_SDE_60_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_60_next_state), .CK(clk), .Q(RoundKey[60]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_60_MUX_inst_U1 ( .A(RoundKeyOutput[60]), .B(
        key[60]), .S(reset), .Z(KeyReg_Inst_ff_SDE_60_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_61_current_state_reg_U1 ( .A(RoundKey[61]), .ZN(
        KeyReg_Inst_ff_SDE_61_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_61_next_state), .CK(clk), .Q(RoundKey[61]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_61_MUX_inst_U1 ( .A(RoundKeyOutput[61]), .B(
        key[61]), .S(reset), .Z(KeyReg_Inst_ff_SDE_61_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_62_current_state_reg_U1 ( .A(RoundKey[62]), .ZN(
        KeyReg_Inst_ff_SDE_62_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_62_next_state), .CK(clk), .Q(RoundKey[62]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_62_MUX_inst_U1 ( .A(RoundKeyOutput[62]), .B(
        key[62]), .S(reset), .Z(KeyReg_Inst_ff_SDE_62_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_63_current_state_reg_U1 ( .A(RoundKey[63]), .ZN(
        KeyReg_Inst_ff_SDE_63_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_63_next_state), .CK(clk), .Q(RoundKey[63]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_63_MUX_inst_U1 ( .A(RoundKeyOutput[63]), .B(
        key[63]), .S(reset), .Z(KeyReg_Inst_ff_SDE_63_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_64_current_state_reg_U1 ( .A(RoundKey[64]), .ZN(
        KeyReg_Inst_ff_SDE_64_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_64_next_state), .CK(clk), .Q(RoundKey[64]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_64_MUX_inst_U1 ( .A(RoundKeyOutput[64]), .B(
        key[64]), .S(reset), .Z(KeyReg_Inst_ff_SDE_64_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_65_current_state_reg_U1 ( .A(RoundKey[65]), .ZN(
        KeyReg_Inst_ff_SDE_65_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_65_next_state), .CK(clk), .Q(RoundKey[65]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_65_MUX_inst_U1 ( .A(RoundKeyOutput[65]), .B(
        key[65]), .S(reset), .Z(KeyReg_Inst_ff_SDE_65_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_66_current_state_reg_U1 ( .A(RoundKey[66]), .ZN(
        KeyReg_Inst_ff_SDE_66_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_66_next_state), .CK(clk), .Q(RoundKey[66]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_66_MUX_inst_U1 ( .A(RoundKeyOutput[66]), .B(
        key[66]), .S(reset), .Z(KeyReg_Inst_ff_SDE_66_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_67_current_state_reg_U1 ( .A(RoundKey[67]), .ZN(
        KeyReg_Inst_ff_SDE_67_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_67_next_state), .CK(clk), .Q(RoundKey[67]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_67_MUX_inst_U1 ( .A(RoundKeyOutput[67]), .B(
        key[67]), .S(reset), .Z(KeyReg_Inst_ff_SDE_67_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_68_current_state_reg_U1 ( .A(RoundKey[68]), .ZN(
        KeyReg_Inst_ff_SDE_68_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_68_next_state), .CK(clk), .Q(RoundKey[68]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_68_MUX_inst_U1 ( .A(RoundKeyOutput[68]), .B(
        key[68]), .S(reset), .Z(KeyReg_Inst_ff_SDE_68_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_69_current_state_reg_U1 ( .A(RoundKey[69]), .ZN(
        KeyReg_Inst_ff_SDE_69_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_69_next_state), .CK(clk), .Q(RoundKey[69]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_69_MUX_inst_U1 ( .A(RoundKeyOutput[69]), .B(
        key[69]), .S(reset), .Z(KeyReg_Inst_ff_SDE_69_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_70_current_state_reg_U1 ( .A(RoundKey[70]), .ZN(
        KeyReg_Inst_ff_SDE_70_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_70_next_state), .CK(clk), .Q(RoundKey[70]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_70_MUX_inst_U1 ( .A(RoundKeyOutput[70]), .B(
        key[70]), .S(reset), .Z(KeyReg_Inst_ff_SDE_70_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_71_current_state_reg_U1 ( .A(RoundKey[71]), .ZN(
        KeyReg_Inst_ff_SDE_71_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_71_next_state), .CK(clk), .Q(RoundKey[71]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_71_MUX_inst_U1 ( .A(RoundKeyOutput[71]), .B(
        key[71]), .S(reset), .Z(KeyReg_Inst_ff_SDE_71_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_72_current_state_reg_U1 ( .A(RoundKey[72]), .ZN(
        KeyReg_Inst_ff_SDE_72_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_72_next_state), .CK(clk), .Q(RoundKey[72]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_72_MUX_inst_U1 ( .A(RoundKeyOutput[72]), .B(
        key[72]), .S(reset), .Z(KeyReg_Inst_ff_SDE_72_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_73_current_state_reg_U1 ( .A(RoundKey[73]), .ZN(
        KeyReg_Inst_ff_SDE_73_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_73_next_state), .CK(clk), .Q(RoundKey[73]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_73_MUX_inst_U1 ( .A(RoundKeyOutput[73]), .B(
        key[73]), .S(reset), .Z(KeyReg_Inst_ff_SDE_73_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_74_current_state_reg_U1 ( .A(RoundKey[74]), .ZN(
        KeyReg_Inst_ff_SDE_74_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_74_next_state), .CK(clk), .Q(RoundKey[74]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_74_MUX_inst_U1 ( .A(RoundKeyOutput[74]), .B(
        key[74]), .S(reset), .Z(KeyReg_Inst_ff_SDE_74_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_75_current_state_reg_U1 ( .A(RoundKey[75]), .ZN(
        KeyReg_Inst_ff_SDE_75_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_75_next_state), .CK(clk), .Q(RoundKey[75]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_75_MUX_inst_U1 ( .A(RoundKeyOutput[75]), .B(
        key[75]), .S(reset), .Z(KeyReg_Inst_ff_SDE_75_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_76_current_state_reg_U1 ( .A(RoundKey[76]), .ZN(
        KeyReg_Inst_ff_SDE_76_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_76_next_state), .CK(clk), .Q(RoundKey[76]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_76_MUX_inst_U1 ( .A(RoundKeyOutput[76]), .B(
        key[76]), .S(reset), .Z(KeyReg_Inst_ff_SDE_76_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_77_current_state_reg_U1 ( .A(RoundKey[77]), .ZN(
        KeyReg_Inst_ff_SDE_77_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_77_next_state), .CK(clk), .Q(RoundKey[77]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_77_MUX_inst_U1 ( .A(RoundKeyOutput[77]), .B(
        key[77]), .S(reset), .Z(KeyReg_Inst_ff_SDE_77_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_78_current_state_reg_U1 ( .A(RoundKey[78]), .ZN(
        KeyReg_Inst_ff_SDE_78_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_78_next_state), .CK(clk), .Q(RoundKey[78]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_78_MUX_inst_U1 ( .A(RoundKeyOutput[78]), .B(
        key[78]), .S(reset), .Z(KeyReg_Inst_ff_SDE_78_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_79_current_state_reg_U1 ( .A(RoundKey[79]), .ZN(
        KeyReg_Inst_ff_SDE_79_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_79_next_state), .CK(clk), .Q(RoundKey[79]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_79_MUX_inst_U1 ( .A(RoundKeyOutput[79]), .B(
        key[79]), .S(reset), .Z(KeyReg_Inst_ff_SDE_79_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_80_current_state_reg_U1 ( .A(RoundKey[80]), .ZN(
        KeyReg_Inst_ff_SDE_80_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_80_next_state), .CK(clk), .Q(RoundKey[80]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_80_MUX_inst_U1 ( .A(RoundKeyOutput[80]), .B(
        key[80]), .S(reset), .Z(KeyReg_Inst_ff_SDE_80_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_81_current_state_reg_U1 ( .A(RoundKey[81]), .ZN(
        KeyReg_Inst_ff_SDE_81_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_81_next_state), .CK(clk), .Q(RoundKey[81]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_81_MUX_inst_U1 ( .A(RoundKeyOutput[81]), .B(
        key[81]), .S(reset), .Z(KeyReg_Inst_ff_SDE_81_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_82_current_state_reg_U1 ( .A(RoundKey[82]), .ZN(
        KeyReg_Inst_ff_SDE_82_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_82_next_state), .CK(clk), .Q(RoundKey[82]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_82_MUX_inst_U1 ( .A(RoundKeyOutput[82]), .B(
        key[82]), .S(reset), .Z(KeyReg_Inst_ff_SDE_82_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_83_current_state_reg_U1 ( .A(RoundKey[83]), .ZN(
        KeyReg_Inst_ff_SDE_83_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_83_next_state), .CK(clk), .Q(RoundKey[83]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_83_MUX_inst_U1 ( .A(RoundKeyOutput[83]), .B(
        key[83]), .S(reset), .Z(KeyReg_Inst_ff_SDE_83_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_84_current_state_reg_U1 ( .A(RoundKey[84]), .ZN(
        KeyReg_Inst_ff_SDE_84_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_84_next_state), .CK(clk), .Q(RoundKey[84]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_84_MUX_inst_U1 ( .A(RoundKeyOutput[84]), .B(
        key[84]), .S(reset), .Z(KeyReg_Inst_ff_SDE_84_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_85_current_state_reg_U1 ( .A(RoundKey[85]), .ZN(
        KeyReg_Inst_ff_SDE_85_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_85_next_state), .CK(clk), .Q(RoundKey[85]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_85_MUX_inst_U1 ( .A(RoundKeyOutput[85]), .B(
        key[85]), .S(reset), .Z(KeyReg_Inst_ff_SDE_85_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_86_current_state_reg_U1 ( .A(RoundKey[86]), .ZN(
        KeyReg_Inst_ff_SDE_86_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_86_next_state), .CK(clk), .Q(RoundKey[86]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_86_MUX_inst_U1 ( .A(RoundKeyOutput[86]), .B(
        key[86]), .S(reset), .Z(KeyReg_Inst_ff_SDE_86_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_87_current_state_reg_U1 ( .A(RoundKey[87]), .ZN(
        KeyReg_Inst_ff_SDE_87_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_87_next_state), .CK(clk), .Q(RoundKey[87]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_87_MUX_inst_U1 ( .A(RoundKeyOutput[87]), .B(
        key[87]), .S(reset), .Z(KeyReg_Inst_ff_SDE_87_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_88_current_state_reg_U1 ( .A(RoundKey[88]), .ZN(
        KeyReg_Inst_ff_SDE_88_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_88_next_state), .CK(clk), .Q(RoundKey[88]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_88_MUX_inst_U1 ( .A(RoundKeyOutput[88]), .B(
        key[88]), .S(reset), .Z(KeyReg_Inst_ff_SDE_88_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_89_current_state_reg_U1 ( .A(RoundKey[89]), .ZN(
        KeyReg_Inst_ff_SDE_89_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_89_next_state), .CK(clk), .Q(RoundKey[89]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_89_MUX_inst_U1 ( .A(RoundKeyOutput[89]), .B(
        key[89]), .S(reset), .Z(KeyReg_Inst_ff_SDE_89_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_90_current_state_reg_U1 ( .A(RoundKey[90]), .ZN(
        KeyReg_Inst_ff_SDE_90_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_90_next_state), .CK(clk), .Q(RoundKey[90]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_90_MUX_inst_U1 ( .A(RoundKeyOutput[90]), .B(
        key[90]), .S(reset), .Z(KeyReg_Inst_ff_SDE_90_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_91_current_state_reg_U1 ( .A(RoundKey[91]), .ZN(
        KeyReg_Inst_ff_SDE_91_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_91_next_state), .CK(clk), .Q(RoundKey[91]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_91_MUX_inst_U1 ( .A(RoundKeyOutput[91]), .B(
        key[91]), .S(reset), .Z(KeyReg_Inst_ff_SDE_91_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_92_current_state_reg_U1 ( .A(RoundKey[92]), .ZN(
        KeyReg_Inst_ff_SDE_92_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_92_next_state), .CK(clk), .Q(RoundKey[92]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_92_MUX_inst_U1 ( .A(RoundKeyOutput[92]), .B(
        key[92]), .S(reset), .Z(KeyReg_Inst_ff_SDE_92_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_93_current_state_reg_U1 ( .A(RoundKey[93]), .ZN(
        KeyReg_Inst_ff_SDE_93_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_93_next_state), .CK(clk), .Q(RoundKey[93]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_93_MUX_inst_U1 ( .A(RoundKeyOutput[93]), .B(
        key[93]), .S(reset), .Z(KeyReg_Inst_ff_SDE_93_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_94_current_state_reg_U1 ( .A(RoundKey[94]), .ZN(
        KeyReg_Inst_ff_SDE_94_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_94_next_state), .CK(clk), .Q(RoundKey[94]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_94_MUX_inst_U1 ( .A(RoundKeyOutput[94]), .B(
        key[94]), .S(reset), .Z(KeyReg_Inst_ff_SDE_94_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_95_current_state_reg_U1 ( .A(RoundKey[95]), .ZN(
        KeyReg_Inst_ff_SDE_95_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_95_next_state), .CK(clk), .Q(RoundKey[95]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_95_MUX_inst_U1 ( .A(RoundKeyOutput[95]), .B(
        key[95]), .S(reset), .Z(KeyReg_Inst_ff_SDE_95_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_96_current_state_reg_U1 ( .A(RoundKey[96]), .ZN(
        KeyReg_Inst_ff_SDE_96_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_96_next_state), .CK(clk), .Q(RoundKey[96]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_96_MUX_inst_U1 ( .A(RoundKeyOutput[96]), .B(
        key[96]), .S(reset), .Z(KeyReg_Inst_ff_SDE_96_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_97_current_state_reg_U1 ( .A(RoundKey[97]), .ZN(
        KeyReg_Inst_ff_SDE_97_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_97_next_state), .CK(clk), .Q(RoundKey[97]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_97_MUX_inst_U1 ( .A(RoundKeyOutput[97]), .B(
        key[97]), .S(reset), .Z(KeyReg_Inst_ff_SDE_97_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_98_current_state_reg_U1 ( .A(RoundKey[98]), .ZN(
        KeyReg_Inst_ff_SDE_98_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_98_next_state), .CK(clk), .Q(RoundKey[98]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_98_MUX_inst_U1 ( .A(RoundKeyOutput[98]), .B(
        key[98]), .S(reset), .Z(KeyReg_Inst_ff_SDE_98_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_99_current_state_reg_U1 ( .A(RoundKey[99]), .ZN(
        KeyReg_Inst_ff_SDE_99_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_99_next_state), .CK(clk), .Q(RoundKey[99]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_99_MUX_inst_U1 ( .A(RoundKeyOutput[99]), .B(
        key[99]), .S(reset), .Z(KeyReg_Inst_ff_SDE_99_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_100_current_state_reg_U1 ( .A(RoundKey[100]), .ZN(
        KeyReg_Inst_ff_SDE_100_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_100_next_state), .CK(clk), .Q(RoundKey[100]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_100_MUX_inst_U1 ( .A(RoundKeyOutput[100]), .B(
        key[100]), .S(reset), .Z(KeyReg_Inst_ff_SDE_100_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_101_current_state_reg_U1 ( .A(RoundKey[101]), .ZN(
        KeyReg_Inst_ff_SDE_101_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_101_next_state), .CK(clk), .Q(RoundKey[101]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_101_MUX_inst_U1 ( .A(RoundKeyOutput[101]), .B(
        key[101]), .S(reset), .Z(KeyReg_Inst_ff_SDE_101_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_102_current_state_reg_U1 ( .A(RoundKey[102]), .ZN(
        KeyReg_Inst_ff_SDE_102_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_102_next_state), .CK(clk), .Q(RoundKey[102]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_102_MUX_inst_U1 ( .A(RoundKeyOutput[102]), .B(
        key[102]), .S(reset), .Z(KeyReg_Inst_ff_SDE_102_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_103_current_state_reg_U1 ( .A(RoundKey[103]), .ZN(
        KeyReg_Inst_ff_SDE_103_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_103_next_state), .CK(clk), .Q(RoundKey[103]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_103_MUX_inst_U1 ( .A(RoundKeyOutput[103]), .B(
        key[103]), .S(reset), .Z(KeyReg_Inst_ff_SDE_103_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_104_current_state_reg_U1 ( .A(RoundKey[104]), .ZN(
        KeyReg_Inst_ff_SDE_104_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_104_next_state), .CK(clk), .Q(RoundKey[104]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_104_MUX_inst_U1 ( .A(RoundKeyOutput[104]), .B(
        key[104]), .S(reset), .Z(KeyReg_Inst_ff_SDE_104_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_105_current_state_reg_U1 ( .A(RoundKey[105]), .ZN(
        KeyReg_Inst_ff_SDE_105_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_105_next_state), .CK(clk), .Q(RoundKey[105]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_105_MUX_inst_U1 ( .A(RoundKeyOutput[105]), .B(
        key[105]), .S(reset), .Z(KeyReg_Inst_ff_SDE_105_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_106_current_state_reg_U1 ( .A(RoundKey[106]), .ZN(
        KeyReg_Inst_ff_SDE_106_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_106_next_state), .CK(clk), .Q(RoundKey[106]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_106_MUX_inst_U1 ( .A(RoundKeyOutput[106]), .B(
        key[106]), .S(reset), .Z(KeyReg_Inst_ff_SDE_106_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_107_current_state_reg_U1 ( .A(RoundKey[107]), .ZN(
        KeyReg_Inst_ff_SDE_107_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_107_next_state), .CK(clk), .Q(RoundKey[107]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_107_MUX_inst_U1 ( .A(RoundKeyOutput[107]), .B(
        key[107]), .S(reset), .Z(KeyReg_Inst_ff_SDE_107_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_108_current_state_reg_U1 ( .A(RoundKey[108]), .ZN(
        KeyReg_Inst_ff_SDE_108_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_108_next_state), .CK(clk), .Q(RoundKey[108]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_108_MUX_inst_U1 ( .A(RoundKeyOutput[108]), .B(
        key[108]), .S(reset), .Z(KeyReg_Inst_ff_SDE_108_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_109_current_state_reg_U1 ( .A(RoundKey[109]), .ZN(
        KeyReg_Inst_ff_SDE_109_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_109_next_state), .CK(clk), .Q(RoundKey[109]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_109_MUX_inst_U1 ( .A(RoundKeyOutput[109]), .B(
        key[109]), .S(reset), .Z(KeyReg_Inst_ff_SDE_109_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_110_current_state_reg_U1 ( .A(RoundKey[110]), .ZN(
        KeyReg_Inst_ff_SDE_110_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_110_next_state), .CK(clk), .Q(RoundKey[110]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_110_MUX_inst_U1 ( .A(RoundKeyOutput[110]), .B(
        key[110]), .S(reset), .Z(KeyReg_Inst_ff_SDE_110_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_111_current_state_reg_U1 ( .A(RoundKey[111]), .ZN(
        KeyReg_Inst_ff_SDE_111_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_111_next_state), .CK(clk), .Q(RoundKey[111]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_111_MUX_inst_U1 ( .A(RoundKeyOutput[111]), .B(
        key[111]), .S(reset), .Z(KeyReg_Inst_ff_SDE_111_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_112_current_state_reg_U1 ( .A(RoundKey[112]), .ZN(
        KeyReg_Inst_ff_SDE_112_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_112_next_state), .CK(clk), .Q(RoundKey[112]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_112_MUX_inst_U1 ( .A(RoundKeyOutput[112]), .B(
        key[112]), .S(reset), .Z(KeyReg_Inst_ff_SDE_112_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_113_current_state_reg_U1 ( .A(RoundKey[113]), .ZN(
        KeyReg_Inst_ff_SDE_113_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_113_next_state), .CK(clk), .Q(RoundKey[113]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_113_MUX_inst_U1 ( .A(RoundKeyOutput[113]), .B(
        key[113]), .S(reset), .Z(KeyReg_Inst_ff_SDE_113_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_114_current_state_reg_U1 ( .A(RoundKey[114]), .ZN(
        KeyReg_Inst_ff_SDE_114_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_114_next_state), .CK(clk), .Q(RoundKey[114]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_114_MUX_inst_U1 ( .A(RoundKeyOutput[114]), .B(
        key[114]), .S(reset), .Z(KeyReg_Inst_ff_SDE_114_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_115_current_state_reg_U1 ( .A(RoundKey[115]), .ZN(
        KeyReg_Inst_ff_SDE_115_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_115_next_state), .CK(clk), .Q(RoundKey[115]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_115_MUX_inst_U1 ( .A(RoundKeyOutput[115]), .B(
        key[115]), .S(reset), .Z(KeyReg_Inst_ff_SDE_115_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_116_current_state_reg_U1 ( .A(RoundKey[116]), .ZN(
        KeyReg_Inst_ff_SDE_116_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_116_next_state), .CK(clk), .Q(RoundKey[116]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_116_MUX_inst_U1 ( .A(RoundKeyOutput[116]), .B(
        key[116]), .S(reset), .Z(KeyReg_Inst_ff_SDE_116_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_117_current_state_reg_U1 ( .A(RoundKey[117]), .ZN(
        KeyReg_Inst_ff_SDE_117_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_117_next_state), .CK(clk), .Q(RoundKey[117]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_117_MUX_inst_U1 ( .A(RoundKeyOutput[117]), .B(
        key[117]), .S(reset), .Z(KeyReg_Inst_ff_SDE_117_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_118_current_state_reg_U1 ( .A(RoundKey[118]), .ZN(
        KeyReg_Inst_ff_SDE_118_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_118_next_state), .CK(clk), .Q(RoundKey[118]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_118_MUX_inst_U1 ( .A(RoundKeyOutput[118]), .B(
        key[118]), .S(reset), .Z(KeyReg_Inst_ff_SDE_118_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_119_current_state_reg_U1 ( .A(RoundKey[119]), .ZN(
        KeyReg_Inst_ff_SDE_119_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_119_next_state), .CK(clk), .Q(RoundKey[119]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_119_MUX_inst_U1 ( .A(RoundKeyOutput[119]), .B(
        key[119]), .S(reset), .Z(KeyReg_Inst_ff_SDE_119_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_120_current_state_reg_U1 ( .A(RoundKey[120]), .ZN(
        KeyReg_Inst_ff_SDE_120_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_120_next_state), .CK(clk), .Q(RoundKey[120]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_120_MUX_inst_U1 ( .A(RoundKeyOutput[120]), .B(
        key[120]), .S(reset), .Z(KeyReg_Inst_ff_SDE_120_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_121_current_state_reg_U1 ( .A(RoundKey[121]), .ZN(
        KeyReg_Inst_ff_SDE_121_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_121_next_state), .CK(clk), .Q(RoundKey[121]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_121_MUX_inst_U1 ( .A(RoundKeyOutput[121]), .B(
        key[121]), .S(reset), .Z(KeyReg_Inst_ff_SDE_121_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_122_current_state_reg_U1 ( .A(RoundKey[122]), .ZN(
        KeyReg_Inst_ff_SDE_122_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_122_next_state), .CK(clk), .Q(RoundKey[122]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_122_MUX_inst_U1 ( .A(RoundKeyOutput[122]), .B(
        key[122]), .S(reset), .Z(KeyReg_Inst_ff_SDE_122_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_123_current_state_reg_U1 ( .A(RoundKey[123]), .ZN(
        KeyReg_Inst_ff_SDE_123_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_123_next_state), .CK(clk), .Q(RoundKey[123]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_123_MUX_inst_U1 ( .A(RoundKeyOutput[123]), .B(
        key[123]), .S(reset), .Z(KeyReg_Inst_ff_SDE_123_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_124_current_state_reg_U1 ( .A(RoundKey[124]), .ZN(
        KeyReg_Inst_ff_SDE_124_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_124_next_state), .CK(clk), .Q(RoundKey[124]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_124_MUX_inst_U1 ( .A(RoundKeyOutput[124]), .B(
        key[124]), .S(reset), .Z(KeyReg_Inst_ff_SDE_124_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_125_current_state_reg_U1 ( .A(RoundKey[125]), .ZN(
        KeyReg_Inst_ff_SDE_125_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_125_next_state), .CK(clk), .Q(RoundKey[125]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_125_MUX_inst_U1 ( .A(RoundKeyOutput[125]), .B(
        key[125]), .S(reset), .Z(KeyReg_Inst_ff_SDE_125_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_126_current_state_reg_U1 ( .A(RoundKey[126]), .ZN(
        KeyReg_Inst_ff_SDE_126_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_126_next_state), .CK(clk), .Q(RoundKey[126]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_126_MUX_inst_U1 ( .A(RoundKeyOutput[126]), .B(
        key[126]), .S(reset), .Z(KeyReg_Inst_ff_SDE_126_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_127_current_state_reg_U1 ( .A(RoundKey[127]), .ZN(
        KeyReg_Inst_ff_SDE_127_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_127_next_state), .CK(clk), .Q(RoundKey[127]), .QN()
         );
  MUX2_X1 KeyReg_Inst_ff_SDE_127_MUX_inst_U1 ( .A(RoundKeyOutput[127]), .B(
        key[127]), .S(reset), .Z(KeyReg_Inst_ff_SDE_127_next_state) );
  XOR2_X1 KeyExpansionIns_U128 ( .A(KSSubBytesInput[9]), .B(
        KeyExpansionOutput[41]), .Z(KeyExpansionOutput[9]) );
  XOR2_X1 KeyExpansionIns_U127 ( .A(KSSubBytesInput[8]), .B(
        KeyExpansionOutput[40]), .Z(KeyExpansionOutput[8]) );
  XOR2_X1 KeyExpansionIns_U126 ( .A(KSSubBytesInput[23]), .B(
        KeyExpansionOutput[39]), .Z(KeyExpansionOutput[7]) );
  XOR2_X1 KeyExpansionIns_U125 ( .A(KSSubBytesInput[22]), .B(
        KeyExpansionOutput[38]), .Z(KeyExpansionOutput[6]) );
  XOR2_X1 KeyExpansionIns_U124 ( .A(KSSubBytesInput[21]), .B(
        KeyExpansionOutput[37]), .Z(KeyExpansionOutput[5]) );
  XOR2_X1 KeyExpansionIns_U123 ( .A(KSSubBytesInput[20]), .B(
        KeyExpansionOutput[36]), .Z(KeyExpansionOutput[4]) );
  XOR2_X1 KeyExpansionIns_U122 ( .A(RoundKey[41]), .B(KeyExpansionOutput[73]), 
        .Z(KeyExpansionOutput[41]) );
  XOR2_X1 KeyExpansionIns_U121 ( .A(RoundKey[73]), .B(KeyExpansionOutput[105]), 
        .Z(KeyExpansionOutput[73]) );
  XOR2_X1 KeyExpansionIns_U120 ( .A(RoundKey[40]), .B(KeyExpansionOutput[72]), 
        .Z(KeyExpansionOutput[40]) );
  XOR2_X1 KeyExpansionIns_U119 ( .A(RoundKey[72]), .B(KeyExpansionOutput[104]), 
        .Z(KeyExpansionOutput[72]) );
  XOR2_X1 KeyExpansionIns_U118 ( .A(KSSubBytesInput[19]), .B(
        KeyExpansionOutput[35]), .Z(KeyExpansionOutput[3]) );
  XOR2_X1 KeyExpansionIns_U117 ( .A(RoundKey[39]), .B(KeyExpansionOutput[71]), 
        .Z(KeyExpansionOutput[39]) );
  XOR2_X1 KeyExpansionIns_U116 ( .A(RoundKey[71]), .B(KeyExpansionOutput[103]), 
        .Z(KeyExpansionOutput[71]) );
  XOR2_X1 KeyExpansionIns_U115 ( .A(RoundKey[38]), .B(KeyExpansionOutput[70]), 
        .Z(KeyExpansionOutput[38]) );
  XOR2_X1 KeyExpansionIns_U114 ( .A(RoundKey[70]), .B(KeyExpansionOutput[102]), 
        .Z(KeyExpansionOutput[70]) );
  XOR2_X1 KeyExpansionIns_U113 ( .A(RoundKey[37]), .B(KeyExpansionOutput[69]), 
        .Z(KeyExpansionOutput[37]) );
  XOR2_X1 KeyExpansionIns_U112 ( .A(RoundKey[69]), .B(KeyExpansionOutput[101]), 
        .Z(KeyExpansionOutput[69]) );
  XOR2_X1 KeyExpansionIns_U111 ( .A(RoundKey[36]), .B(KeyExpansionOutput[68]), 
        .Z(KeyExpansionOutput[36]) );
  XOR2_X1 KeyExpansionIns_U110 ( .A(RoundKey[68]), .B(KeyExpansionOutput[100]), 
        .Z(KeyExpansionOutput[68]) );
  XOR2_X1 KeyExpansionIns_U109 ( .A(RoundKey[35]), .B(KeyExpansionOutput[67]), 
        .Z(KeyExpansionOutput[35]) );
  XOR2_X1 KeyExpansionIns_U108 ( .A(RoundKey[67]), .B(KeyExpansionOutput[99]), 
        .Z(KeyExpansionOutput[67]) );
  XOR2_X1 KeyExpansionIns_U107 ( .A(RoundKey[99]), .B(KeyExpansionIns_tmp[3]), 
        .Z(KeyExpansionOutput[99]) );
  XOR2_X1 KeyExpansionIns_U106 ( .A(KSSubBytesInput[31]), .B(
        KeyExpansionOutput[63]), .Z(KeyExpansionOutput[31]) );
  XOR2_X1 KeyExpansionIns_U105 ( .A(RoundKey[63]), .B(KeyExpansionOutput[95]), 
        .Z(KeyExpansionOutput[63]) );
  XOR2_X1 KeyExpansionIns_U104 ( .A(RoundKey[95]), .B(KeyExpansionOutput[127]), 
        .Z(KeyExpansionOutput[95]) );
  XOR2_X1 KeyExpansionIns_U103 ( .A(KSSubBytesInput[30]), .B(
        KeyExpansionOutput[62]), .Z(KeyExpansionOutput[30]) );
  XOR2_X1 KeyExpansionIns_U102 ( .A(RoundKey[62]), .B(KeyExpansionOutput[94]), 
        .Z(KeyExpansionOutput[62]) );
  XOR2_X1 KeyExpansionIns_U101 ( .A(RoundKey[94]), .B(KeyExpansionOutput[126]), 
        .Z(KeyExpansionOutput[94]) );
  XOR2_X1 KeyExpansionIns_U100 ( .A(KSSubBytesInput[18]), .B(
        KeyExpansionOutput[34]), .Z(KeyExpansionOutput[2]) );
  XOR2_X1 KeyExpansionIns_U99 ( .A(RoundKey[34]), .B(KeyExpansionOutput[66]), 
        .Z(KeyExpansionOutput[34]) );
  XOR2_X1 KeyExpansionIns_U98 ( .A(RoundKey[66]), .B(KeyExpansionOutput[98]), 
        .Z(KeyExpansionOutput[66]) );
  XOR2_X1 KeyExpansionIns_U97 ( .A(RoundKey[98]), .B(KeyExpansionIns_tmp[2]), 
        .Z(KeyExpansionOutput[98]) );
  XOR2_X1 KeyExpansionIns_U96 ( .A(KSSubBytesInput[29]), .B(
        KeyExpansionOutput[61]), .Z(KeyExpansionOutput[29]) );
  XOR2_X1 KeyExpansionIns_U95 ( .A(RoundKey[61]), .B(KeyExpansionOutput[93]), 
        .Z(KeyExpansionOutput[61]) );
  XOR2_X1 KeyExpansionIns_U94 ( .A(RoundKey[93]), .B(KeyExpansionOutput[125]), 
        .Z(KeyExpansionOutput[93]) );
  XOR2_X1 KeyExpansionIns_U93 ( .A(KSSubBytesInput[28]), .B(
        KeyExpansionOutput[60]), .Z(KeyExpansionOutput[28]) );
  XOR2_X1 KeyExpansionIns_U92 ( .A(RoundKey[60]), .B(KeyExpansionOutput[92]), 
        .Z(KeyExpansionOutput[60]) );
  XOR2_X1 KeyExpansionIns_U91 ( .A(RoundKey[92]), .B(KeyExpansionOutput[124]), 
        .Z(KeyExpansionOutput[92]) );
  XOR2_X1 KeyExpansionIns_U90 ( .A(KSSubBytesInput[27]), .B(
        KeyExpansionOutput[59]), .Z(KeyExpansionOutput[27]) );
  XOR2_X1 KeyExpansionIns_U89 ( .A(RoundKey[59]), .B(KeyExpansionOutput[91]), 
        .Z(KeyExpansionOutput[59]) );
  XOR2_X1 KeyExpansionIns_U88 ( .A(RoundKey[91]), .B(KeyExpansionOutput[123]), 
        .Z(KeyExpansionOutput[91]) );
  XOR2_X1 KeyExpansionIns_U87 ( .A(KSSubBytesInput[26]), .B(
        KeyExpansionOutput[58]), .Z(KeyExpansionOutput[26]) );
  XOR2_X1 KeyExpansionIns_U86 ( .A(RoundKey[58]), .B(KeyExpansionOutput[90]), 
        .Z(KeyExpansionOutput[58]) );
  XOR2_X1 KeyExpansionIns_U85 ( .A(RoundKey[90]), .B(KeyExpansionOutput[122]), 
        .Z(KeyExpansionOutput[90]) );
  XOR2_X1 KeyExpansionIns_U84 ( .A(KSSubBytesInput[25]), .B(
        KeyExpansionOutput[57]), .Z(KeyExpansionOutput[25]) );
  XOR2_X1 KeyExpansionIns_U83 ( .A(RoundKey[57]), .B(KeyExpansionOutput[89]), 
        .Z(KeyExpansionOutput[57]) );
  XOR2_X1 KeyExpansionIns_U82 ( .A(RoundKey[89]), .B(KeyExpansionOutput[121]), 
        .Z(KeyExpansionOutput[89]) );
  XOR2_X1 KeyExpansionIns_U81 ( .A(KSSubBytesInput[24]), .B(
        KeyExpansionOutput[56]), .Z(KeyExpansionOutput[24]) );
  XOR2_X1 KeyExpansionIns_U80 ( .A(RoundKey[56]), .B(KeyExpansionOutput[88]), 
        .Z(KeyExpansionOutput[56]) );
  XOR2_X1 KeyExpansionIns_U79 ( .A(RoundKey[88]), .B(KeyExpansionOutput[120]), 
        .Z(KeyExpansionOutput[88]) );
  XOR2_X1 KeyExpansionIns_U78 ( .A(KSSubBytesInput[7]), .B(
        KeyExpansionOutput[55]), .Z(KeyExpansionOutput[23]) );
  XOR2_X1 KeyExpansionIns_U77 ( .A(RoundKey[55]), .B(KeyExpansionOutput[87]), 
        .Z(KeyExpansionOutput[55]) );
  XOR2_X1 KeyExpansionIns_U76 ( .A(RoundKey[87]), .B(KeyExpansionOutput[119]), 
        .Z(KeyExpansionOutput[87]) );
  XOR2_X1 KeyExpansionIns_U75 ( .A(KSSubBytesInput[6]), .B(
        KeyExpansionOutput[54]), .Z(KeyExpansionOutput[22]) );
  XOR2_X1 KeyExpansionIns_U74 ( .A(RoundKey[54]), .B(KeyExpansionOutput[86]), 
        .Z(KeyExpansionOutput[54]) );
  XOR2_X1 KeyExpansionIns_U73 ( .A(RoundKey[86]), .B(KeyExpansionOutput[118]), 
        .Z(KeyExpansionOutput[86]) );
  XOR2_X1 KeyExpansionIns_U72 ( .A(KSSubBytesInput[5]), .B(
        KeyExpansionOutput[53]), .Z(KeyExpansionOutput[21]) );
  XOR2_X1 KeyExpansionIns_U71 ( .A(RoundKey[53]), .B(KeyExpansionOutput[85]), 
        .Z(KeyExpansionOutput[53]) );
  XOR2_X1 KeyExpansionIns_U70 ( .A(RoundKey[85]), .B(KeyExpansionOutput[117]), 
        .Z(KeyExpansionOutput[85]) );
  XOR2_X1 KeyExpansionIns_U69 ( .A(KSSubBytesInput[4]), .B(
        KeyExpansionOutput[52]), .Z(KeyExpansionOutput[20]) );
  XOR2_X1 KeyExpansionIns_U68 ( .A(RoundKey[52]), .B(KeyExpansionOutput[84]), 
        .Z(KeyExpansionOutput[52]) );
  XOR2_X1 KeyExpansionIns_U67 ( .A(RoundKey[84]), .B(KeyExpansionOutput[116]), 
        .Z(KeyExpansionOutput[84]) );
  XOR2_X1 KeyExpansionIns_U66 ( .A(KSSubBytesInput[17]), .B(
        KeyExpansionOutput[33]), .Z(KeyExpansionOutput[1]) );
  XOR2_X1 KeyExpansionIns_U65 ( .A(RoundKey[33]), .B(KeyExpansionOutput[65]), 
        .Z(KeyExpansionOutput[33]) );
  XOR2_X1 KeyExpansionIns_U64 ( .A(RoundKey[65]), .B(KeyExpansionOutput[97]), 
        .Z(KeyExpansionOutput[65]) );
  XOR2_X1 KeyExpansionIns_U63 ( .A(RoundKey[97]), .B(KeyExpansionIns_tmp[1]), 
        .Z(KeyExpansionOutput[97]) );
  XOR2_X1 KeyExpansionIns_U62 ( .A(KSSubBytesInput[3]), .B(
        KeyExpansionOutput[51]), .Z(KeyExpansionOutput[19]) );
  XOR2_X1 KeyExpansionIns_U61 ( .A(RoundKey[51]), .B(KeyExpansionOutput[83]), 
        .Z(KeyExpansionOutput[51]) );
  XOR2_X1 KeyExpansionIns_U60 ( .A(RoundKey[83]), .B(KeyExpansionOutput[115]), 
        .Z(KeyExpansionOutput[83]) );
  XOR2_X1 KeyExpansionIns_U59 ( .A(KSSubBytesInput[2]), .B(
        KeyExpansionOutput[50]), .Z(KeyExpansionOutput[18]) );
  XOR2_X1 KeyExpansionIns_U58 ( .A(RoundKey[50]), .B(KeyExpansionOutput[82]), 
        .Z(KeyExpansionOutput[50]) );
  XOR2_X1 KeyExpansionIns_U57 ( .A(RoundKey[82]), .B(KeyExpansionOutput[114]), 
        .Z(KeyExpansionOutput[82]) );
  XOR2_X1 KeyExpansionIns_U56 ( .A(KSSubBytesInput[1]), .B(
        KeyExpansionOutput[49]), .Z(KeyExpansionOutput[17]) );
  XOR2_X1 KeyExpansionIns_U55 ( .A(RoundKey[49]), .B(KeyExpansionOutput[81]), 
        .Z(KeyExpansionOutput[49]) );
  XOR2_X1 KeyExpansionIns_U54 ( .A(RoundKey[81]), .B(KeyExpansionOutput[113]), 
        .Z(KeyExpansionOutput[81]) );
  XOR2_X1 KeyExpansionIns_U53 ( .A(KSSubBytesInput[0]), .B(
        KeyExpansionOutput[48]), .Z(KeyExpansionOutput[16]) );
  XOR2_X1 KeyExpansionIns_U52 ( .A(RoundKey[48]), .B(KeyExpansionOutput[80]), 
        .Z(KeyExpansionOutput[48]) );
  XOR2_X1 KeyExpansionIns_U51 ( .A(RoundKey[80]), .B(KeyExpansionOutput[112]), 
        .Z(KeyExpansionOutput[80]) );
  XOR2_X1 KeyExpansionIns_U50 ( .A(KSSubBytesInput[15]), .B(
        KeyExpansionOutput[47]), .Z(KeyExpansionOutput[15]) );
  XOR2_X1 KeyExpansionIns_U49 ( .A(RoundKey[47]), .B(KeyExpansionOutput[79]), 
        .Z(KeyExpansionOutput[47]) );
  XOR2_X1 KeyExpansionIns_U48 ( .A(RoundKey[79]), .B(KeyExpansionOutput[111]), 
        .Z(KeyExpansionOutput[79]) );
  XOR2_X1 KeyExpansionIns_U47 ( .A(KSSubBytesInput[14]), .B(
        KeyExpansionOutput[46]), .Z(KeyExpansionOutput[14]) );
  XOR2_X1 KeyExpansionIns_U46 ( .A(RoundKey[46]), .B(KeyExpansionOutput[78]), 
        .Z(KeyExpansionOutput[46]) );
  XOR2_X1 KeyExpansionIns_U45 ( .A(RoundKey[78]), .B(KeyExpansionOutput[110]), 
        .Z(KeyExpansionOutput[78]) );
  XOR2_X1 KeyExpansionIns_U44 ( .A(KSSubBytesInput[13]), .B(
        KeyExpansionOutput[45]), .Z(KeyExpansionOutput[13]) );
  XOR2_X1 KeyExpansionIns_U43 ( .A(RoundKey[45]), .B(KeyExpansionOutput[77]), 
        .Z(KeyExpansionOutput[45]) );
  XOR2_X1 KeyExpansionIns_U42 ( .A(RoundKey[77]), .B(KeyExpansionOutput[109]), 
        .Z(KeyExpansionOutput[77]) );
  XOR2_X1 KeyExpansionIns_U41 ( .A(KSSubBytesInput[12]), .B(
        KeyExpansionOutput[44]), .Z(KeyExpansionOutput[12]) );
  XOR2_X1 KeyExpansionIns_U40 ( .A(RoundKey[44]), .B(KeyExpansionOutput[76]), 
        .Z(KeyExpansionOutput[44]) );
  XOR2_X1 KeyExpansionIns_U39 ( .A(RoundKey[76]), .B(KeyExpansionOutput[108]), 
        .Z(KeyExpansionOutput[76]) );
  XOR2_X1 KeyExpansionIns_U38 ( .A(RoundKey[127]), .B(KeyExpansionIns_tmp[31]), 
        .Z(KeyExpansionOutput[127]) );
  XOR2_X1 KeyExpansionIns_U37 ( .A(RoundKey[126]), .B(KeyExpansionIns_tmp[30]), 
        .Z(KeyExpansionOutput[126]) );
  XOR2_X1 KeyExpansionIns_U36 ( .A(RoundKey[125]), .B(KeyExpansionIns_tmp[29]), 
        .Z(KeyExpansionOutput[125]) );
  XOR2_X1 KeyExpansionIns_U35 ( .A(RoundKey[124]), .B(KeyExpansionIns_tmp[28]), 
        .Z(KeyExpansionOutput[124]) );
  XOR2_X1 KeyExpansionIns_U34 ( .A(RoundKey[123]), .B(KeyExpansionIns_tmp[27]), 
        .Z(KeyExpansionOutput[123]) );
  XOR2_X1 KeyExpansionIns_U33 ( .A(RoundKey[122]), .B(KeyExpansionIns_tmp[26]), 
        .Z(KeyExpansionOutput[122]) );
  XOR2_X1 KeyExpansionIns_U32 ( .A(RoundKey[121]), .B(KeyExpansionIns_tmp[25]), 
        .Z(KeyExpansionOutput[121]) );
  XOR2_X1 KeyExpansionIns_U31 ( .A(RoundKey[120]), .B(KeyExpansionIns_tmp[24]), 
        .Z(KeyExpansionOutput[120]) );
  XOR2_X1 KeyExpansionIns_U30 ( .A(KSSubBytesInput[11]), .B(
        KeyExpansionOutput[43]), .Z(KeyExpansionOutput[11]) );
  XOR2_X1 KeyExpansionIns_U29 ( .A(RoundKey[43]), .B(KeyExpansionOutput[75]), 
        .Z(KeyExpansionOutput[43]) );
  XOR2_X1 KeyExpansionIns_U28 ( .A(RoundKey[75]), .B(KeyExpansionOutput[107]), 
        .Z(KeyExpansionOutput[75]) );
  XOR2_X1 KeyExpansionIns_U27 ( .A(RoundKey[119]), .B(KeyExpansionIns_tmp[23]), 
        .Z(KeyExpansionOutput[119]) );
  XOR2_X1 KeyExpansionIns_U26 ( .A(RoundKey[118]), .B(KeyExpansionIns_tmp[22]), 
        .Z(KeyExpansionOutput[118]) );
  XOR2_X1 KeyExpansionIns_U25 ( .A(RoundKey[117]), .B(KeyExpansionIns_tmp[21]), 
        .Z(KeyExpansionOutput[117]) );
  XOR2_X1 KeyExpansionIns_U24 ( .A(RoundKey[116]), .B(KeyExpansionIns_tmp[20]), 
        .Z(KeyExpansionOutput[116]) );
  XOR2_X1 KeyExpansionIns_U23 ( .A(RoundKey[115]), .B(KeyExpansionIns_tmp[19]), 
        .Z(KeyExpansionOutput[115]) );
  XOR2_X1 KeyExpansionIns_U22 ( .A(RoundKey[114]), .B(KeyExpansionIns_tmp[18]), 
        .Z(KeyExpansionOutput[114]) );
  XOR2_X1 KeyExpansionIns_U21 ( .A(RoundKey[113]), .B(KeyExpansionIns_tmp[17]), 
        .Z(KeyExpansionOutput[113]) );
  XOR2_X1 KeyExpansionIns_U20 ( .A(RoundKey[112]), .B(KeyExpansionIns_tmp[16]), 
        .Z(KeyExpansionOutput[112]) );
  XOR2_X1 KeyExpansionIns_U19 ( .A(RoundKey[111]), .B(KeyExpansionIns_tmp[15]), 
        .Z(KeyExpansionOutput[111]) );
  XOR2_X1 KeyExpansionIns_U18 ( .A(RoundKey[110]), .B(KeyExpansionIns_tmp[14]), 
        .Z(KeyExpansionOutput[110]) );
  XOR2_X1 KeyExpansionIns_U17 ( .A(KSSubBytesInput[10]), .B(
        KeyExpansionOutput[42]), .Z(KeyExpansionOutput[10]) );
  XOR2_X1 KeyExpansionIns_U16 ( .A(RoundKey[42]), .B(KeyExpansionOutput[74]), 
        .Z(KeyExpansionOutput[42]) );
  XOR2_X1 KeyExpansionIns_U15 ( .A(RoundKey[74]), .B(KeyExpansionOutput[106]), 
        .Z(KeyExpansionOutput[74]) );
  XOR2_X1 KeyExpansionIns_U14 ( .A(RoundKey[109]), .B(KeyExpansionIns_tmp[13]), 
        .Z(KeyExpansionOutput[109]) );
  XOR2_X1 KeyExpansionIns_U13 ( .A(RoundKey[108]), .B(KeyExpansionIns_tmp[12]), 
        .Z(KeyExpansionOutput[108]) );
  XOR2_X1 KeyExpansionIns_U12 ( .A(RoundKey[107]), .B(KeyExpansionIns_tmp[11]), 
        .Z(KeyExpansionOutput[107]) );
  XOR2_X1 KeyExpansionIns_U11 ( .A(RoundKey[106]), .B(KeyExpansionIns_tmp[10]), 
        .Z(KeyExpansionOutput[106]) );
  XOR2_X1 KeyExpansionIns_U10 ( .A(RoundKey[105]), .B(KeyExpansionIns_tmp[9]), 
        .Z(KeyExpansionOutput[105]) );
  XOR2_X1 KeyExpansionIns_U9 ( .A(RoundKey[104]), .B(KeyExpansionIns_tmp[8]), 
        .Z(KeyExpansionOutput[104]) );
  XOR2_X1 KeyExpansionIns_U8 ( .A(RoundKey[103]), .B(KeyExpansionIns_tmp[7]), 
        .Z(KeyExpansionOutput[103]) );
  XOR2_X1 KeyExpansionIns_U7 ( .A(RoundKey[102]), .B(KeyExpansionIns_tmp[6]), 
        .Z(KeyExpansionOutput[102]) );
  XOR2_X1 KeyExpansionIns_U6 ( .A(RoundKey[101]), .B(KeyExpansionIns_tmp[5]), 
        .Z(KeyExpansionOutput[101]) );
  XOR2_X1 KeyExpansionIns_U5 ( .A(RoundKey[100]), .B(KeyExpansionIns_tmp[4]), 
        .Z(KeyExpansionOutput[100]) );
  XOR2_X1 KeyExpansionIns_U4 ( .A(KSSubBytesInput[16]), .B(
        KeyExpansionOutput[32]), .Z(KeyExpansionOutput[0]) );
  XOR2_X1 KeyExpansionIns_U3 ( .A(RoundKey[32]), .B(KeyExpansionOutput[64]), 
        .Z(KeyExpansionOutput[32]) );
  XOR2_X1 KeyExpansionIns_U2 ( .A(RoundKey[64]), .B(KeyExpansionOutput[96]), 
        .Z(KeyExpansionOutput[64]) );
  XOR2_X1 KeyExpansionIns_U1 ( .A(RoundKey[96]), .B(KeyExpansionIns_tmp[0]), 
        .Z(KeyExpansionOutput[96]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U8 ( .A(Rcon[7]), .B(
        MixColumnsIns_DoubleBytes[0]), .Z(KeyExpansionIns_tmp[31]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U7 ( .A(Rcon[6]), .B(
        MixColumnsIns_DoubleBytes[7]), .Z(KeyExpansionIns_tmp[30]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U6 ( .A(Rcon[5]), .B(
        MixColumnsIns_DoubleBytes[6]), .Z(KeyExpansionIns_tmp[29]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U5 ( .A(Rcon[4]), .B(
        MixColumnsIns_DoubleBytes[5]), .Z(KeyExpansionIns_tmp[28]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U4 ( .A(Rcon[3]), .B(
        SubBytesOutput[3]), .Z(KeyExpansionIns_tmp[27]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U3 ( .A(Rcon[2]), .B(
        SubBytesOutput[2]), .Z(KeyExpansionIns_tmp[26]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U2 ( .A(Rcon[1]), .B(
        MixColumnsIns_DoubleBytes[2]), .Z(KeyExpansionIns_tmp[25]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U1 ( .A(Rcon[0]), .B(
        SubBytesOutput[0]), .Z(KeyExpansionIns_tmp[24]) );
  INV_X1 MuxKeyExpansion_U8 ( .A(MuxKeyExpansion_n21), .ZN(MuxKeyExpansion_n14) );
  INV_X1 MuxKeyExpansion_U7 ( .A(AKSRnotDone), .ZN(MuxKeyExpansion_n21) );
  INV_X1 MuxKeyExpansion_U6 ( .A(MuxKeyExpansion_n21), .ZN(MuxKeyExpansion_n16) );
  INV_X1 MuxKeyExpansion_U5 ( .A(MuxKeyExpansion_n21), .ZN(MuxKeyExpansion_n17) );
  INV_X1 MuxKeyExpansion_U4 ( .A(MuxKeyExpansion_n21), .ZN(MuxKeyExpansion_n18) );
  INV_X1 MuxKeyExpansion_U3 ( .A(MuxKeyExpansion_n21), .ZN(MuxKeyExpansion_n19) );
  INV_X1 MuxKeyExpansion_U2 ( .A(MuxKeyExpansion_n21), .ZN(MuxKeyExpansion_n20) );
  INV_X1 MuxKeyExpansion_U1 ( .A(MuxKeyExpansion_n21), .ZN(MuxKeyExpansion_n15) );
  MUX2_X1 MuxKeyExpansion_mux_inst_0_U1 ( .A(KSSubBytesInput[16]), .B(
        KeyExpansionOutput[0]), .S(MuxKeyExpansion_n15), .Z(RoundKeyOutput[0])
         );
  MUX2_X1 MuxKeyExpansion_mux_inst_1_U1 ( .A(KSSubBytesInput[17]), .B(
        KeyExpansionOutput[1]), .S(MuxKeyExpansion_n16), .Z(RoundKeyOutput[1])
         );
  MUX2_X1 MuxKeyExpansion_mux_inst_2_U1 ( .A(KSSubBytesInput[18]), .B(
        KeyExpansionOutput[2]), .S(MuxKeyExpansion_n17), .Z(RoundKeyOutput[2])
         );
  MUX2_X1 MuxKeyExpansion_mux_inst_3_U1 ( .A(KSSubBytesInput[19]), .B(
        KeyExpansionOutput[3]), .S(MuxKeyExpansion_n18), .Z(RoundKeyOutput[3])
         );
  MUX2_X1 MuxKeyExpansion_mux_inst_4_U1 ( .A(KSSubBytesInput[20]), .B(
        KeyExpansionOutput[4]), .S(MuxKeyExpansion_n19), .Z(RoundKeyOutput[4])
         );
  MUX2_X1 MuxKeyExpansion_mux_inst_5_U1 ( .A(KSSubBytesInput[21]), .B(
        KeyExpansionOutput[5]), .S(MuxKeyExpansion_n20), .Z(RoundKeyOutput[5])
         );
  MUX2_X1 MuxKeyExpansion_mux_inst_6_U1 ( .A(KSSubBytesInput[22]), .B(
        KeyExpansionOutput[6]), .S(MuxKeyExpansion_n16), .Z(RoundKeyOutput[6])
         );
  MUX2_X1 MuxKeyExpansion_mux_inst_7_U1 ( .A(KSSubBytesInput[23]), .B(
        KeyExpansionOutput[7]), .S(MuxKeyExpansion_n18), .Z(RoundKeyOutput[7])
         );
  MUX2_X1 MuxKeyExpansion_mux_inst_8_U1 ( .A(KSSubBytesInput[8]), .B(
        KeyExpansionOutput[8]), .S(MuxKeyExpansion_n15), .Z(RoundKeyOutput[8])
         );
  MUX2_X1 MuxKeyExpansion_mux_inst_9_U1 ( .A(KSSubBytesInput[9]), .B(
        KeyExpansionOutput[9]), .S(MuxKeyExpansion_n16), .Z(RoundKeyOutput[9])
         );
  MUX2_X1 MuxKeyExpansion_mux_inst_10_U1 ( .A(KSSubBytesInput[10]), .B(
        KeyExpansionOutput[10]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[10]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_11_U1 ( .A(KSSubBytesInput[11]), .B(
        KeyExpansionOutput[11]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[11]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_12_U1 ( .A(KSSubBytesInput[12]), .B(
        KeyExpansionOutput[12]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[12]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_13_U1 ( .A(KSSubBytesInput[13]), .B(
        KeyExpansionOutput[13]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[13]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_14_U1 ( .A(KSSubBytesInput[14]), .B(
        KeyExpansionOutput[14]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[14]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_15_U1 ( .A(KSSubBytesInput[15]), .B(
        KeyExpansionOutput[15]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[15]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_16_U1 ( .A(KSSubBytesInput[0]), .B(
        KeyExpansionOutput[16]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[16]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_17_U1 ( .A(KSSubBytesInput[1]), .B(
        KeyExpansionOutput[17]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[17]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_18_U1 ( .A(KSSubBytesInput[2]), .B(
        KeyExpansionOutput[18]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[18]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_19_U1 ( .A(KSSubBytesInput[3]), .B(
        KeyExpansionOutput[19]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[19]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_20_U1 ( .A(KSSubBytesInput[4]), .B(
        KeyExpansionOutput[20]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[20]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_21_U1 ( .A(KSSubBytesInput[5]), .B(
        KeyExpansionOutput[21]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[21]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_22_U1 ( .A(KSSubBytesInput[6]), .B(
        KeyExpansionOutput[22]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[22]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_23_U1 ( .A(KSSubBytesInput[7]), .B(
        KeyExpansionOutput[23]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[23]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_24_U1 ( .A(KSSubBytesInput[24]), .B(
        KeyExpansionOutput[24]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[24]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_25_U1 ( .A(KSSubBytesInput[25]), .B(
        KeyExpansionOutput[25]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[25]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_26_U1 ( .A(KSSubBytesInput[26]), .B(
        KeyExpansionOutput[26]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[26]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_27_U1 ( .A(KSSubBytesInput[27]), .B(
        KeyExpansionOutput[27]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[27]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_28_U1 ( .A(KSSubBytesInput[28]), .B(
        KeyExpansionOutput[28]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[28]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_29_U1 ( .A(KSSubBytesInput[29]), .B(
        KeyExpansionOutput[29]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[29]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_30_U1 ( .A(KSSubBytesInput[30]), .B(
        KeyExpansionOutput[30]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[30]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_31_U1 ( .A(KSSubBytesInput[31]), .B(
        KeyExpansionOutput[31]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[31]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_32_U1 ( .A(RoundKey[32]), .B(
        KeyExpansionOutput[32]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[32]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_33_U1 ( .A(RoundKey[33]), .B(
        KeyExpansionOutput[33]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[33]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_34_U1 ( .A(RoundKey[34]), .B(
        KeyExpansionOutput[34]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[34]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_35_U1 ( .A(RoundKey[35]), .B(
        KeyExpansionOutput[35]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[35]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_36_U1 ( .A(RoundKey[36]), .B(
        KeyExpansionOutput[36]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[36]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_37_U1 ( .A(RoundKey[37]), .B(
        KeyExpansionOutput[37]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[37]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_38_U1 ( .A(RoundKey[38]), .B(
        KeyExpansionOutput[38]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[38]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_39_U1 ( .A(RoundKey[39]), .B(
        KeyExpansionOutput[39]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[39]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_40_U1 ( .A(RoundKey[40]), .B(
        KeyExpansionOutput[40]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[40]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_41_U1 ( .A(RoundKey[41]), .B(
        KeyExpansionOutput[41]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[41]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_42_U1 ( .A(RoundKey[42]), .B(
        KeyExpansionOutput[42]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[42]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_43_U1 ( .A(RoundKey[43]), .B(
        KeyExpansionOutput[43]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[43]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_44_U1 ( .A(RoundKey[44]), .B(
        KeyExpansionOutput[44]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[44]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_45_U1 ( .A(RoundKey[45]), .B(
        KeyExpansionOutput[45]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[45]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_46_U1 ( .A(RoundKey[46]), .B(
        KeyExpansionOutput[46]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[46]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_47_U1 ( .A(RoundKey[47]), .B(
        KeyExpansionOutput[47]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[47]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_48_U1 ( .A(RoundKey[48]), .B(
        KeyExpansionOutput[48]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[48]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_49_U1 ( .A(RoundKey[49]), .B(
        KeyExpansionOutput[49]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[49]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_50_U1 ( .A(RoundKey[50]), .B(
        KeyExpansionOutput[50]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[50]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_51_U1 ( .A(RoundKey[51]), .B(
        KeyExpansionOutput[51]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[51]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_52_U1 ( .A(RoundKey[52]), .B(
        KeyExpansionOutput[52]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[52]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_53_U1 ( .A(RoundKey[53]), .B(
        KeyExpansionOutput[53]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[53]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_54_U1 ( .A(RoundKey[54]), .B(
        KeyExpansionOutput[54]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[54]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_55_U1 ( .A(RoundKey[55]), .B(
        KeyExpansionOutput[55]), .S(MuxKeyExpansion_n20), .Z(
        RoundKeyOutput[55]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_56_U1 ( .A(RoundKey[56]), .B(
        KeyExpansionOutput[56]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[56]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_57_U1 ( .A(RoundKey[57]), .B(
        KeyExpansionOutput[57]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[57]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_58_U1 ( .A(RoundKey[58]), .B(
        KeyExpansionOutput[58]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[58]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_59_U1 ( .A(RoundKey[59]), .B(
        KeyExpansionOutput[59]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[59]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_60_U1 ( .A(RoundKey[60]), .B(
        KeyExpansionOutput[60]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[60]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_61_U1 ( .A(RoundKey[61]), .B(
        KeyExpansionOutput[61]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[61]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_62_U1 ( .A(RoundKey[62]), .B(
        KeyExpansionOutput[62]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[62]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_63_U1 ( .A(RoundKey[63]), .B(
        KeyExpansionOutput[63]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[63]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_64_U1 ( .A(RoundKey[64]), .B(
        KeyExpansionOutput[64]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[64]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_65_U1 ( .A(RoundKey[65]), .B(
        KeyExpansionOutput[65]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[65]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_66_U1 ( .A(RoundKey[66]), .B(
        KeyExpansionOutput[66]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[66]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_67_U1 ( .A(RoundKey[67]), .B(
        KeyExpansionOutput[67]), .S(MuxKeyExpansion_n19), .Z(
        RoundKeyOutput[67]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_68_U1 ( .A(RoundKey[68]), .B(
        KeyExpansionOutput[68]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[68]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_69_U1 ( .A(RoundKey[69]), .B(
        KeyExpansionOutput[69]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[69]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_70_U1 ( .A(RoundKey[70]), .B(
        KeyExpansionOutput[70]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[70]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_71_U1 ( .A(RoundKey[71]), .B(
        KeyExpansionOutput[71]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[71]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_72_U1 ( .A(RoundKey[72]), .B(
        KeyExpansionOutput[72]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[72]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_73_U1 ( .A(RoundKey[73]), .B(
        KeyExpansionOutput[73]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[73]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_74_U1 ( .A(RoundKey[74]), .B(
        KeyExpansionOutput[74]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[74]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_75_U1 ( .A(RoundKey[75]), .B(
        KeyExpansionOutput[75]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[75]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_76_U1 ( .A(RoundKey[76]), .B(
        KeyExpansionOutput[76]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[76]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_77_U1 ( .A(RoundKey[77]), .B(
        KeyExpansionOutput[77]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[77]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_78_U1 ( .A(RoundKey[78]), .B(
        KeyExpansionOutput[78]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[78]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_79_U1 ( .A(RoundKey[79]), .B(
        KeyExpansionOutput[79]), .S(MuxKeyExpansion_n18), .Z(
        RoundKeyOutput[79]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_80_U1 ( .A(RoundKey[80]), .B(
        KeyExpansionOutput[80]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[80]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_81_U1 ( .A(RoundKey[81]), .B(
        KeyExpansionOutput[81]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[81]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_82_U1 ( .A(RoundKey[82]), .B(
        KeyExpansionOutput[82]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[82]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_83_U1 ( .A(RoundKey[83]), .B(
        KeyExpansionOutput[83]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[83]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_84_U1 ( .A(RoundKey[84]), .B(
        KeyExpansionOutput[84]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[84]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_85_U1 ( .A(RoundKey[85]), .B(
        KeyExpansionOutput[85]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[85]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_86_U1 ( .A(RoundKey[86]), .B(
        KeyExpansionOutput[86]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[86]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_87_U1 ( .A(RoundKey[87]), .B(
        KeyExpansionOutput[87]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[87]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_88_U1 ( .A(RoundKey[88]), .B(
        KeyExpansionOutput[88]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[88]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_89_U1 ( .A(RoundKey[89]), .B(
        KeyExpansionOutput[89]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[89]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_90_U1 ( .A(RoundKey[90]), .B(
        KeyExpansionOutput[90]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[90]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_91_U1 ( .A(RoundKey[91]), .B(
        KeyExpansionOutput[91]), .S(MuxKeyExpansion_n17), .Z(
        RoundKeyOutput[91]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_92_U1 ( .A(RoundKey[92]), .B(
        KeyExpansionOutput[92]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[92]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_93_U1 ( .A(RoundKey[93]), .B(
        KeyExpansionOutput[93]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[93]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_94_U1 ( .A(RoundKey[94]), .B(
        KeyExpansionOutput[94]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[94]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_95_U1 ( .A(RoundKey[95]), .B(
        KeyExpansionOutput[95]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[95]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_96_U1 ( .A(RoundKey[96]), .B(
        KeyExpansionOutput[96]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[96]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_97_U1 ( .A(RoundKey[97]), .B(
        KeyExpansionOutput[97]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[97]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_98_U1 ( .A(RoundKey[98]), .B(
        KeyExpansionOutput[98]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[98]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_99_U1 ( .A(RoundKey[99]), .B(
        KeyExpansionOutput[99]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[99]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_100_U1 ( .A(RoundKey[100]), .B(
        KeyExpansionOutput[100]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[100]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_101_U1 ( .A(RoundKey[101]), .B(
        KeyExpansionOutput[101]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[101]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_102_U1 ( .A(RoundKey[102]), .B(
        KeyExpansionOutput[102]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[102]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_103_U1 ( .A(RoundKey[103]), .B(
        KeyExpansionOutput[103]), .S(MuxKeyExpansion_n16), .Z(
        RoundKeyOutput[103]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_104_U1 ( .A(RoundKey[104]), .B(
        KeyExpansionOutput[104]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[104]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_105_U1 ( .A(RoundKey[105]), .B(
        KeyExpansionOutput[105]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[105]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_106_U1 ( .A(RoundKey[106]), .B(
        KeyExpansionOutput[106]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[106]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_107_U1 ( .A(RoundKey[107]), .B(
        KeyExpansionOutput[107]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[107]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_108_U1 ( .A(RoundKey[108]), .B(
        KeyExpansionOutput[108]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[108]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_109_U1 ( .A(RoundKey[109]), .B(
        KeyExpansionOutput[109]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[109]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_110_U1 ( .A(RoundKey[110]), .B(
        KeyExpansionOutput[110]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[110]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_111_U1 ( .A(RoundKey[111]), .B(
        KeyExpansionOutput[111]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[111]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_112_U1 ( .A(RoundKey[112]), .B(
        KeyExpansionOutput[112]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[112]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_113_U1 ( .A(RoundKey[113]), .B(
        KeyExpansionOutput[113]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[113]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_114_U1 ( .A(RoundKey[114]), .B(
        KeyExpansionOutput[114]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[114]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_115_U1 ( .A(RoundKey[115]), .B(
        KeyExpansionOutput[115]), .S(MuxKeyExpansion_n15), .Z(
        RoundKeyOutput[115]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_116_U1 ( .A(RoundKey[116]), .B(
        KeyExpansionOutput[116]), .S(MuxKeyExpansion_n14), .Z(
        RoundKeyOutput[116]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_117_U1 ( .A(RoundKey[117]), .B(
        KeyExpansionOutput[117]), .S(MuxKeyExpansion_n14), .Z(
        RoundKeyOutput[117]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_118_U1 ( .A(RoundKey[118]), .B(
        KeyExpansionOutput[118]), .S(MuxKeyExpansion_n14), .Z(
        RoundKeyOutput[118]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_119_U1 ( .A(RoundKey[119]), .B(
        KeyExpansionOutput[119]), .S(MuxKeyExpansion_n14), .Z(
        RoundKeyOutput[119]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_120_U1 ( .A(RoundKey[120]), .B(
        KeyExpansionOutput[120]), .S(MuxKeyExpansion_n14), .Z(
        RoundKeyOutput[120]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_121_U1 ( .A(RoundKey[121]), .B(
        KeyExpansionOutput[121]), .S(MuxKeyExpansion_n14), .Z(
        RoundKeyOutput[121]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_122_U1 ( .A(RoundKey[122]), .B(
        KeyExpansionOutput[122]), .S(MuxKeyExpansion_n14), .Z(
        RoundKeyOutput[122]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_123_U1 ( .A(RoundKey[123]), .B(
        KeyExpansionOutput[123]), .S(MuxKeyExpansion_n14), .Z(
        RoundKeyOutput[123]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_124_U1 ( .A(RoundKey[124]), .B(
        KeyExpansionOutput[124]), .S(MuxKeyExpansion_n14), .Z(
        RoundKeyOutput[124]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_125_U1 ( .A(RoundKey[125]), .B(
        KeyExpansionOutput[125]), .S(MuxKeyExpansion_n14), .Z(
        RoundKeyOutput[125]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_126_U1 ( .A(RoundKey[126]), .B(
        KeyExpansionOutput[126]), .S(MuxKeyExpansion_n14), .Z(
        RoundKeyOutput[126]) );
  MUX2_X1 MuxKeyExpansion_mux_inst_127_U1 ( .A(RoundKey[127]), .B(
        KeyExpansionOutput[127]), .S(MuxKeyExpansion_n14), .Z(
        RoundKeyOutput[127]) );
  NOR2_X1 RoundCounterIns_U11 ( .A1(reset), .A2(RoundCounterIns_n10), .ZN(
        RoundCounterIns_n45) );
  XNOR2_X1 RoundCounterIns_U10 ( .A(RoundCounter[0]), .B(AKSRnotDone), .ZN(
        RoundCounterIns_n10) );
  NOR2_X1 RoundCounterIns_U9 ( .A1(reset), .A2(RoundCounterIns_n9), .ZN(
        RoundCounterIns_n44) );
  XOR2_X1 RoundCounterIns_U8 ( .A(RoundCounter[1]), .B(RoundCounterIns_n8), 
        .Z(RoundCounterIns_n9) );
  NOR2_X1 RoundCounterIns_U7 ( .A1(reset), .A2(RoundCounterIns_n7), .ZN(
        RoundCounterIns_n42) );
  XOR2_X1 RoundCounterIns_U6 ( .A(RoundCounter[3]), .B(RoundCounterIns_n6), 
        .Z(RoundCounterIns_n7) );
  NAND2_X1 RoundCounterIns_U5 ( .A1(RoundCounterIns_n5), .A2(RoundCounter[2]), 
        .ZN(RoundCounterIns_n6) );
  NOR2_X1 RoundCounterIns_U4 ( .A1(reset), .A2(RoundCounterIns_n4), .ZN(
        RoundCounterIns_n1) );
  XNOR2_X1 RoundCounterIns_U3 ( .A(RoundCounter[2]), .B(RoundCounterIns_n5), 
        .ZN(RoundCounterIns_n4) );
  NOR2_X1 RoundCounterIns_U2 ( .A1(RoundCounterIns_n2), .A2(RoundCounterIns_n8), .ZN(RoundCounterIns_n5) );
  NAND2_X1 RoundCounterIns_U1 ( .A1(AKSRnotDone), .A2(RoundCounter[0]), .ZN(
        RoundCounterIns_n8) );
  INV_X1 RoundCounterIns_count_reg_0__U1 ( .A(RoundCounter[0]), .ZN(
        RoundCounterIns_count_reg_0__QN) );
  DFF_X1 RoundCounterIns_count_reg_0__FF_FF ( .D(RoundCounterIns_n45), .CK(clk), .Q(RoundCounter[0]), .QN() );
  INV_X1 RoundCounterIns_count_reg_1__U1 ( .A(RoundCounter[1]), .ZN(
        RoundCounterIns_n2) );
  DFF_X1 RoundCounterIns_count_reg_1__FF_FF ( .D(RoundCounterIns_n44), .CK(clk), .Q(RoundCounter[1]), .QN() );
  INV_X1 RoundCounterIns_count_reg_2__U1 ( .A(RoundCounter[2]), .ZN(
        RoundCounterIns_count_reg_2__QN) );
  DFF_X1 RoundCounterIns_count_reg_2__FF_FF ( .D(RoundCounterIns_n1), .CK(clk), 
        .Q(RoundCounter[2]), .QN() );
  INV_X1 RoundCounterIns_count_reg_3__U1 ( .A(RoundCounter[3]), .ZN(
        RoundCounterIns_count_reg_3__QN) );
  DFF_X1 RoundCounterIns_count_reg_3__FF_FF ( .D(RoundCounterIns_n42), .CK(clk), .Q(RoundCounter[3]), .QN() );
  NOR2_X1 InRoundCounterIns_U13 ( .A1(reset), .A2(InRoundCounterIns_n12), .ZN(
        InRoundCounterIns_n41) );
  XOR2_X1 InRoundCounterIns_U12 ( .A(InRoundCounter[0]), .B(
        InRoundCounterIns_n11), .Z(InRoundCounterIns_n12) );
  NAND2_X1 InRoundCounterIns_U11 ( .A1(InRoundCounterIns_n10), .A2(1'b1), .ZN(
        InRoundCounterIns_n11) );
  NAND2_X1 InRoundCounterIns_U10 ( .A1(InRoundCounterIns_n9), .A2(
        InRoundCounter[2]), .ZN(InRoundCounterIns_n10) );
  NAND2_X1 InRoundCounterIns_U9 ( .A1(InRoundCounter[0]), .A2(
        InRoundCounter[1]), .ZN(InRoundCounterIns_n9) );
  NOR2_X1 InRoundCounterIns_U8 ( .A1(reset), .A2(InRoundCounterIns_n8), .ZN(
        InRoundCounterIns_n40) );
  MUX2_X1 InRoundCounterIns_U7 ( .A(InRoundCounterIns_n7), .B(
        InRoundCounterIns_n5), .S(InRoundCounter[1]), .Z(InRoundCounterIns_n8)
         );
  NOR2_X1 InRoundCounterIns_U6 ( .A1(reset), .A2(InRoundCounterIns_n4), .ZN(
        InRoundCounterIns_n39) );
  NOR2_X1 InRoundCounterIns_U5 ( .A1(InRoundCounterIns_n3), .A2(
        InRoundCounterIns_n2), .ZN(InRoundCounterIns_n4) );
  NOR2_X1 InRoundCounterIns_U4 ( .A1(InRoundCounterIns_n1), .A2(
        InRoundCounterIns_n7), .ZN(InRoundCounterIns_n2) );
  NAND2_X1 InRoundCounterIns_U3 ( .A1(InRoundCounterIns_n5), .A2(
        InRoundCounterIns_n6), .ZN(InRoundCounterIns_n7) );
  AND2_X1 InRoundCounterIns_U2 ( .A1(InRoundCounter[0]), .A2(1'b1), .ZN(
        InRoundCounterIns_n5) );
  NOR2_X1 InRoundCounterIns_U1 ( .A1(1'b1), .A2(InRoundCounterIns_n6), .ZN(
        InRoundCounterIns_n3) );
  INV_X1 InRoundCounterIns_count_reg_0__U1 ( .A(InRoundCounter[0]), .ZN(
        InRoundCounterIns_count_reg_0__QN) );
  DFF_X1 InRoundCounterIns_count_reg_0__FF_FF ( .D(InRoundCounterIns_n41), 
        .CK(clk), .Q(InRoundCounter[0]), .QN() );
  INV_X1 InRoundCounterIns_count_reg_1__U1 ( .A(InRoundCounter[1]), .ZN(
        InRoundCounterIns_n1) );
  DFF_X1 InRoundCounterIns_count_reg_1__FF_FF ( .D(InRoundCounterIns_n40), 
        .CK(clk), .Q(InRoundCounter[1]), .QN() );
  INV_X1 InRoundCounterIns_count_reg_2__U1 ( .A(InRoundCounter[2]), .ZN(
        InRoundCounterIns_n6) );
  DFF_X1 InRoundCounterIns_count_reg_2__FF_FF ( .D(InRoundCounterIns_n39), 
        .CK(clk), .Q(InRoundCounter[2]), .QN() );
endmodule

