/* modified netlist. Source: module AES in file AES.v */
/* clock gating is added to the circuit, the latency increased 2 time(s)  */

module AES_GHPC_ANF_ClockGating_d1 (plaintext_s0, key_s0, clk, reset, plaintext_s1, key_s1, Fresh, ciphertext_s0, done, ciphertext_s1, Synch);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [31:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output Synch ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_416 ;
    wire signal_418 ;
    wire signal_420 ;
    wire signal_422 ;
    wire signal_424 ;
    wire signal_426 ;
    wire signal_428 ;
    wire signal_430 ;
    wire signal_432 ;
    wire signal_434 ;
    wire signal_436 ;
    wire signal_438 ;
    wire signal_440 ;
    wire signal_442 ;
    wire signal_444 ;
    wire signal_446 ;
    wire signal_448 ;
    wire signal_450 ;
    wire signal_452 ;
    wire signal_454 ;
    wire signal_456 ;
    wire signal_458 ;
    wire signal_460 ;
    wire signal_462 ;
    wire signal_464 ;
    wire signal_466 ;
    wire signal_468 ;
    wire signal_470 ;
    wire signal_472 ;
    wire signal_474 ;
    wire signal_476 ;
    wire signal_478 ;
    wire signal_480 ;
    wire signal_482 ;
    wire signal_484 ;
    wire signal_486 ;
    wire signal_488 ;
    wire signal_490 ;
    wire signal_492 ;
    wire signal_494 ;
    wire signal_496 ;
    wire signal_498 ;
    wire signal_500 ;
    wire signal_502 ;
    wire signal_504 ;
    wire signal_506 ;
    wire signal_508 ;
    wire signal_510 ;
    wire signal_512 ;
    wire signal_514 ;
    wire signal_516 ;
    wire signal_518 ;
    wire signal_520 ;
    wire signal_522 ;
    wire signal_524 ;
    wire signal_526 ;
    wire signal_528 ;
    wire signal_530 ;
    wire signal_532 ;
    wire signal_534 ;
    wire signal_536 ;
    wire signal_538 ;
    wire signal_540 ;
    wire signal_542 ;
    wire signal_544 ;
    wire signal_546 ;
    wire signal_548 ;
    wire signal_550 ;
    wire signal_552 ;
    wire signal_554 ;
    wire signal_556 ;
    wire signal_558 ;
    wire signal_560 ;
    wire signal_562 ;
    wire signal_564 ;
    wire signal_566 ;
    wire signal_568 ;
    wire signal_570 ;
    wire signal_572 ;
    wire signal_574 ;
    wire signal_576 ;
    wire signal_578 ;
    wire signal_580 ;
    wire signal_582 ;
    wire signal_584 ;
    wire signal_586 ;
    wire signal_588 ;
    wire signal_590 ;
    wire signal_592 ;
    wire signal_594 ;
    wire signal_596 ;
    wire signal_598 ;
    wire signal_600 ;
    wire signal_602 ;
    wire signal_604 ;
    wire signal_606 ;
    wire signal_608 ;
    wire signal_610 ;
    wire signal_612 ;
    wire signal_614 ;
    wire signal_616 ;
    wire signal_618 ;
    wire signal_620 ;
    wire signal_622 ;
    wire signal_624 ;
    wire signal_626 ;
    wire signal_628 ;
    wire signal_630 ;
    wire signal_632 ;
    wire signal_634 ;
    wire signal_636 ;
    wire signal_638 ;
    wire signal_640 ;
    wire signal_642 ;
    wire signal_644 ;
    wire signal_646 ;
    wire signal_648 ;
    wire signal_650 ;
    wire signal_652 ;
    wire signal_654 ;
    wire signal_656 ;
    wire signal_658 ;
    wire signal_660 ;
    wire signal_662 ;
    wire signal_664 ;
    wire signal_666 ;
    wire signal_668 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_788 ;
    wire signal_908 ;
    wire signal_1028 ;
    wire signal_1148 ;
    wire signal_1153 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1229 ;
    wire signal_1231 ;
    wire signal_1233 ;
    wire signal_1235 ;
    wire signal_1237 ;
    wire signal_1239 ;
    wire signal_1241 ;
    wire signal_1243 ;
    wire signal_1245 ;
    wire signal_1247 ;
    wire signal_1249 ;
    wire signal_1251 ;
    wire signal_1253 ;
    wire signal_1255 ;
    wire signal_1257 ;
    wire signal_1259 ;
    wire signal_1261 ;
    wire signal_1263 ;
    wire signal_1265 ;
    wire signal_1267 ;
    wire signal_1269 ;
    wire signal_1271 ;
    wire signal_1273 ;
    wire signal_1275 ;
    wire signal_1277 ;
    wire signal_1279 ;
    wire signal_1281 ;
    wire signal_1283 ;
    wire signal_1285 ;
    wire signal_1287 ;
    wire signal_1289 ;
    wire signal_1291 ;
    wire signal_1293 ;
    wire signal_1295 ;
    wire signal_1297 ;
    wire signal_1299 ;
    wire signal_1301 ;
    wire signal_1303 ;
    wire signal_1305 ;
    wire signal_1307 ;
    wire signal_1309 ;
    wire signal_1311 ;
    wire signal_1313 ;
    wire signal_1315 ;
    wire signal_1317 ;
    wire signal_1319 ;
    wire signal_1321 ;
    wire signal_1323 ;
    wire signal_1325 ;
    wire signal_1327 ;
    wire signal_1329 ;
    wire signal_1331 ;
    wire signal_1333 ;
    wire signal_1335 ;
    wire signal_1337 ;
    wire signal_1339 ;
    wire signal_1341 ;
    wire signal_1343 ;
    wire signal_1345 ;
    wire signal_1347 ;
    wire signal_1349 ;
    wire signal_1351 ;
    wire signal_1353 ;
    wire signal_1355 ;
    wire signal_1357 ;
    wire signal_1359 ;
    wire signal_1361 ;
    wire signal_1363 ;
    wire signal_1365 ;
    wire signal_1367 ;
    wire signal_1369 ;
    wire signal_1371 ;
    wire signal_1373 ;
    wire signal_1375 ;
    wire signal_1377 ;
    wire signal_1379 ;
    wire signal_1381 ;
    wire signal_1383 ;
    wire signal_1385 ;
    wire signal_1387 ;
    wire signal_1389 ;
    wire signal_1391 ;
    wire signal_1393 ;
    wire signal_1395 ;
    wire signal_1397 ;
    wire signal_1399 ;
    wire signal_1401 ;
    wire signal_1403 ;
    wire signal_1405 ;
    wire signal_1407 ;
    wire signal_1409 ;
    wire signal_1411 ;
    wire signal_1413 ;
    wire signal_1415 ;
    wire signal_1417 ;
    wire signal_1419 ;
    wire signal_1421 ;
    wire signal_1423 ;
    wire signal_1425 ;
    wire signal_1427 ;
    wire signal_1429 ;
    wire signal_1431 ;
    wire signal_1433 ;
    wire signal_1435 ;
    wire signal_1437 ;
    wire signal_1439 ;
    wire signal_1441 ;
    wire signal_1443 ;
    wire signal_1445 ;
    wire signal_1447 ;
    wire signal_1449 ;
    wire signal_1451 ;
    wire signal_1453 ;
    wire signal_1455 ;
    wire signal_1457 ;
    wire signal_1459 ;
    wire signal_1461 ;
    wire signal_1463 ;
    wire signal_1465 ;
    wire signal_1467 ;
    wire signal_1469 ;
    wire signal_1471 ;
    wire signal_1473 ;
    wire signal_1475 ;
    wire signal_1477 ;
    wire signal_1479 ;
    wire signal_1481 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2303 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2851 ;
    wire signal_2853 ;
    wire signal_2855 ;
    wire signal_2857 ;
    wire signal_2859 ;
    wire signal_2861 ;
    wire signal_2863 ;
    wire signal_2865 ;
    wire signal_2867 ;
    wire signal_2869 ;
    wire signal_2871 ;
    wire signal_2873 ;
    wire signal_2875 ;
    wire signal_2877 ;
    wire signal_2879 ;
    wire signal_2881 ;
    wire signal_2883 ;
    wire signal_2885 ;
    wire signal_2887 ;
    wire signal_2889 ;
    wire signal_2891 ;
    wire signal_2893 ;
    wire signal_2895 ;
    wire signal_2897 ;
    wire signal_2899 ;
    wire signal_2901 ;
    wire signal_2903 ;
    wire signal_2905 ;
    wire signal_2907 ;
    wire signal_2909 ;
    wire signal_2911 ;
    wire signal_2913 ;
    wire signal_2915 ;
    wire signal_2917 ;
    wire signal_2919 ;
    wire signal_2921 ;
    wire signal_2923 ;
    wire signal_2925 ;
    wire signal_2927 ;
    wire signal_2929 ;
    wire signal_2931 ;
    wire signal_2933 ;
    wire signal_2935 ;
    wire signal_2937 ;
    wire signal_2939 ;
    wire signal_2941 ;
    wire signal_2943 ;
    wire signal_2945 ;
    wire signal_2947 ;
    wire signal_2949 ;
    wire signal_2951 ;
    wire signal_2953 ;
    wire signal_2955 ;
    wire signal_2957 ;
    wire signal_2959 ;
    wire signal_2961 ;
    wire signal_2963 ;
    wire signal_2965 ;
    wire signal_2967 ;
    wire signal_2969 ;
    wire signal_2971 ;
    wire signal_2973 ;
    wire signal_2975 ;
    wire signal_2977 ;
    wire signal_2979 ;
    wire signal_2981 ;
    wire signal_2983 ;
    wire signal_2985 ;
    wire signal_2987 ;
    wire signal_2989 ;
    wire signal_2991 ;
    wire signal_2993 ;
    wire signal_2995 ;
    wire signal_2997 ;
    wire signal_2999 ;
    wire signal_3001 ;
    wire signal_3003 ;
    wire signal_3005 ;
    wire signal_3007 ;
    wire signal_3009 ;
    wire signal_3011 ;
    wire signal_3013 ;
    wire signal_3015 ;
    wire signal_3017 ;
    wire signal_3019 ;
    wire signal_3021 ;
    wire signal_3023 ;
    wire signal_3025 ;
    wire signal_3027 ;
    wire signal_3029 ;
    wire signal_3031 ;
    wire signal_3033 ;
    wire signal_3035 ;
    wire signal_3037 ;
    wire signal_3039 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_3066 ;
    wire signal_3067 ;
    wire signal_3068 ;
    wire signal_3069 ;
    wire signal_3070 ;
    wire signal_3071 ;
    wire signal_3072 ;
    wire signal_3073 ;
    wire signal_3074 ;
    wire signal_3075 ;
    wire signal_3076 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3263 ;
    wire signal_3265 ;
    wire signal_3267 ;
    wire signal_3269 ;
    wire signal_3271 ;
    wire signal_3273 ;
    wire signal_3275 ;
    wire signal_3277 ;
    wire signal_3279 ;
    wire signal_3281 ;
    wire signal_3283 ;
    wire signal_3285 ;
    wire signal_3287 ;
    wire signal_3289 ;
    wire signal_3291 ;
    wire signal_3293 ;
    wire signal_3295 ;
    wire signal_3297 ;
    wire signal_3299 ;
    wire signal_3301 ;
    wire signal_3303 ;
    wire signal_3305 ;
    wire signal_3307 ;
    wire signal_3309 ;
    wire signal_3311 ;
    wire signal_3313 ;
    wire signal_3315 ;
    wire signal_3317 ;
    wire signal_3319 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3325 ;
    wire signal_3327 ;
    wire signal_3329 ;
    wire signal_3331 ;
    wire signal_3333 ;
    wire signal_3335 ;
    wire signal_3337 ;
    wire signal_3339 ;
    wire signal_3341 ;
    wire signal_3343 ;
    wire signal_3345 ;
    wire signal_3347 ;
    wire signal_3349 ;
    wire signal_3351 ;
    wire signal_3353 ;
    wire signal_3355 ;
    wire signal_3357 ;
    wire signal_3359 ;
    wire signal_3361 ;
    wire signal_3363 ;
    wire signal_3365 ;
    wire signal_3367 ;
    wire signal_3369 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3437 ;
    wire signal_3439 ;
    wire signal_3441 ;
    wire signal_3443 ;
    wire signal_3445 ;
    wire signal_3447 ;
    wire signal_3449 ;
    wire signal_3451 ;
    wire signal_3453 ;
    wire signal_3455 ;
    wire signal_3457 ;
    wire signal_3459 ;
    wire signal_3461 ;
    wire signal_3463 ;
    wire signal_3465 ;
    wire signal_3467 ;
    wire signal_3469 ;
    wire signal_3471 ;
    wire signal_3473 ;
    wire signal_3475 ;
    wire signal_3477 ;
    wire signal_3479 ;
    wire signal_3481 ;
    wire signal_3483 ;
    wire signal_3485 ;
    wire signal_3487 ;
    wire signal_3489 ;
    wire signal_3491 ;
    wire signal_3493 ;
    wire signal_3495 ;
    wire signal_3497 ;
    wire signal_3499 ;
    wire signal_3501 ;
    wire signal_3503 ;
    wire signal_3504 ;
    wire signal_3505 ;
    wire signal_3506 ;
    wire signal_3507 ;
    wire signal_3508 ;
    wire signal_3509 ;
    wire signal_3510 ;
    wire signal_3511 ;
    wire signal_3512 ;
    wire signal_3513 ;
    wire signal_3514 ;
    wire signal_3515 ;
    wire signal_3516 ;
    wire signal_3517 ;
    wire signal_3518 ;
    wire signal_3519 ;
    wire signal_3520 ;
    wire signal_3521 ;
    wire signal_3522 ;
    wire signal_3523 ;
    wire signal_3524 ;
    wire signal_3525 ;
    wire signal_3526 ;
    wire signal_3527 ;
    wire signal_3528 ;
    wire signal_3529 ;
    wire signal_3530 ;
    wire signal_3531 ;
    wire signal_3532 ;
    wire signal_3533 ;
    wire signal_3534 ;
    wire signal_3535 ;
    wire signal_3536 ;
    wire signal_3537 ;
    wire signal_3538 ;
    wire signal_3539 ;
    wire signal_3540 ;
    wire signal_3541 ;
    wire signal_3542 ;
    wire signal_3543 ;
    wire signal_3544 ;
    wire signal_3545 ;
    wire signal_3546 ;
    wire signal_3547 ;
    wire signal_3548 ;
    wire signal_3549 ;
    wire signal_3550 ;
    wire signal_3551 ;
    wire signal_3552 ;
    wire signal_3553 ;
    wire signal_3554 ;
    wire signal_3555 ;
    wire signal_3556 ;
    wire signal_3557 ;
    wire signal_3558 ;
    wire signal_3559 ;
    wire signal_3560 ;
    wire signal_3561 ;
    wire signal_3562 ;
    wire signal_3563 ;
    wire signal_3564 ;
    wire signal_3565 ;
    wire signal_3566 ;
    wire signal_3567 ;
    wire signal_3569 ;
    wire signal_3571 ;
    wire signal_3573 ;
    wire signal_3575 ;
    wire signal_3577 ;
    wire signal_3579 ;
    wire signal_3581 ;
    wire signal_3583 ;
    wire signal_3585 ;
    wire signal_3587 ;
    wire signal_3589 ;
    wire signal_3591 ;
    wire signal_3593 ;
    wire signal_3595 ;
    wire signal_3597 ;
    wire signal_3599 ;
    wire signal_3601 ;
    wire signal_3603 ;
    wire signal_3605 ;
    wire signal_3607 ;
    wire signal_3609 ;
    wire signal_3611 ;
    wire signal_3613 ;
    wire signal_3615 ;
    wire signal_3617 ;
    wire signal_3619 ;
    wire signal_3621 ;
    wire signal_3623 ;
    wire signal_3625 ;
    wire signal_3627 ;
    wire signal_3629 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3673 ;
    wire signal_3675 ;
    wire signal_3677 ;
    wire signal_3679 ;
    wire signal_3681 ;
    wire signal_3683 ;
    wire signal_3685 ;
    wire signal_3687 ;
    wire signal_3689 ;
    wire signal_3691 ;
    wire signal_3693 ;
    wire signal_3695 ;
    wire signal_3697 ;
    wire signal_3699 ;
    wire signal_3701 ;
    wire signal_3703 ;
    wire signal_3705 ;
    wire signal_3707 ;
    wire signal_3709 ;
    wire signal_3711 ;
    wire signal_3713 ;
    wire signal_3715 ;
    wire signal_3717 ;
    wire signal_3719 ;
    wire signal_3721 ;
    wire signal_3723 ;
    wire signal_3725 ;
    wire signal_3727 ;
    wire signal_3729 ;
    wire signal_3731 ;
    wire signal_3733 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3745 ;
    wire signal_3747 ;
    wire signal_3749 ;
    wire signal_3751 ;
    wire signal_3753 ;
    wire signal_3755 ;
    wire signal_3757 ;
    wire signal_3759 ;
    wire signal_3792 ;

    /* cells in depth 0 */
    AND2_X1 cell_0 ( .A1 (signal_396), .A2 (signal_395), .ZN (signal_393) ) ;
    NOR2_X1 cell_1 ( .A1 (signal_411), .A2 (signal_400), .ZN (signal_394) ) ;
    AND2_X1 cell_2 ( .A1 (signal_2273), .A2 (signal_394), .ZN (done) ) ;
    INV_X1 cell_3 ( .A (signal_2270), .ZN (signal_411) ) ;
    NOR2_X1 cell_4 ( .A1 (signal_2276), .A2 (signal_2275), .ZN (signal_396) ) ;
    INV_X1 cell_5 ( .A (signal_2271), .ZN (signal_397) ) ;
    NAND2_X1 cell_6 ( .A1 (signal_2272), .A2 (signal_397), .ZN (signal_400) ) ;
    NOR2_X1 cell_7 ( .A1 (done), .A2 (signal_2274), .ZN (signal_395) ) ;
    INV_X1 cell_8 ( .A (signal_2272), .ZN (signal_406) ) ;
    NAND2_X1 cell_9 ( .A1 (signal_406), .A2 (signal_397), .ZN (signal_398) ) ;
    NOR2_X1 cell_10 ( .A1 (signal_2273), .A2 (signal_398), .ZN (signal_2141) ) ;
    NOR2_X1 cell_11 ( .A1 (signal_2273), .A2 (signal_2270), .ZN (signal_409) ) ;
    NOR2_X1 cell_12 ( .A1 (signal_409), .A2 (signal_398), .ZN (signal_2140) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_2270), .A2 (signal_400), .ZN (signal_399) ) ;
    NOR2_X1 cell_14 ( .A1 (signal_411), .A2 (signal_398), .ZN (signal_405) ) ;
    MUX2_X1 cell_15 ( .S (signal_2273), .A (signal_399), .B (signal_405), .Z (signal_2139) ) ;
    INV_X1 cell_16 ( .A (signal_2273), .ZN (signal_401) ) ;
    NOR2_X1 cell_17 ( .A1 (signal_401), .A2 (signal_400), .ZN (signal_402) ) ;
    MUX2_X1 cell_18 ( .S (signal_2270), .A (signal_402), .B (signal_2141), .Z (signal_2138) ) ;
    NAND2_X1 cell_19 ( .A1 (signal_2271), .A2 (signal_409), .ZN (signal_403) ) ;
    NOR2_X1 cell_20 ( .A1 (signal_2272), .A2 (signal_403), .ZN (signal_404) ) ;
    OR2_X1 cell_21 ( .A1 (signal_405), .A2 (signal_404), .ZN (signal_2137) ) ;
    XNOR2_X1 cell_22 ( .A (signal_2271), .B (signal_2270), .ZN (signal_408) ) ;
    NAND2_X1 cell_23 ( .A1 (signal_2273), .A2 (signal_406), .ZN (signal_407) ) ;
    NOR2_X1 cell_24 ( .A1 (signal_408), .A2 (signal_407), .ZN (signal_2136) ) ;
    INV_X1 cell_25 ( .A (signal_409), .ZN (signal_410) ) ;
    NAND2_X1 cell_26 ( .A1 (signal_2272), .A2 (signal_2271), .ZN (signal_412) ) ;
    NOR2_X1 cell_27 ( .A1 (signal_410), .A2 (signal_412), .ZN (signal_2135) ) ;
    NAND2_X1 cell_28 ( .A1 (signal_2273), .A2 (signal_411), .ZN (signal_413) ) ;
    NOR2_X1 cell_29 ( .A1 (signal_413), .A2 (signal_412), .ZN (signal_2134) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_30 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_2339, signal_1793}), .c ({signal_2340, signal_1681}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_31 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({signal_2342, signal_2065}), .c ({signal_2343, signal_1709}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_32 ( .a ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({signal_2345, signal_2064}), .c ({signal_2346, signal_1708}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_33 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({signal_2348, signal_2063}), .c ({signal_2349, signal_1707}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_34 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({signal_2351, signal_2062}), .c ({signal_2352, signal_1706}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_35 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_2354, signal_2061}), .c ({signal_2355, signal_1737}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_36 ( .a ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({signal_2357, signal_2060}), .c ({signal_2358, signal_1736}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_37 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({signal_2360, signal_2059}), .c ({signal_2361, signal_1735}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_38 ( .a ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({signal_2363, signal_2058}), .c ({signal_2364, signal_1734}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_39 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({signal_2366, signal_2057}), .c ({signal_2367, signal_1733}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_40 ( .a ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({signal_2369, signal_2056}), .c ({signal_2370, signal_1732}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_41 ( .a ({ciphertext_s1[74], ciphertext_s0[74]}), .b ({signal_2372, signal_1799}), .c ({signal_2373, signal_1703}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_42 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({signal_2375, signal_2055}), .c ({signal_2376, signal_1731}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_43 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({signal_2378, signal_2054}), .c ({signal_2379, signal_1730}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_44 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({signal_2381, signal_2053}), .c ({signal_2382, signal_1761}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_45 ( .a ({ciphertext_s1[81], ciphertext_s0[81]}), .b ({signal_2384, signal_2052}), .c ({signal_2385, signal_1760}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_46 ( .a ({ciphertext_s1[82], ciphertext_s0[82]}), .b ({signal_2387, signal_2051}), .c ({signal_2388, signal_1759}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_47 ( .a ({ciphertext_s1[83], ciphertext_s0[83]}), .b ({signal_2390, signal_2050}), .c ({signal_2391, signal_1758}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_48 ( .a ({ciphertext_s1[84], ciphertext_s0[84]}), .b ({signal_2393, signal_2049}), .c ({signal_2394, signal_1757}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_49 ( .a ({ciphertext_s1[85], ciphertext_s0[85]}), .b ({signal_2396, signal_2048}), .c ({signal_2397, signal_1756}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_50 ( .a ({ciphertext_s1[86], ciphertext_s0[86]}), .b ({signal_2399, signal_2047}), .c ({signal_2400, signal_1755}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_51 ( .a ({ciphertext_s1[87], ciphertext_s0[87]}), .b ({signal_2402, signal_2046}), .c ({signal_2403, signal_1754}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_52 ( .a ({ciphertext_s1[75], ciphertext_s0[75]}), .b ({signal_2405, signal_1798}), .c ({signal_2406, signal_1702}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_53 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({signal_2408, signal_2045}), .c ({signal_2409, signal_1657}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_54 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({signal_2411, signal_2044}), .c ({signal_2412, signal_1656}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_55 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({signal_2414, signal_2043}), .c ({signal_2415, signal_1655}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_56 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({signal_2417, signal_2042}), .c ({signal_2418, signal_1654}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_57 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({signal_2420, signal_2041}), .c ({signal_2421, signal_1653}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_58 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({signal_2423, signal_2040}), .c ({signal_2424, signal_1652}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_59 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({signal_2426, signal_2039}), .c ({signal_2427, signal_1651}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_60 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({signal_2429, signal_2038}), .c ({signal_2430, signal_1650}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_61 ( .a ({ciphertext_s1[76], ciphertext_s0[76]}), .b ({signal_2432, signal_1797}), .c ({signal_2433, signal_1701}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_62 ( .a ({ciphertext_s1[77], ciphertext_s0[77]}), .b ({signal_2435, signal_1796}), .c ({signal_2436, signal_1700}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_63 ( .a ({ciphertext_s1[78], ciphertext_s0[78]}), .b ({signal_2438, signal_1795}), .c ({signal_2439, signal_1699}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_64 ( .a ({ciphertext_s1[79], ciphertext_s0[79]}), .b ({signal_2441, signal_1794}), .c ({signal_2442, signal_1698}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_65 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({signal_2444, signal_1809}), .c ({signal_2445, signal_1729}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_66 ( .a ({ciphertext_s1[113], ciphertext_s0[113]}), .b ({signal_2447, signal_1808}), .c ({signal_2448, signal_1728}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_67 ( .a ({ciphertext_s1[114], ciphertext_s0[114]}), .b ({signal_2450, signal_1807}), .c ({signal_2451, signal_1727}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_68 ( .a ({ciphertext_s1[115], ciphertext_s0[115]}), .b ({signal_2453, signal_1806}), .c ({signal_2454, signal_1726}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_69 ( .a ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({signal_2456, signal_1792}), .c ({signal_2457, signal_1680}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_70 ( .a ({ciphertext_s1[116], ciphertext_s0[116]}), .b ({signal_2459, signal_1805}), .c ({signal_2460, signal_1725}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_71 ( .a ({ciphertext_s1[117], ciphertext_s0[117]}), .b ({signal_2462, signal_1804}), .c ({signal_2463, signal_1724}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_72 ( .a ({ciphertext_s1[118], ciphertext_s0[118]}), .b ({signal_2465, signal_1803}), .c ({signal_2466, signal_1723}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_73 ( .a ({ciphertext_s1[119], ciphertext_s0[119]}), .b ({signal_2468, signal_1802}), .c ({signal_2469, signal_1722}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_74 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_2471, signal_1785}), .c ({signal_2472, signal_1753}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_75 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({signal_2474, signal_1784}), .c ({signal_2475, signal_1752}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_76 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({signal_2477, signal_1783}), .c ({signal_2478, signal_1751}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_77 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({signal_2480, signal_1782}), .c ({signal_2481, signal_1750}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_78 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_2483, signal_1781}), .c ({signal_2484, signal_1749}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_79 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({signal_2486, signal_1780}), .c ({signal_2487, signal_1748}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_80 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({signal_2489, signal_1791}), .c ({signal_2490, signal_1679}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_81 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({signal_2492, signal_1779}), .c ({signal_2493, signal_1747}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_82 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({signal_2495, signal_1778}), .c ({signal_2496, signal_1746}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_83 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({signal_2498, signal_2133}), .c ({signal_2499, signal_1777}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_84 ( .a ({ciphertext_s1[65], ciphertext_s0[65]}), .b ({signal_2501, signal_2132}), .c ({signal_2502, signal_1776}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_85 ( .a ({ciphertext_s1[66], ciphertext_s0[66]}), .b ({signal_2504, signal_2131}), .c ({signal_2505, signal_1775}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_86 ( .a ({ciphertext_s1[67], ciphertext_s0[67]}), .b ({signal_2507, signal_2130}), .c ({signal_2508, signal_1774}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_87 ( .a ({ciphertext_s1[68], ciphertext_s0[68]}), .b ({signal_2510, signal_2129}), .c ({signal_2511, signal_1773}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_88 ( .a ({ciphertext_s1[69], ciphertext_s0[69]}), .b ({signal_2513, signal_2128}), .c ({signal_2514, signal_1772}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_89 ( .a ({ciphertext_s1[70], ciphertext_s0[70]}), .b ({signal_2516, signal_2127}), .c ({signal_2517, signal_1771}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_90 ( .a ({ciphertext_s1[71], ciphertext_s0[71]}), .b ({signal_2519, signal_2126}), .c ({signal_2520, signal_1770}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_91 ( .a ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({signal_2522, signal_1790}), .c ({signal_2523, signal_1678}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_92 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({signal_2525, signal_2125}), .c ({signal_2526, signal_1673}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_93 ( .a ({ciphertext_s1[105], ciphertext_s0[105]}), .b ({signal_2528, signal_2124}), .c ({signal_2529, signal_1672}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_94 ( .a ({ciphertext_s1[106], ciphertext_s0[106]}), .b ({signal_2531, signal_2123}), .c ({signal_2532, signal_1671}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_95 ( .a ({ciphertext_s1[107], ciphertext_s0[107]}), .b ({signal_2534, signal_2122}), .c ({signal_2535, signal_1670}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_96 ( .a ({ciphertext_s1[108], ciphertext_s0[108]}), .b ({signal_2537, signal_2121}), .c ({signal_2538, signal_1669}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_97 ( .a ({ciphertext_s1[109], ciphertext_s0[109]}), .b ({signal_2540, signal_2120}), .c ({signal_2541, signal_1668}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_98 ( .a ({ciphertext_s1[110], ciphertext_s0[110]}), .b ({signal_2543, signal_2119}), .c ({signal_2544, signal_1667}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_99 ( .a ({ciphertext_s1[111], ciphertext_s0[111]}), .b ({signal_2546, signal_2118}), .c ({signal_2547, signal_1666}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_100 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_2549, signal_2117}), .c ({signal_2550, signal_1697}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_101 ( .a ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({signal_2552, signal_2116}), .c ({signal_2553, signal_1696}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_102 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({signal_2555, signal_1789}), .c ({signal_2556, signal_1677}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_103 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({signal_2558, signal_2115}), .c ({signal_2559, signal_1695}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_104 ( .a ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({signal_2561, signal_2114}), .c ({signal_2562, signal_1694}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_105 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({signal_2564, signal_2113}), .c ({signal_2565, signal_1693}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_106 ( .a ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({signal_2567, signal_2112}), .c ({signal_2568, signal_1692}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_107 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({signal_2570, signal_2111}), .c ({signal_2571, signal_1691}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_108 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({signal_2573, signal_2110}), .c ({signal_2574, signal_1690}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_109 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_2576, signal_2109}), .c ({signal_2577, signal_1721}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_110 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({signal_2579, signal_2108}), .c ({signal_2580, signal_1720}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_111 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({signal_2582, signal_2107}), .c ({signal_2583, signal_1719}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_112 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({signal_2585, signal_2106}), .c ({signal_2586, signal_1718}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_113 ( .a ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({signal_2588, signal_1788}), .c ({signal_2589, signal_1676}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_114 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_2591, signal_2105}), .c ({signal_2592, signal_1717}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_115 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({signal_2594, signal_2104}), .c ({signal_2595, signal_1716}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_116 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({signal_2597, signal_2103}), .c ({signal_2598, signal_1715}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_117 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({signal_2600, signal_2102}), .c ({signal_2601, signal_1714}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_118 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({signal_2603, signal_2101}), .c ({signal_2604, signal_1745}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_119 ( .a ({ciphertext_s1[97], ciphertext_s0[97]}), .b ({signal_2606, signal_2100}), .c ({signal_2607, signal_1744}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_120 ( .a ({ciphertext_s1[98], ciphertext_s0[98]}), .b ({signal_2609, signal_2099}), .c ({signal_2610, signal_1743}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_121 ( .a ({ciphertext_s1[99], ciphertext_s0[99]}), .b ({signal_2612, signal_2098}), .c ({signal_2613, signal_1742}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_122 ( .a ({ciphertext_s1[100], ciphertext_s0[100]}), .b ({signal_2615, signal_2097}), .c ({signal_2616, signal_1741}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_123 ( .a ({ciphertext_s1[101], ciphertext_s0[101]}), .b ({signal_2618, signal_2096}), .c ({signal_2619, signal_1740}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_124 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({signal_2621, signal_1787}), .c ({signal_2622, signal_1675}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_125 ( .a ({ciphertext_s1[102], ciphertext_s0[102]}), .b ({signal_2624, signal_2095}), .c ({signal_2625, signal_1739}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_126 ( .a ({ciphertext_s1[103], ciphertext_s0[103]}), .b ({signal_2627, signal_2094}), .c ({signal_2628, signal_1738}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_127 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_2630, signal_2093}), .c ({signal_2631, signal_1769}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_128 ( .a ({ciphertext_s1[9], ciphertext_s0[9]}), .b ({signal_2633, signal_2092}), .c ({signal_2634, signal_1768}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_129 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({signal_2636, signal_2091}), .c ({signal_2637, signal_1767}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_130 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({signal_2639, signal_2090}), .c ({signal_2640, signal_1766}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_131 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({signal_2642, signal_2089}), .c ({signal_2643, signal_1765}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_132 ( .a ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({signal_2645, signal_2088}), .c ({signal_2646, signal_1764}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_133 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({signal_2648, signal_2087}), .c ({signal_2649, signal_1763}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_134 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({signal_2651, signal_2086}), .c ({signal_2652, signal_1762}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_135 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({signal_2654, signal_1786}), .c ({signal_2655, signal_1674}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_136 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_2657, signal_2085}), .c ({signal_2658, signal_1665}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_137 ( .a ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({signal_2660, signal_2084}), .c ({signal_2661, signal_1664}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_138 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({signal_2663, signal_2083}), .c ({signal_2664, signal_1663}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_139 ( .a ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({signal_2666, signal_2082}), .c ({signal_2667, signal_1662}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_140 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({signal_2669, signal_2081}), .c ({signal_2670, signal_1661}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_141 ( .a ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({signal_2672, signal_2080}), .c ({signal_2673, signal_1660}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_142 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({signal_2675, signal_2079}), .c ({signal_2676, signal_1659}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_143 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({signal_2678, signal_2078}), .c ({signal_2679, signal_1658}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_144 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({signal_2681, signal_2077}), .c ({signal_2682, signal_1689}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_145 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({signal_2684, signal_2076}), .c ({signal_2685, signal_1688}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_146 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({signal_2687, signal_1801}), .c ({signal_2688, signal_1705}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_147 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({signal_2690, signal_2075}), .c ({signal_2691, signal_1687}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_148 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({signal_2693, signal_2074}), .c ({signal_2694, signal_1686}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_149 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({signal_2696, signal_2073}), .c ({signal_2697, signal_1685}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_150 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({signal_2699, signal_2072}), .c ({signal_2700, signal_1684}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_151 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({signal_2702, signal_2071}), .c ({signal_2703, signal_1683}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_152 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({signal_2705, signal_2070}), .c ({signal_2706, signal_1682}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_153 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_2708, signal_2069}), .c ({signal_2709, signal_1713}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_154 ( .a ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({signal_2711, signal_2068}), .c ({signal_2712, signal_1712}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_155 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({signal_2714, signal_2067}), .c ({signal_2715, signal_1711}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_156 ( .a ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({signal_2717, signal_2066}), .c ({signal_2718, signal_1710}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_157 ( .a ({ciphertext_s1[73], ciphertext_s0[73]}), .b ({signal_2720, signal_1800}), .c ({signal_2721, signal_1704}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_256 ( .s (reset), .b ({signal_2754, signal_1617}), .a ({plaintext_s1[32], plaintext_s0[32]}), .c ({signal_2851, signal_478}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_259 ( .s (reset), .b ({signal_2755, signal_1616}), .a ({plaintext_s1[33], plaintext_s0[33]}), .c ({signal_2853, signal_480}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_262 ( .s (reset), .b ({signal_2756, signal_1615}), .a ({plaintext_s1[34], plaintext_s0[34]}), .c ({signal_2855, signal_482}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_265 ( .s (reset), .b ({signal_2757, signal_1614}), .a ({plaintext_s1[35], plaintext_s0[35]}), .c ({signal_2857, signal_484}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_268 ( .s (reset), .b ({signal_2758, signal_1613}), .a ({plaintext_s1[36], plaintext_s0[36]}), .c ({signal_2859, signal_486}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_271 ( .s (reset), .b ({signal_2759, signal_1612}), .a ({plaintext_s1[37], plaintext_s0[37]}), .c ({signal_2861, signal_488}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_274 ( .s (reset), .b ({signal_2760, signal_1611}), .a ({plaintext_s1[38], plaintext_s0[38]}), .c ({signal_2863, signal_490}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_277 ( .s (reset), .b ({signal_2761, signal_1610}), .a ({plaintext_s1[39], plaintext_s0[39]}), .c ({signal_2865, signal_492}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_280 ( .s (reset), .b ({signal_2762, signal_1609}), .a ({plaintext_s1[40], plaintext_s0[40]}), .c ({signal_2867, signal_494}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_283 ( .s (reset), .b ({signal_2763, signal_1608}), .a ({plaintext_s1[41], plaintext_s0[41]}), .c ({signal_2869, signal_496}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_286 ( .s (reset), .b ({signal_2764, signal_1607}), .a ({plaintext_s1[42], plaintext_s0[42]}), .c ({signal_2871, signal_498}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_289 ( .s (reset), .b ({signal_2765, signal_1606}), .a ({plaintext_s1[43], plaintext_s0[43]}), .c ({signal_2873, signal_500}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_292 ( .s (reset), .b ({signal_2766, signal_1605}), .a ({plaintext_s1[44], plaintext_s0[44]}), .c ({signal_2875, signal_502}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_295 ( .s (reset), .b ({signal_2767, signal_1604}), .a ({plaintext_s1[45], plaintext_s0[45]}), .c ({signal_2877, signal_504}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_298 ( .s (reset), .b ({signal_2768, signal_1603}), .a ({plaintext_s1[46], plaintext_s0[46]}), .c ({signal_2879, signal_506}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_301 ( .s (reset), .b ({signal_2769, signal_1602}), .a ({plaintext_s1[47], plaintext_s0[47]}), .c ({signal_2881, signal_508}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_304 ( .s (reset), .b ({signal_2770, signal_1601}), .a ({plaintext_s1[48], plaintext_s0[48]}), .c ({signal_2883, signal_510}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_307 ( .s (reset), .b ({signal_2771, signal_1600}), .a ({plaintext_s1[49], plaintext_s0[49]}), .c ({signal_2885, signal_512}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_310 ( .s (reset), .b ({signal_2772, signal_1599}), .a ({plaintext_s1[50], plaintext_s0[50]}), .c ({signal_2887, signal_514}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_313 ( .s (reset), .b ({signal_2773, signal_1598}), .a ({plaintext_s1[51], plaintext_s0[51]}), .c ({signal_2889, signal_516}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_316 ( .s (reset), .b ({signal_2774, signal_1597}), .a ({plaintext_s1[52], plaintext_s0[52]}), .c ({signal_2891, signal_518}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_319 ( .s (reset), .b ({signal_2775, signal_1596}), .a ({plaintext_s1[53], plaintext_s0[53]}), .c ({signal_2893, signal_520}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_322 ( .s (reset), .b ({signal_2776, signal_1595}), .a ({plaintext_s1[54], plaintext_s0[54]}), .c ({signal_2895, signal_522}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_325 ( .s (reset), .b ({signal_2777, signal_1594}), .a ({plaintext_s1[55], plaintext_s0[55]}), .c ({signal_2897, signal_524}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_328 ( .s (reset), .b ({signal_2778, signal_1593}), .a ({plaintext_s1[56], plaintext_s0[56]}), .c ({signal_2899, signal_526}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_331 ( .s (reset), .b ({signal_2779, signal_1592}), .a ({plaintext_s1[57], plaintext_s0[57]}), .c ({signal_2901, signal_528}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_334 ( .s (reset), .b ({signal_2780, signal_1591}), .a ({plaintext_s1[58], plaintext_s0[58]}), .c ({signal_2903, signal_530}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_337 ( .s (reset), .b ({signal_2781, signal_1590}), .a ({plaintext_s1[59], plaintext_s0[59]}), .c ({signal_2905, signal_532}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_340 ( .s (reset), .b ({signal_2782, signal_1589}), .a ({plaintext_s1[60], plaintext_s0[60]}), .c ({signal_2907, signal_534}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_343 ( .s (reset), .b ({signal_2783, signal_1588}), .a ({plaintext_s1[61], plaintext_s0[61]}), .c ({signal_2909, signal_536}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_346 ( .s (reset), .b ({signal_2784, signal_1587}), .a ({plaintext_s1[62], plaintext_s0[62]}), .c ({signal_2911, signal_538}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_349 ( .s (reset), .b ({signal_2785, signal_1586}), .a ({plaintext_s1[63], plaintext_s0[63]}), .c ({signal_2913, signal_540}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_352 ( .s (reset), .b ({signal_2786, signal_1585}), .a ({plaintext_s1[64], plaintext_s0[64]}), .c ({signal_2915, signal_542}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_355 ( .s (reset), .b ({signal_2787, signal_1584}), .a ({plaintext_s1[65], plaintext_s0[65]}), .c ({signal_2917, signal_544}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_358 ( .s (reset), .b ({signal_2788, signal_1583}), .a ({plaintext_s1[66], plaintext_s0[66]}), .c ({signal_2919, signal_546}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_361 ( .s (reset), .b ({signal_2789, signal_1582}), .a ({plaintext_s1[67], plaintext_s0[67]}), .c ({signal_2921, signal_548}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_364 ( .s (reset), .b ({signal_2790, signal_1581}), .a ({plaintext_s1[68], plaintext_s0[68]}), .c ({signal_2923, signal_550}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_367 ( .s (reset), .b ({signal_2791, signal_1580}), .a ({plaintext_s1[69], plaintext_s0[69]}), .c ({signal_2925, signal_552}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_370 ( .s (reset), .b ({signal_2792, signal_1579}), .a ({plaintext_s1[70], plaintext_s0[70]}), .c ({signal_2927, signal_554}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_373 ( .s (reset), .b ({signal_2793, signal_1578}), .a ({plaintext_s1[71], plaintext_s0[71]}), .c ({signal_2929, signal_556}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_376 ( .s (reset), .b ({signal_2794, signal_1577}), .a ({plaintext_s1[72], plaintext_s0[72]}), .c ({signal_2931, signal_558}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_379 ( .s (reset), .b ({signal_2795, signal_1576}), .a ({plaintext_s1[73], plaintext_s0[73]}), .c ({signal_2933, signal_560}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_382 ( .s (reset), .b ({signal_2796, signal_1575}), .a ({plaintext_s1[74], plaintext_s0[74]}), .c ({signal_2935, signal_562}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_385 ( .s (reset), .b ({signal_2797, signal_1574}), .a ({plaintext_s1[75], plaintext_s0[75]}), .c ({signal_2937, signal_564}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_388 ( .s (reset), .b ({signal_2798, signal_1573}), .a ({plaintext_s1[76], plaintext_s0[76]}), .c ({signal_2939, signal_566}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_391 ( .s (reset), .b ({signal_2799, signal_1572}), .a ({plaintext_s1[77], plaintext_s0[77]}), .c ({signal_2941, signal_568}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_394 ( .s (reset), .b ({signal_2800, signal_1571}), .a ({plaintext_s1[78], plaintext_s0[78]}), .c ({signal_2943, signal_570}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_397 ( .s (reset), .b ({signal_2801, signal_1570}), .a ({plaintext_s1[79], plaintext_s0[79]}), .c ({signal_2945, signal_572}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_400 ( .s (reset), .b ({signal_2802, signal_1569}), .a ({plaintext_s1[80], plaintext_s0[80]}), .c ({signal_2947, signal_574}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_403 ( .s (reset), .b ({signal_2803, signal_1568}), .a ({plaintext_s1[81], plaintext_s0[81]}), .c ({signal_2949, signal_576}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_406 ( .s (reset), .b ({signal_2804, signal_1567}), .a ({plaintext_s1[82], plaintext_s0[82]}), .c ({signal_2951, signal_578}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_409 ( .s (reset), .b ({signal_2805, signal_1566}), .a ({plaintext_s1[83], plaintext_s0[83]}), .c ({signal_2953, signal_580}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_412 ( .s (reset), .b ({signal_2806, signal_1565}), .a ({plaintext_s1[84], plaintext_s0[84]}), .c ({signal_2955, signal_582}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_415 ( .s (reset), .b ({signal_2807, signal_1564}), .a ({plaintext_s1[85], plaintext_s0[85]}), .c ({signal_2957, signal_584}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_418 ( .s (reset), .b ({signal_2808, signal_1563}), .a ({plaintext_s1[86], plaintext_s0[86]}), .c ({signal_2959, signal_586}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_421 ( .s (reset), .b ({signal_2809, signal_1562}), .a ({plaintext_s1[87], plaintext_s0[87]}), .c ({signal_2961, signal_588}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_424 ( .s (reset), .b ({signal_2810, signal_1561}), .a ({plaintext_s1[88], plaintext_s0[88]}), .c ({signal_2963, signal_590}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_427 ( .s (reset), .b ({signal_2811, signal_1560}), .a ({plaintext_s1[89], plaintext_s0[89]}), .c ({signal_2965, signal_592}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_430 ( .s (reset), .b ({signal_2812, signal_1559}), .a ({plaintext_s1[90], plaintext_s0[90]}), .c ({signal_2967, signal_594}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_433 ( .s (reset), .b ({signal_2813, signal_1558}), .a ({plaintext_s1[91], plaintext_s0[91]}), .c ({signal_2969, signal_596}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_436 ( .s (reset), .b ({signal_2814, signal_1557}), .a ({plaintext_s1[92], plaintext_s0[92]}), .c ({signal_2971, signal_598}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_439 ( .s (reset), .b ({signal_2815, signal_1556}), .a ({plaintext_s1[93], plaintext_s0[93]}), .c ({signal_2973, signal_600}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_442 ( .s (reset), .b ({signal_2816, signal_1555}), .a ({plaintext_s1[94], plaintext_s0[94]}), .c ({signal_2975, signal_602}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_445 ( .s (reset), .b ({signal_2817, signal_1554}), .a ({plaintext_s1[95], plaintext_s0[95]}), .c ({signal_2977, signal_604}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_448 ( .s (reset), .b ({signal_2818, signal_1553}), .a ({plaintext_s1[96], plaintext_s0[96]}), .c ({signal_2979, signal_606}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_451 ( .s (reset), .b ({signal_2819, signal_1552}), .a ({plaintext_s1[97], plaintext_s0[97]}), .c ({signal_2981, signal_608}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_454 ( .s (reset), .b ({signal_2820, signal_1551}), .a ({plaintext_s1[98], plaintext_s0[98]}), .c ({signal_2983, signal_610}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_457 ( .s (reset), .b ({signal_2821, signal_1550}), .a ({plaintext_s1[99], plaintext_s0[99]}), .c ({signal_2985, signal_612}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_460 ( .s (reset), .b ({signal_2822, signal_1549}), .a ({plaintext_s1[100], plaintext_s0[100]}), .c ({signal_2987, signal_614}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_463 ( .s (reset), .b ({signal_2823, signal_1548}), .a ({plaintext_s1[101], plaintext_s0[101]}), .c ({signal_2989, signal_616}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_466 ( .s (reset), .b ({signal_2824, signal_1547}), .a ({plaintext_s1[102], plaintext_s0[102]}), .c ({signal_2991, signal_618}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_469 ( .s (reset), .b ({signal_2825, signal_1546}), .a ({plaintext_s1[103], plaintext_s0[103]}), .c ({signal_2993, signal_620}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_472 ( .s (reset), .b ({signal_2826, signal_1545}), .a ({plaintext_s1[104], plaintext_s0[104]}), .c ({signal_2995, signal_622}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_475 ( .s (reset), .b ({signal_2827, signal_1544}), .a ({plaintext_s1[105], plaintext_s0[105]}), .c ({signal_2997, signal_624}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_478 ( .s (reset), .b ({signal_2828, signal_1543}), .a ({plaintext_s1[106], plaintext_s0[106]}), .c ({signal_2999, signal_626}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_481 ( .s (reset), .b ({signal_2829, signal_1542}), .a ({plaintext_s1[107], plaintext_s0[107]}), .c ({signal_3001, signal_628}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_484 ( .s (reset), .b ({signal_2830, signal_1541}), .a ({plaintext_s1[108], plaintext_s0[108]}), .c ({signal_3003, signal_630}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_487 ( .s (reset), .b ({signal_2831, signal_1540}), .a ({plaintext_s1[109], plaintext_s0[109]}), .c ({signal_3005, signal_632}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_490 ( .s (reset), .b ({signal_2832, signal_1539}), .a ({plaintext_s1[110], plaintext_s0[110]}), .c ({signal_3007, signal_634}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_493 ( .s (reset), .b ({signal_2833, signal_1538}), .a ({plaintext_s1[111], plaintext_s0[111]}), .c ({signal_3009, signal_636}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_496 ( .s (reset), .b ({signal_2834, signal_1537}), .a ({plaintext_s1[112], plaintext_s0[112]}), .c ({signal_3011, signal_638}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_499 ( .s (reset), .b ({signal_2835, signal_1536}), .a ({plaintext_s1[113], plaintext_s0[113]}), .c ({signal_3013, signal_640}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_502 ( .s (reset), .b ({signal_2836, signal_1535}), .a ({plaintext_s1[114], plaintext_s0[114]}), .c ({signal_3015, signal_642}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_505 ( .s (reset), .b ({signal_2837, signal_1534}), .a ({plaintext_s1[115], plaintext_s0[115]}), .c ({signal_3017, signal_644}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_508 ( .s (reset), .b ({signal_2838, signal_1533}), .a ({plaintext_s1[116], plaintext_s0[116]}), .c ({signal_3019, signal_646}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_511 ( .s (reset), .b ({signal_2839, signal_1532}), .a ({plaintext_s1[117], plaintext_s0[117]}), .c ({signal_3021, signal_648}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_514 ( .s (reset), .b ({signal_2840, signal_1531}), .a ({plaintext_s1[118], plaintext_s0[118]}), .c ({signal_3023, signal_650}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_517 ( .s (reset), .b ({signal_2841, signal_1530}), .a ({plaintext_s1[119], plaintext_s0[119]}), .c ({signal_3025, signal_652}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_520 ( .s (reset), .b ({signal_2842, signal_1529}), .a ({plaintext_s1[120], plaintext_s0[120]}), .c ({signal_3027, signal_654}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_523 ( .s (reset), .b ({signal_2843, signal_1528}), .a ({plaintext_s1[121], plaintext_s0[121]}), .c ({signal_3029, signal_656}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_526 ( .s (reset), .b ({signal_2844, signal_1527}), .a ({plaintext_s1[122], plaintext_s0[122]}), .c ({signal_3031, signal_658}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_529 ( .s (reset), .b ({signal_2845, signal_1526}), .a ({plaintext_s1[123], plaintext_s0[123]}), .c ({signal_3033, signal_660}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_532 ( .s (reset), .b ({signal_2846, signal_1525}), .a ({plaintext_s1[124], plaintext_s0[124]}), .c ({signal_3035, signal_662}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_535 ( .s (reset), .b ({signal_2847, signal_1524}), .a ({plaintext_s1[125], plaintext_s0[125]}), .c ({signal_3037, signal_664}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_538 ( .s (reset), .b ({signal_2848, signal_1523}), .a ({plaintext_s1[126], plaintext_s0[126]}), .c ({signal_3039, signal_666}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_541 ( .s (reset), .b ({signal_2849, signal_1522}), .a ({plaintext_s1[127], plaintext_s0[127]}), .c ({signal_3041, signal_668}) ) ;
    INV_X1 cell_542 ( .A (signal_393), .ZN (signal_670) ) ;
    INV_X1 cell_543 ( .A (signal_670), .ZN (signal_672) ) ;
    INV_X1 cell_544 ( .A (signal_670), .ZN (signal_671) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_545 ( .s (signal_671), .b ({ciphertext_s1[0], ciphertext_s0[0]}), .a ({signal_2444, signal_1809}), .c ({signal_2723, signal_1841}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_546 ( .s (signal_671), .b ({ciphertext_s1[1], ciphertext_s0[1]}), .a ({signal_2447, signal_1808}), .c ({signal_2724, signal_1840}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_547 ( .s (signal_671), .b ({ciphertext_s1[2], ciphertext_s0[2]}), .a ({signal_2450, signal_1807}), .c ({signal_2725, signal_1839}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_548 ( .s (signal_671), .b ({ciphertext_s1[3], ciphertext_s0[3]}), .a ({signal_2453, signal_1806}), .c ({signal_2726, signal_1838}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_549 ( .s (signal_671), .b ({ciphertext_s1[4], ciphertext_s0[4]}), .a ({signal_2459, signal_1805}), .c ({signal_2727, signal_1837}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_550 ( .s (signal_671), .b ({ciphertext_s1[5], ciphertext_s0[5]}), .a ({signal_2462, signal_1804}), .c ({signal_2728, signal_1836}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_551 ( .s (signal_671), .b ({ciphertext_s1[6], ciphertext_s0[6]}), .a ({signal_2465, signal_1803}), .c ({signal_2729, signal_1835}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_552 ( .s (signal_671), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .a ({signal_2468, signal_1802}), .c ({signal_2730, signal_1834}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_553 ( .s (signal_393), .b ({ciphertext_s1[40], ciphertext_s0[40]}), .a ({signal_2687, signal_1801}), .c ({signal_2722, signal_1833}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_554 ( .s (signal_672), .b ({ciphertext_s1[41], ciphertext_s0[41]}), .a ({signal_2720, signal_1800}), .c ({signal_2731, signal_1832}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_555 ( .s (signal_672), .b ({ciphertext_s1[42], ciphertext_s0[42]}), .a ({signal_2372, signal_1799}), .c ({signal_2732, signal_1831}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_556 ( .s (signal_672), .b ({ciphertext_s1[43], ciphertext_s0[43]}), .a ({signal_2405, signal_1798}), .c ({signal_2733, signal_1830}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_557 ( .s (signal_672), .b ({ciphertext_s1[44], ciphertext_s0[44]}), .a ({signal_2432, signal_1797}), .c ({signal_2734, signal_1829}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_558 ( .s (signal_671), .b ({ciphertext_s1[45], ciphertext_s0[45]}), .a ({signal_2435, signal_1796}), .c ({signal_2735, signal_1828}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_559 ( .s (signal_671), .b ({ciphertext_s1[46], ciphertext_s0[46]}), .a ({signal_2438, signal_1795}), .c ({signal_2736, signal_1827}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_560 ( .s (signal_672), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .a ({signal_2441, signal_1794}), .c ({signal_2737, signal_1826}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_561 ( .s (signal_671), .b ({ciphertext_s1[80], ciphertext_s0[80]}), .a ({signal_2339, signal_1793}), .c ({signal_2738, signal_1825}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_562 ( .s (signal_672), .b ({ciphertext_s1[81], ciphertext_s0[81]}), .a ({signal_2456, signal_1792}), .c ({signal_2739, signal_1824}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_563 ( .s (signal_672), .b ({ciphertext_s1[82], ciphertext_s0[82]}), .a ({signal_2489, signal_1791}), .c ({signal_2740, signal_1823}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_564 ( .s (signal_672), .b ({ciphertext_s1[83], ciphertext_s0[83]}), .a ({signal_2522, signal_1790}), .c ({signal_2741, signal_1822}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_565 ( .s (signal_672), .b ({ciphertext_s1[84], ciphertext_s0[84]}), .a ({signal_2555, signal_1789}), .c ({signal_2742, signal_1821}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_566 ( .s (signal_672), .b ({ciphertext_s1[85], ciphertext_s0[85]}), .a ({signal_2588, signal_1788}), .c ({signal_2743, signal_1820}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_567 ( .s (signal_672), .b ({ciphertext_s1[86], ciphertext_s0[86]}), .a ({signal_2621, signal_1787}), .c ({signal_2744, signal_1819}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_568 ( .s (signal_672), .b ({ciphertext_s1[87], ciphertext_s0[87]}), .a ({signal_2654, signal_1786}), .c ({signal_2745, signal_1818}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_569 ( .s (signal_672), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .a ({signal_2471, signal_1785}), .c ({signal_2746, signal_1817}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_570 ( .s (signal_672), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .a ({signal_2474, signal_1784}), .c ({signal_2747, signal_1816}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_571 ( .s (signal_672), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .a ({signal_2477, signal_1783}), .c ({signal_2748, signal_1815}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_572 ( .s (signal_672), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .a ({signal_2480, signal_1782}), .c ({signal_2749, signal_1814}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_573 ( .s (signal_672), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .a ({signal_2483, signal_1781}), .c ({signal_2750, signal_1813}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_574 ( .s (signal_672), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .a ({signal_2486, signal_1780}), .c ({signal_2751, signal_1812}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_575 ( .s (signal_672), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .a ({signal_2492, signal_1779}), .c ({signal_2752, signal_1811}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_576 ( .s (signal_672), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .a ({signal_2495, signal_1778}), .c ({signal_2753, signal_1810}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_581 ( .a ({signal_2726, signal_1838}), .b ({signal_2724, signal_1840}), .c ({signal_3042, signal_788}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_709 ( .a ({signal_2733, signal_1830}), .b ({signal_2731, signal_1832}), .c ({signal_3043, signal_908}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_837 ( .a ({signal_2741, signal_1822}), .b ({signal_2739, signal_1824}), .c ({signal_3044, signal_1028}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_965 ( .a ({signal_2749, signal_1814}), .b ({signal_2747, signal_1816}), .c ({signal_3045, signal_1148}) ) ;
    INV_X1 cell_1197 ( .A (signal_394), .ZN (signal_1217) ) ;
    INV_X1 cell_1198 ( .A (signal_1217), .ZN (signal_1218) ) ;
    INV_X1 cell_1199 ( .A (signal_1217), .ZN (signal_1219) ) ;
    INV_X1 cell_1232 ( .A (signal_393), .ZN (signal_1220) ) ;
    INV_X1 cell_1233 ( .A (signal_1220), .ZN (signal_1223) ) ;
    INV_X1 cell_1234 ( .A (signal_1220), .ZN (signal_1225) ) ;
    INV_X1 cell_1235 ( .A (signal_1220), .ZN (signal_1226) ) ;
    INV_X1 cell_1236 ( .A (signal_1220), .ZN (signal_1224) ) ;
    INV_X1 cell_1237 ( .A (signal_1220), .ZN (signal_1221) ) ;
    INV_X1 cell_1238 ( .A (signal_1220), .ZN (signal_1222) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1271 ( .s (signal_1221), .b ({ciphertext_s1[32], ciphertext_s0[32]}), .a ({signal_2604, signal_1745}), .c ({signal_2754, signal_1617}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1272 ( .s (signal_1222), .b ({ciphertext_s1[33], ciphertext_s0[33]}), .a ({signal_2607, signal_1744}), .c ({signal_2755, signal_1616}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1273 ( .s (signal_1226), .b ({ciphertext_s1[34], ciphertext_s0[34]}), .a ({signal_2610, signal_1743}), .c ({signal_2756, signal_1615}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1274 ( .s (signal_1225), .b ({ciphertext_s1[35], ciphertext_s0[35]}), .a ({signal_2613, signal_1742}), .c ({signal_2757, signal_1614}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1275 ( .s (signal_1224), .b ({ciphertext_s1[36], ciphertext_s0[36]}), .a ({signal_2616, signal_1741}), .c ({signal_2758, signal_1613}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1276 ( .s (signal_1223), .b ({ciphertext_s1[37], ciphertext_s0[37]}), .a ({signal_2619, signal_1740}), .c ({signal_2759, signal_1612}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1277 ( .s (signal_1222), .b ({ciphertext_s1[38], ciphertext_s0[38]}), .a ({signal_2625, signal_1739}), .c ({signal_2760, signal_1611}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1278 ( .s (signal_1221), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .a ({signal_2628, signal_1738}), .c ({signal_2761, signal_1610}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1279 ( .s (signal_1221), .b ({ciphertext_s1[72], ciphertext_s0[72]}), .a ({signal_2355, signal_1737}), .c ({signal_2762, signal_1609}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1280 ( .s (signal_1226), .b ({ciphertext_s1[73], ciphertext_s0[73]}), .a ({signal_2358, signal_1736}), .c ({signal_2763, signal_1608}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1281 ( .s (signal_1225), .b ({ciphertext_s1[74], ciphertext_s0[74]}), .a ({signal_2361, signal_1735}), .c ({signal_2764, signal_1607}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1282 ( .s (signal_1224), .b ({ciphertext_s1[75], ciphertext_s0[75]}), .a ({signal_2364, signal_1734}), .c ({signal_2765, signal_1606}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1283 ( .s (signal_1226), .b ({ciphertext_s1[76], ciphertext_s0[76]}), .a ({signal_2367, signal_1733}), .c ({signal_2766, signal_1605}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1284 ( .s (signal_1225), .b ({ciphertext_s1[77], ciphertext_s0[77]}), .a ({signal_2370, signal_1732}), .c ({signal_2767, signal_1604}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1285 ( .s (signal_1224), .b ({ciphertext_s1[78], ciphertext_s0[78]}), .a ({signal_2376, signal_1731}), .c ({signal_2768, signal_1603}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1286 ( .s (signal_1223), .b ({ciphertext_s1[79], ciphertext_s0[79]}), .a ({signal_2379, signal_1730}), .c ({signal_2769, signal_1602}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1287 ( .s (signal_1222), .b ({ciphertext_s1[112], ciphertext_s0[112]}), .a ({signal_2445, signal_1729}), .c ({signal_2770, signal_1601}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1288 ( .s (signal_1221), .b ({ciphertext_s1[113], ciphertext_s0[113]}), .a ({signal_2448, signal_1728}), .c ({signal_2771, signal_1600}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1289 ( .s (signal_1226), .b ({ciphertext_s1[114], ciphertext_s0[114]}), .a ({signal_2451, signal_1727}), .c ({signal_2772, signal_1599}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1290 ( .s (signal_1225), .b ({ciphertext_s1[115], ciphertext_s0[115]}), .a ({signal_2454, signal_1726}), .c ({signal_2773, signal_1598}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1291 ( .s (signal_1224), .b ({ciphertext_s1[116], ciphertext_s0[116]}), .a ({signal_2460, signal_1725}), .c ({signal_2774, signal_1597}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1292 ( .s (signal_1223), .b ({ciphertext_s1[117], ciphertext_s0[117]}), .a ({signal_2463, signal_1724}), .c ({signal_2775, signal_1596}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1293 ( .s (signal_1222), .b ({ciphertext_s1[118], ciphertext_s0[118]}), .a ({signal_2466, signal_1723}), .c ({signal_2776, signal_1595}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1294 ( .s (signal_1221), .b ({ciphertext_s1[119], ciphertext_s0[119]}), .a ({signal_2469, signal_1722}), .c ({signal_2777, signal_1594}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1295 ( .s (signal_1221), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .a ({signal_2577, signal_1721}), .c ({signal_2778, signal_1593}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1296 ( .s (signal_1221), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .a ({signal_2580, signal_1720}), .c ({signal_2779, signal_1592}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1297 ( .s (signal_1221), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .a ({signal_2583, signal_1719}), .c ({signal_2780, signal_1591}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1298 ( .s (signal_1221), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .a ({signal_2586, signal_1718}), .c ({signal_2781, signal_1590}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1299 ( .s (signal_1221), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .a ({signal_2592, signal_1717}), .c ({signal_2782, signal_1589}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1300 ( .s (signal_1221), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .a ({signal_2595, signal_1716}), .c ({signal_2783, signal_1588}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1301 ( .s (signal_1221), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .a ({signal_2598, signal_1715}), .c ({signal_2784, signal_1587}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1302 ( .s (signal_1221), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .a ({signal_2601, signal_1714}), .c ({signal_2785, signal_1586}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1303 ( .s (signal_1221), .b ({ciphertext_s1[64], ciphertext_s0[64]}), .a ({signal_2709, signal_1713}), .c ({signal_2786, signal_1585}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1304 ( .s (signal_1221), .b ({ciphertext_s1[65], ciphertext_s0[65]}), .a ({signal_2712, signal_1712}), .c ({signal_2787, signal_1584}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1305 ( .s (signal_1221), .b ({ciphertext_s1[66], ciphertext_s0[66]}), .a ({signal_2715, signal_1711}), .c ({signal_2788, signal_1583}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1306 ( .s (signal_1221), .b ({ciphertext_s1[67], ciphertext_s0[67]}), .a ({signal_2718, signal_1710}), .c ({signal_2789, signal_1582}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1307 ( .s (signal_1222), .b ({ciphertext_s1[68], ciphertext_s0[68]}), .a ({signal_2343, signal_1709}), .c ({signal_2790, signal_1581}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1308 ( .s (signal_1222), .b ({ciphertext_s1[69], ciphertext_s0[69]}), .a ({signal_2346, signal_1708}), .c ({signal_2791, signal_1580}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1309 ( .s (signal_1222), .b ({ciphertext_s1[70], ciphertext_s0[70]}), .a ({signal_2349, signal_1707}), .c ({signal_2792, signal_1579}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1310 ( .s (signal_1222), .b ({ciphertext_s1[71], ciphertext_s0[71]}), .a ({signal_2352, signal_1706}), .c ({signal_2793, signal_1578}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1311 ( .s (signal_1222), .b ({ciphertext_s1[104], ciphertext_s0[104]}), .a ({signal_2688, signal_1705}), .c ({signal_2794, signal_1577}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1312 ( .s (signal_1222), .b ({ciphertext_s1[105], ciphertext_s0[105]}), .a ({signal_2721, signal_1704}), .c ({signal_2795, signal_1576}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1313 ( .s (signal_1222), .b ({ciphertext_s1[106], ciphertext_s0[106]}), .a ({signal_2373, signal_1703}), .c ({signal_2796, signal_1575}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1314 ( .s (signal_1222), .b ({ciphertext_s1[107], ciphertext_s0[107]}), .a ({signal_2406, signal_1702}), .c ({signal_2797, signal_1574}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1315 ( .s (signal_1222), .b ({ciphertext_s1[108], ciphertext_s0[108]}), .a ({signal_2433, signal_1701}), .c ({signal_2798, signal_1573}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1316 ( .s (signal_1222), .b ({ciphertext_s1[109], ciphertext_s0[109]}), .a ({signal_2436, signal_1700}), .c ({signal_2799, signal_1572}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1317 ( .s (signal_1222), .b ({ciphertext_s1[110], ciphertext_s0[110]}), .a ({signal_2439, signal_1699}), .c ({signal_2800, signal_1571}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1318 ( .s (signal_1222), .b ({ciphertext_s1[111], ciphertext_s0[111]}), .a ({signal_2442, signal_1698}), .c ({signal_2801, signal_1570}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1319 ( .s (signal_1223), .b ({ciphertext_s1[16], ciphertext_s0[16]}), .a ({signal_2550, signal_1697}), .c ({signal_2802, signal_1569}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1320 ( .s (signal_1223), .b ({ciphertext_s1[17], ciphertext_s0[17]}), .a ({signal_2553, signal_1696}), .c ({signal_2803, signal_1568}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1321 ( .s (signal_1223), .b ({ciphertext_s1[18], ciphertext_s0[18]}), .a ({signal_2559, signal_1695}), .c ({signal_2804, signal_1567}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1322 ( .s (signal_1223), .b ({ciphertext_s1[19], ciphertext_s0[19]}), .a ({signal_2562, signal_1694}), .c ({signal_2805, signal_1566}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1323 ( .s (signal_1223), .b ({ciphertext_s1[20], ciphertext_s0[20]}), .a ({signal_2565, signal_1693}), .c ({signal_2806, signal_1565}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1324 ( .s (signal_1223), .b ({ciphertext_s1[21], ciphertext_s0[21]}), .a ({signal_2568, signal_1692}), .c ({signal_2807, signal_1564}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1325 ( .s (signal_1223), .b ({ciphertext_s1[22], ciphertext_s0[22]}), .a ({signal_2571, signal_1691}), .c ({signal_2808, signal_1563}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1326 ( .s (signal_1223), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .a ({signal_2574, signal_1690}), .c ({signal_2809, signal_1562}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1327 ( .s (signal_1223), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .a ({signal_2682, signal_1689}), .c ({signal_2810, signal_1561}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1328 ( .s (signal_1223), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .a ({signal_2685, signal_1688}), .c ({signal_2811, signal_1560}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1329 ( .s (signal_1223), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .a ({signal_2691, signal_1687}), .c ({signal_2812, signal_1559}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1330 ( .s (signal_1223), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .a ({signal_2694, signal_1686}), .c ({signal_2813, signal_1558}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1331 ( .s (signal_1224), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .a ({signal_2697, signal_1685}), .c ({signal_2814, signal_1557}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1332 ( .s (signal_1224), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .a ({signal_2700, signal_1684}), .c ({signal_2815, signal_1556}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1333 ( .s (signal_1224), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .a ({signal_2703, signal_1683}), .c ({signal_2816, signal_1555}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1334 ( .s (signal_1224), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .a ({signal_2706, signal_1682}), .c ({signal_2817, signal_1554}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1335 ( .s (signal_1224), .b ({ciphertext_s1[96], ciphertext_s0[96]}), .a ({signal_2340, signal_1681}), .c ({signal_2818, signal_1553}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1336 ( .s (signal_1224), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .a ({signal_2457, signal_1680}), .c ({signal_2819, signal_1552}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1337 ( .s (signal_1224), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .a ({signal_2490, signal_1679}), .c ({signal_2820, signal_1551}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1338 ( .s (signal_1224), .b ({ciphertext_s1[99], ciphertext_s0[99]}), .a ({signal_2523, signal_1678}), .c ({signal_2821, signal_1550}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1339 ( .s (signal_1224), .b ({ciphertext_s1[100], ciphertext_s0[100]}), .a ({signal_2556, signal_1677}), .c ({signal_2822, signal_1549}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1340 ( .s (signal_1224), .b ({ciphertext_s1[101], ciphertext_s0[101]}), .a ({signal_2589, signal_1676}), .c ({signal_2823, signal_1548}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1341 ( .s (signal_1224), .b ({ciphertext_s1[102], ciphertext_s0[102]}), .a ({signal_2622, signal_1675}), .c ({signal_2824, signal_1547}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1342 ( .s (signal_1224), .b ({ciphertext_s1[103], ciphertext_s0[103]}), .a ({signal_2655, signal_1674}), .c ({signal_2825, signal_1546}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1343 ( .s (signal_1225), .b ({ciphertext_s1[8], ciphertext_s0[8]}), .a ({signal_2526, signal_1673}), .c ({signal_2826, signal_1545}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1344 ( .s (signal_1225), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .a ({signal_2529, signal_1672}), .c ({signal_2827, signal_1544}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1345 ( .s (signal_1225), .b ({ciphertext_s1[10], ciphertext_s0[10]}), .a ({signal_2532, signal_1671}), .c ({signal_2828, signal_1543}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1346 ( .s (signal_1225), .b ({ciphertext_s1[11], ciphertext_s0[11]}), .a ({signal_2535, signal_1670}), .c ({signal_2829, signal_1542}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1347 ( .s (signal_1225), .b ({ciphertext_s1[12], ciphertext_s0[12]}), .a ({signal_2538, signal_1669}), .c ({signal_2830, signal_1541}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1348 ( .s (signal_1225), .b ({ciphertext_s1[13], ciphertext_s0[13]}), .a ({signal_2541, signal_1668}), .c ({signal_2831, signal_1540}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1349 ( .s (signal_1225), .b ({ciphertext_s1[14], ciphertext_s0[14]}), .a ({signal_2544, signal_1667}), .c ({signal_2832, signal_1539}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1350 ( .s (signal_1225), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .a ({signal_2547, signal_1666}), .c ({signal_2833, signal_1538}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1351 ( .s (signal_1225), .b ({ciphertext_s1[48], ciphertext_s0[48]}), .a ({signal_2658, signal_1665}), .c ({signal_2834, signal_1537}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1352 ( .s (signal_1225), .b ({ciphertext_s1[49], ciphertext_s0[49]}), .a ({signal_2661, signal_1664}), .c ({signal_2835, signal_1536}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1353 ( .s (signal_1225), .b ({ciphertext_s1[50], ciphertext_s0[50]}), .a ({signal_2664, signal_1663}), .c ({signal_2836, signal_1535}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1354 ( .s (signal_1225), .b ({ciphertext_s1[51], ciphertext_s0[51]}), .a ({signal_2667, signal_1662}), .c ({signal_2837, signal_1534}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1355 ( .s (signal_1226), .b ({ciphertext_s1[52], ciphertext_s0[52]}), .a ({signal_2670, signal_1661}), .c ({signal_2838, signal_1533}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1356 ( .s (signal_1226), .b ({ciphertext_s1[53], ciphertext_s0[53]}), .a ({signal_2673, signal_1660}), .c ({signal_2839, signal_1532}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1357 ( .s (signal_1226), .b ({ciphertext_s1[54], ciphertext_s0[54]}), .a ({signal_2676, signal_1659}), .c ({signal_2840, signal_1531}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1358 ( .s (signal_1226), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .a ({signal_2679, signal_1658}), .c ({signal_2841, signal_1530}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1359 ( .s (signal_1226), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .a ({signal_2409, signal_1657}), .c ({signal_2842, signal_1529}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1360 ( .s (signal_1226), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .a ({signal_2412, signal_1656}), .c ({signal_2843, signal_1528}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1361 ( .s (signal_1226), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .a ({signal_2415, signal_1655}), .c ({signal_2844, signal_1527}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1362 ( .s (signal_1226), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .a ({signal_2418, signal_1654}), .c ({signal_2845, signal_1526}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1363 ( .s (signal_1226), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .a ({signal_2421, signal_1653}), .c ({signal_2846, signal_1525}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1364 ( .s (signal_1226), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .a ({signal_2424, signal_1652}), .c ({signal_2847, signal_1524}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1365 ( .s (signal_1226), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .a ({signal_2427, signal_1651}), .c ({signal_2848, signal_1523}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1366 ( .s (signal_1226), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .a ({signal_2430, signal_1650}), .c ({signal_2849, signal_1522}) ) ;
    INV_X1 cell_1887 ( .A (signal_1483), .ZN (signal_1490) ) ;
    INV_X1 cell_1888 ( .A (signal_393), .ZN (signal_1483) ) ;
    INV_X1 cell_1889 ( .A (signal_1483), .ZN (signal_1488) ) ;
    INV_X1 cell_1890 ( .A (signal_1483), .ZN (signal_1487) ) ;
    INV_X1 cell_1891 ( .A (signal_1483), .ZN (signal_1486) ) ;
    INV_X1 cell_1892 ( .A (signal_1483), .ZN (signal_1485) ) ;
    INV_X1 cell_1893 ( .A (signal_1483), .ZN (signal_1484) ) ;
    INV_X1 cell_1894 ( .A (signal_1483), .ZN (signal_1489) ) ;
    NOR2_X1 cell_2023 ( .A1 (reset), .A2 (signal_1491), .ZN (signal_1502) ) ;
    XNOR2_X1 cell_2024 ( .A (signal_2273), .B (signal_393), .ZN (signal_1491) ) ;
    NOR2_X1 cell_2025 ( .A1 (reset), .A2 (signal_1492), .ZN (signal_1501) ) ;
    XOR2_X1 cell_2026 ( .A (signal_2272), .B (signal_1493), .Z (signal_1492) ) ;
    NOR2_X1 cell_2027 ( .A1 (reset), .A2 (signal_1494), .ZN (signal_1498) ) ;
    XOR2_X1 cell_2028 ( .A (signal_2270), .B (signal_1495), .Z (signal_1494) ) ;
    NAND2_X1 cell_2029 ( .A1 (signal_1496), .A2 (signal_2271), .ZN (signal_1495) ) ;
    NOR2_X1 cell_2030 ( .A1 (reset), .A2 (signal_1497), .ZN (signal_1499) ) ;
    XNOR2_X1 cell_2031 ( .A (signal_2271), .B (signal_1496), .ZN (signal_1497) ) ;
    NOR2_X1 cell_2032 ( .A1 (signal_1500), .A2 (signal_1493), .ZN (signal_1496) ) ;
    NAND2_X1 cell_2033 ( .A1 (signal_393), .A2 (signal_2273), .ZN (signal_1493) ) ;
    INV_X1 cell_2036 ( .A (signal_2272), .ZN (signal_1500) ) ;
    NOR2_X1 cell_2042 ( .A1 (reset), .A2 (signal_1506), .ZN (signal_1520) ) ;
    XOR2_X1 cell_2043 ( .A (signal_2276), .B (signal_1507), .Z (signal_1506) ) ;
    NAND2_X1 cell_2044 ( .A1 (signal_1508), .A2 (1'b1), .ZN (signal_1507) ) ;
    NAND2_X1 cell_2045 ( .A1 (signal_1509), .A2 (signal_2274), .ZN (signal_1508) ) ;
    NAND2_X1 cell_2046 ( .A1 (signal_2276), .A2 (signal_2275), .ZN (signal_1509) ) ;
    NOR2_X1 cell_2047 ( .A1 (reset), .A2 (signal_1510), .ZN (signal_1519) ) ;
    MUX2_X1 cell_2048 ( .S (signal_2275), .A (signal_1511), .B (signal_1512), .Z (signal_1510) ) ;
    NOR2_X1 cell_2049 ( .A1 (reset), .A2 (signal_1513), .ZN (signal_1518) ) ;
    NOR2_X1 cell_2050 ( .A1 (signal_1514), .A2 (signal_1515), .ZN (signal_1513) ) ;
    NOR2_X1 cell_2051 ( .A1 (signal_1516), .A2 (signal_1511), .ZN (signal_1515) ) ;
    NAND2_X1 cell_2052 ( .A1 (signal_1512), .A2 (signal_1517), .ZN (signal_1511) ) ;
    AND2_X1 cell_2053 ( .A1 (signal_2276), .A2 (1'b1), .ZN (signal_1512) ) ;
    NOR2_X1 cell_2054 ( .A1 (1'b1), .A2 (signal_1517), .ZN (signal_1514) ) ;
    INV_X1 cell_2057 ( .A (signal_2275), .ZN (signal_1516) ) ;
    INV_X1 cell_2059 ( .A (signal_2274), .ZN (signal_1517) ) ;
    ClockGatingController #(3) cell_2062 ( .clk (clk), .rst (reset), .GatedClk (signal_3792), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_160 ( .s (reset), .b ({signal_3322, signal_1649}), .a ({plaintext_s1[0], plaintext_s0[0]}), .c ({signal_3437, signal_414}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_163 ( .s (reset), .b ({signal_3176, signal_1648}), .a ({plaintext_s1[1], plaintext_s0[1]}), .c ({signal_3263, signal_416}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_166 ( .s (reset), .b ({signal_3177, signal_1647}), .a ({plaintext_s1[2], plaintext_s0[2]}), .c ({signal_3265, signal_418}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_169 ( .s (reset), .b ({signal_3178, signal_1646}), .a ({plaintext_s1[3], plaintext_s0[3]}), .c ({signal_3267, signal_420}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_172 ( .s (reset), .b ({signal_3179, signal_1645}), .a ({plaintext_s1[4], plaintext_s0[4]}), .c ({signal_3269, signal_422}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_175 ( .s (reset), .b ({signal_3180, signal_1644}), .a ({plaintext_s1[5], plaintext_s0[5]}), .c ({signal_3271, signal_424}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_178 ( .s (reset), .b ({signal_3181, signal_1643}), .a ({plaintext_s1[6], plaintext_s0[6]}), .c ({signal_3273, signal_426}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_181 ( .s (reset), .b ({signal_3182, signal_1642}), .a ({plaintext_s1[7], plaintext_s0[7]}), .c ({signal_3275, signal_428}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_184 ( .s (reset), .b ({signal_3183, signal_1641}), .a ({plaintext_s1[8], plaintext_s0[8]}), .c ({signal_3277, signal_430}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_187 ( .s (reset), .b ({signal_3323, signal_1640}), .a ({plaintext_s1[9], plaintext_s0[9]}), .c ({signal_3439, signal_432}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_190 ( .s (reset), .b ({signal_3184, signal_1639}), .a ({plaintext_s1[10], plaintext_s0[10]}), .c ({signal_3279, signal_434}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_193 ( .s (reset), .b ({signal_3185, signal_1638}), .a ({plaintext_s1[11], plaintext_s0[11]}), .c ({signal_3281, signal_436}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_196 ( .s (reset), .b ({signal_3186, signal_1637}), .a ({plaintext_s1[12], plaintext_s0[12]}), .c ({signal_3283, signal_438}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_199 ( .s (reset), .b ({signal_3187, signal_1636}), .a ({plaintext_s1[13], plaintext_s0[13]}), .c ({signal_3285, signal_440}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_202 ( .s (reset), .b ({signal_3188, signal_1635}), .a ({plaintext_s1[14], plaintext_s0[14]}), .c ({signal_3287, signal_442}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_205 ( .s (reset), .b ({signal_3189, signal_1634}), .a ({plaintext_s1[15], plaintext_s0[15]}), .c ({signal_3289, signal_444}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_208 ( .s (reset), .b ({signal_3190, signal_1633}), .a ({plaintext_s1[16], plaintext_s0[16]}), .c ({signal_3291, signal_446}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_211 ( .s (reset), .b ({signal_3191, signal_1632}), .a ({plaintext_s1[17], plaintext_s0[17]}), .c ({signal_3293, signal_448}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_214 ( .s (reset), .b ({signal_3192, signal_1631}), .a ({plaintext_s1[18], plaintext_s0[18]}), .c ({signal_3295, signal_450}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_217 ( .s (reset), .b ({signal_3193, signal_1630}), .a ({plaintext_s1[19], plaintext_s0[19]}), .c ({signal_3297, signal_452}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_220 ( .s (reset), .b ({signal_3194, signal_1629}), .a ({plaintext_s1[20], plaintext_s0[20]}), .c ({signal_3299, signal_454}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_223 ( .s (reset), .b ({signal_3195, signal_1628}), .a ({plaintext_s1[21], plaintext_s0[21]}), .c ({signal_3301, signal_456}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_226 ( .s (reset), .b ({signal_3196, signal_1627}), .a ({plaintext_s1[22], plaintext_s0[22]}), .c ({signal_3303, signal_458}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_229 ( .s (reset), .b ({signal_3197, signal_1626}), .a ({plaintext_s1[23], plaintext_s0[23]}), .c ({signal_3305, signal_460}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_232 ( .s (reset), .b ({signal_3198, signal_1625}), .a ({plaintext_s1[24], plaintext_s0[24]}), .c ({signal_3307, signal_462}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_235 ( .s (reset), .b ({signal_3199, signal_1624}), .a ({plaintext_s1[25], plaintext_s0[25]}), .c ({signal_3309, signal_464}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_238 ( .s (reset), .b ({signal_3200, signal_1623}), .a ({plaintext_s1[26], plaintext_s0[26]}), .c ({signal_3311, signal_466}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_241 ( .s (reset), .b ({signal_3201, signal_1622}), .a ({plaintext_s1[27], plaintext_s0[27]}), .c ({signal_3313, signal_468}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_244 ( .s (reset), .b ({signal_3202, signal_1621}), .a ({plaintext_s1[28], plaintext_s0[28]}), .c ({signal_3315, signal_470}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_247 ( .s (reset), .b ({signal_3203, signal_1620}), .a ({plaintext_s1[29], plaintext_s0[29]}), .c ({signal_3317, signal_472}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_250 ( .s (reset), .b ({signal_3204, signal_1619}), .a ({plaintext_s1[30], plaintext_s0[30]}), .c ({signal_3319, signal_474}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_253 ( .s (reset), .b ({signal_3205, signal_1618}), .a ({plaintext_s1[31], plaintext_s0[31]}), .c ({signal_3321, signal_476}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1089 ( .a ({signal_3046, signal_1153}), .b ({signal_3100, signal_2328}), .c ({signal_3110, signal_1868}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) cell_1181 ( .a ({signal_3047, signal_1216}), .b ({signal_3093, signal_2321}), .c ({signal_3111, signal_1877}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1200 ( .s (signal_1218), .b ({signal_3111, signal_1877}), .a ({signal_3050, signal_1845}), .c ({signal_3174, signal_1909}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1201 ( .s (signal_394), .b ({signal_3080, signal_1876}), .a ({signal_3084, signal_2303}), .c ({signal_3112, signal_1908}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1202 ( .s (signal_394), .b ({signal_3079, signal_1875}), .a ({signal_3049, signal_1843}), .c ({signal_3113, signal_1907}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1203 ( .s (signal_394), .b ({signal_3078, signal_1874}), .a ({signal_3048, signal_1842}), .c ({signal_3114, signal_1906}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1204 ( .s (signal_394), .b ({signal_3077, signal_1873}), .a ({signal_3083, signal_2300}), .c ({signal_3115, signal_1905}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1205 ( .s (signal_394), .b ({signal_3076, signal_1872}), .a ({signal_3082, signal_2299}), .c ({signal_3116, signal_1904}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1206 ( .s (signal_394), .b ({signal_3075, signal_1871}), .a ({signal_3081, signal_2298}), .c ({signal_3117, signal_1903}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1207 ( .s (signal_1219), .b ({signal_3074, signal_1870}), .a ({signal_3085, signal_2305}), .c ({signal_3118, signal_1902}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1208 ( .s (signal_1218), .b ({signal_3073, signal_1869}), .a ({signal_3093, signal_2321}), .c ({signal_3119, signal_1901}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1209 ( .s (signal_1218), .b ({signal_3110, signal_1868}), .a ({signal_3092, signal_2320}), .c ({signal_3175, signal_1900}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1210 ( .s (signal_1218), .b ({signal_3072, signal_1867}), .a ({signal_3091, signal_2319}), .c ({signal_3120, signal_1899}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1211 ( .s (signal_1218), .b ({signal_3071, signal_1866}), .a ({signal_3090, signal_2318}), .c ({signal_3121, signal_1898}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1212 ( .s (signal_1218), .b ({signal_3070, signal_1865}), .a ({signal_3089, signal_2317}), .c ({signal_3122, signal_1897}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1213 ( .s (signal_1218), .b ({signal_3069, signal_1864}), .a ({signal_3088, signal_2316}), .c ({signal_3123, signal_1896}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1214 ( .s (signal_1218), .b ({signal_3068, signal_1863}), .a ({signal_3087, signal_2315}), .c ({signal_3124, signal_1895}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1215 ( .s (signal_1218), .b ({signal_3067, signal_1862}), .a ({signal_3086, signal_2314}), .c ({signal_3125, signal_1894}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1216 ( .s (signal_1218), .b ({signal_3066, signal_1861}), .a ({signal_3101, signal_2329}), .c ({signal_3126, signal_1893}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1217 ( .s (signal_1218), .b ({signal_3065, signal_1860}), .a ({signal_3100, signal_2328}), .c ({signal_3127, signal_1892}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1218 ( .s (signal_1218), .b ({signal_3064, signal_1859}), .a ({signal_3099, signal_2327}), .c ({signal_3128, signal_1891}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1219 ( .s (signal_1218), .b ({signal_3063, signal_1858}), .a ({signal_3098, signal_2326}), .c ({signal_3129, signal_1890}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1220 ( .s (signal_1219), .b ({signal_3062, signal_1857}), .a ({signal_3097, signal_2325}), .c ({signal_3130, signal_1889}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1221 ( .s (signal_1219), .b ({signal_3061, signal_1856}), .a ({signal_3096, signal_2324}), .c ({signal_3131, signal_1888}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1222 ( .s (signal_1219), .b ({signal_3060, signal_1855}), .a ({signal_3095, signal_2323}), .c ({signal_3132, signal_1887}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1223 ( .s (signal_1219), .b ({signal_3059, signal_1854}), .a ({signal_3094, signal_2322}), .c ({signal_3133, signal_1886}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1224 ( .s (signal_1219), .b ({signal_3058, signal_1853}), .a ({signal_3109, signal_2337}), .c ({signal_3134, signal_1885}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1225 ( .s (signal_1219), .b ({signal_3057, signal_1852}), .a ({signal_3108, signal_2336}), .c ({signal_3135, signal_1884}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1226 ( .s (signal_1219), .b ({signal_3056, signal_1851}), .a ({signal_3107, signal_2335}), .c ({signal_3136, signal_1883}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1227 ( .s (signal_1219), .b ({signal_3055, signal_1850}), .a ({signal_3106, signal_2334}), .c ({signal_3137, signal_1882}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1228 ( .s (signal_1219), .b ({signal_3054, signal_1849}), .a ({signal_3105, signal_2333}), .c ({signal_3138, signal_1881}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1229 ( .s (signal_1219), .b ({signal_3053, signal_1848}), .a ({signal_3104, signal_2332}), .c ({signal_3139, signal_1880}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1230 ( .s (signal_1219), .b ({signal_3052, signal_1847}), .a ({signal_3103, signal_2331}), .c ({signal_3140, signal_1879}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1231 ( .s (signal_1219), .b ({signal_3051, signal_1846}), .a ({signal_3102, signal_2330}), .c ({signal_3141, signal_1878}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1239 ( .s (signal_393), .b ({signal_3174, signal_1909}), .a ({signal_2499, signal_1777}), .c ({signal_3322, signal_1649}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1240 ( .s (signal_1226), .b ({signal_3112, signal_1908}), .a ({signal_2502, signal_1776}), .c ({signal_3176, signal_1648}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1241 ( .s (signal_1225), .b ({signal_3113, signal_1907}), .a ({signal_2505, signal_1775}), .c ({signal_3177, signal_1647}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1242 ( .s (signal_1224), .b ({signal_3114, signal_1906}), .a ({signal_2508, signal_1774}), .c ({signal_3178, signal_1646}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1243 ( .s (signal_1223), .b ({signal_3115, signal_1905}), .a ({signal_2511, signal_1773}), .c ({signal_3179, signal_1645}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1244 ( .s (signal_1222), .b ({signal_3116, signal_1904}), .a ({signal_2514, signal_1772}), .c ({signal_3180, signal_1644}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1245 ( .s (signal_1221), .b ({signal_3117, signal_1903}), .a ({signal_2517, signal_1771}), .c ({signal_3181, signal_1643}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1246 ( .s (signal_1226), .b ({signal_3118, signal_1902}), .a ({signal_2520, signal_1770}), .c ({signal_3182, signal_1642}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1247 ( .s (signal_1223), .b ({signal_3119, signal_1901}), .a ({signal_2631, signal_1769}), .c ({signal_3183, signal_1641}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1248 ( .s (signal_1226), .b ({signal_3175, signal_1900}), .a ({signal_2634, signal_1768}), .c ({signal_3323, signal_1640}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1249 ( .s (signal_393), .b ({signal_3120, signal_1899}), .a ({signal_2637, signal_1767}), .c ({signal_3184, signal_1639}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1250 ( .s (signal_393), .b ({signal_3121, signal_1898}), .a ({signal_2640, signal_1766}), .c ({signal_3185, signal_1638}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1251 ( .s (signal_393), .b ({signal_3122, signal_1897}), .a ({signal_2643, signal_1765}), .c ({signal_3186, signal_1637}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1252 ( .s (signal_393), .b ({signal_3123, signal_1896}), .a ({signal_2646, signal_1764}), .c ({signal_3187, signal_1636}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1253 ( .s (signal_393), .b ({signal_3124, signal_1895}), .a ({signal_2649, signal_1763}), .c ({signal_3188, signal_1635}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1254 ( .s (signal_393), .b ({signal_3125, signal_1894}), .a ({signal_2652, signal_1762}), .c ({signal_3189, signal_1634}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1255 ( .s (signal_393), .b ({signal_3126, signal_1893}), .a ({signal_2382, signal_1761}), .c ({signal_3190, signal_1633}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1256 ( .s (signal_393), .b ({signal_3127, signal_1892}), .a ({signal_2385, signal_1760}), .c ({signal_3191, signal_1632}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1257 ( .s (signal_393), .b ({signal_3128, signal_1891}), .a ({signal_2388, signal_1759}), .c ({signal_3192, signal_1631}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1258 ( .s (signal_393), .b ({signal_3129, signal_1890}), .a ({signal_2391, signal_1758}), .c ({signal_3193, signal_1630}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1259 ( .s (signal_1225), .b ({signal_3130, signal_1889}), .a ({signal_2394, signal_1757}), .c ({signal_3194, signal_1629}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1260 ( .s (signal_1224), .b ({signal_3131, signal_1888}), .a ({signal_2397, signal_1756}), .c ({signal_3195, signal_1628}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1261 ( .s (signal_1223), .b ({signal_3132, signal_1887}), .a ({signal_2400, signal_1755}), .c ({signal_3196, signal_1627}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1262 ( .s (signal_1222), .b ({signal_3133, signal_1886}), .a ({signal_2403, signal_1754}), .c ({signal_3197, signal_1626}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1263 ( .s (signal_1221), .b ({signal_3134, signal_1885}), .a ({signal_2472, signal_1753}), .c ({signal_3198, signal_1625}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1264 ( .s (signal_1223), .b ({signal_3135, signal_1884}), .a ({signal_2475, signal_1752}), .c ({signal_3199, signal_1624}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1265 ( .s (signal_1222), .b ({signal_3136, signal_1883}), .a ({signal_2478, signal_1751}), .c ({signal_3200, signal_1623}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1266 ( .s (signal_393), .b ({signal_3137, signal_1882}), .a ({signal_2481, signal_1750}), .c ({signal_3201, signal_1622}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1267 ( .s (signal_393), .b ({signal_3138, signal_1881}), .a ({signal_2484, signal_1749}), .c ({signal_3202, signal_1621}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1268 ( .s (signal_1226), .b ({signal_3139, signal_1880}), .a ({signal_2487, signal_1748}), .c ({signal_3203, signal_1620}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1269 ( .s (signal_1225), .b ({signal_3140, signal_1879}), .a ({signal_2493, signal_1747}), .c ({signal_3204, signal_1619}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1270 ( .s (signal_1224), .b ({signal_3141, signal_1878}), .a ({signal_2496, signal_1746}), .c ({signal_3205, signal_1618}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1369 ( .s (reset), .b ({signal_3640, signal_2037}), .a ({key_s1[0], key_s0[0]}), .c ({signal_3673, signal_1227}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1372 ( .s (reset), .b ({signal_3641, signal_2036}), .a ({key_s1[1], key_s0[1]}), .c ({signal_3675, signal_1229}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1375 ( .s (reset), .b ({signal_3642, signal_2035}), .a ({key_s1[2], key_s0[2]}), .c ({signal_3677, signal_1231}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1378 ( .s (reset), .b ({signal_3643, signal_2034}), .a ({key_s1[3], key_s0[3]}), .c ({signal_3679, signal_1233}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1381 ( .s (reset), .b ({signal_3644, signal_2033}), .a ({key_s1[4], key_s0[4]}), .c ({signal_3681, signal_1235}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1384 ( .s (reset), .b ({signal_3645, signal_2032}), .a ({key_s1[5], key_s0[5]}), .c ({signal_3683, signal_1237}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1387 ( .s (reset), .b ({signal_3646, signal_2031}), .a ({key_s1[6], key_s0[6]}), .c ({signal_3685, signal_1239}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1390 ( .s (reset), .b ({signal_3647, signal_2030}), .a ({key_s1[7], key_s0[7]}), .c ({signal_3687, signal_1241}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1393 ( .s (reset), .b ({signal_3648, signal_2029}), .a ({key_s1[8], key_s0[8]}), .c ({signal_3689, signal_1243}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1396 ( .s (reset), .b ({signal_3649, signal_2028}), .a ({key_s1[9], key_s0[9]}), .c ({signal_3691, signal_1245}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1399 ( .s (reset), .b ({signal_3650, signal_2027}), .a ({key_s1[10], key_s0[10]}), .c ({signal_3693, signal_1247}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1402 ( .s (reset), .b ({signal_3651, signal_2026}), .a ({key_s1[11], key_s0[11]}), .c ({signal_3695, signal_1249}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1405 ( .s (reset), .b ({signal_3652, signal_2025}), .a ({key_s1[12], key_s0[12]}), .c ({signal_3697, signal_1251}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1408 ( .s (reset), .b ({signal_3653, signal_2024}), .a ({key_s1[13], key_s0[13]}), .c ({signal_3699, signal_1253}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1411 ( .s (reset), .b ({signal_3654, signal_2023}), .a ({key_s1[14], key_s0[14]}), .c ({signal_3701, signal_1255}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1414 ( .s (reset), .b ({signal_3655, signal_2022}), .a ({key_s1[15], key_s0[15]}), .c ({signal_3703, signal_1257}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1417 ( .s (reset), .b ({signal_3656, signal_2021}), .a ({key_s1[16], key_s0[16]}), .c ({signal_3705, signal_1259}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1420 ( .s (reset), .b ({signal_3657, signal_2020}), .a ({key_s1[17], key_s0[17]}), .c ({signal_3707, signal_1261}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1423 ( .s (reset), .b ({signal_3658, signal_2019}), .a ({key_s1[18], key_s0[18]}), .c ({signal_3709, signal_1263}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1426 ( .s (reset), .b ({signal_3659, signal_2018}), .a ({key_s1[19], key_s0[19]}), .c ({signal_3711, signal_1265}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1429 ( .s (reset), .b ({signal_3660, signal_2017}), .a ({key_s1[20], key_s0[20]}), .c ({signal_3713, signal_1267}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1432 ( .s (reset), .b ({signal_3661, signal_2016}), .a ({key_s1[21], key_s0[21]}), .c ({signal_3715, signal_1269}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1435 ( .s (reset), .b ({signal_3662, signal_2015}), .a ({key_s1[22], key_s0[22]}), .c ({signal_3717, signal_1271}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1438 ( .s (reset), .b ({signal_3663, signal_2014}), .a ({key_s1[23], key_s0[23]}), .c ({signal_3719, signal_1273}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1441 ( .s (reset), .b ({signal_3736, signal_2013}), .a ({key_s1[24], key_s0[24]}), .c ({signal_3745, signal_1275}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1444 ( .s (reset), .b ({signal_3737, signal_2012}), .a ({key_s1[25], key_s0[25]}), .c ({signal_3747, signal_1277}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1447 ( .s (reset), .b ({signal_3738, signal_2011}), .a ({key_s1[26], key_s0[26]}), .c ({signal_3749, signal_1279}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1450 ( .s (reset), .b ({signal_3739, signal_2010}), .a ({key_s1[27], key_s0[27]}), .c ({signal_3751, signal_1281}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1453 ( .s (reset), .b ({signal_3740, signal_2009}), .a ({key_s1[28], key_s0[28]}), .c ({signal_3753, signal_1283}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1456 ( .s (reset), .b ({signal_3741, signal_2008}), .a ({key_s1[29], key_s0[29]}), .c ({signal_3755, signal_1285}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1459 ( .s (reset), .b ({signal_3742, signal_2007}), .a ({key_s1[30], key_s0[30]}), .c ({signal_3757, signal_1287}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1462 ( .s (reset), .b ({signal_3743, signal_2006}), .a ({key_s1[31], key_s0[31]}), .c ({signal_3759, signal_1289}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1465 ( .s (reset), .b ({signal_3536, signal_2005}), .a ({key_s1[32], key_s0[32]}), .c ({signal_3569, signal_1291}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1468 ( .s (reset), .b ({signal_3537, signal_2004}), .a ({key_s1[33], key_s0[33]}), .c ({signal_3571, signal_1293}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1471 ( .s (reset), .b ({signal_3538, signal_2003}), .a ({key_s1[34], key_s0[34]}), .c ({signal_3573, signal_1295}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1474 ( .s (reset), .b ({signal_3539, signal_2002}), .a ({key_s1[35], key_s0[35]}), .c ({signal_3575, signal_1297}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1477 ( .s (reset), .b ({signal_3540, signal_2001}), .a ({key_s1[36], key_s0[36]}), .c ({signal_3577, signal_1299}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1480 ( .s (reset), .b ({signal_3541, signal_2000}), .a ({key_s1[37], key_s0[37]}), .c ({signal_3579, signal_1301}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1483 ( .s (reset), .b ({signal_3542, signal_1999}), .a ({key_s1[38], key_s0[38]}), .c ({signal_3581, signal_1303}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1486 ( .s (reset), .b ({signal_3543, signal_1998}), .a ({key_s1[39], key_s0[39]}), .c ({signal_3583, signal_1305}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1489 ( .s (reset), .b ({signal_3544, signal_1997}), .a ({key_s1[40], key_s0[40]}), .c ({signal_3585, signal_1307}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1492 ( .s (reset), .b ({signal_3545, signal_1996}), .a ({key_s1[41], key_s0[41]}), .c ({signal_3587, signal_1309}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1495 ( .s (reset), .b ({signal_3546, signal_1995}), .a ({key_s1[42], key_s0[42]}), .c ({signal_3589, signal_1311}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1498 ( .s (reset), .b ({signal_3547, signal_1994}), .a ({key_s1[43], key_s0[43]}), .c ({signal_3591, signal_1313}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1501 ( .s (reset), .b ({signal_3548, signal_1993}), .a ({key_s1[44], key_s0[44]}), .c ({signal_3593, signal_1315}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1504 ( .s (reset), .b ({signal_3549, signal_1992}), .a ({key_s1[45], key_s0[45]}), .c ({signal_3595, signal_1317}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1507 ( .s (reset), .b ({signal_3550, signal_1991}), .a ({key_s1[46], key_s0[46]}), .c ({signal_3597, signal_1319}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1510 ( .s (reset), .b ({signal_3551, signal_1990}), .a ({key_s1[47], key_s0[47]}), .c ({signal_3599, signal_1321}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1513 ( .s (reset), .b ({signal_3552, signal_1989}), .a ({key_s1[48], key_s0[48]}), .c ({signal_3601, signal_1323}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1516 ( .s (reset), .b ({signal_3553, signal_1988}), .a ({key_s1[49], key_s0[49]}), .c ({signal_3603, signal_1325}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1519 ( .s (reset), .b ({signal_3554, signal_1987}), .a ({key_s1[50], key_s0[50]}), .c ({signal_3605, signal_1327}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1522 ( .s (reset), .b ({signal_3555, signal_1986}), .a ({key_s1[51], key_s0[51]}), .c ({signal_3607, signal_1329}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1525 ( .s (reset), .b ({signal_3556, signal_1985}), .a ({key_s1[52], key_s0[52]}), .c ({signal_3609, signal_1331}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1528 ( .s (reset), .b ({signal_3557, signal_1984}), .a ({key_s1[53], key_s0[53]}), .c ({signal_3611, signal_1333}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1531 ( .s (reset), .b ({signal_3558, signal_1983}), .a ({key_s1[54], key_s0[54]}), .c ({signal_3613, signal_1335}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1534 ( .s (reset), .b ({signal_3559, signal_1982}), .a ({key_s1[55], key_s0[55]}), .c ({signal_3615, signal_1337}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1537 ( .s (reset), .b ({signal_3664, signal_1981}), .a ({key_s1[56], key_s0[56]}), .c ({signal_3721, signal_1339}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1540 ( .s (reset), .b ({signal_3665, signal_1980}), .a ({key_s1[57], key_s0[57]}), .c ({signal_3723, signal_1341}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1543 ( .s (reset), .b ({signal_3666, signal_1979}), .a ({key_s1[58], key_s0[58]}), .c ({signal_3725, signal_1343}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1546 ( .s (reset), .b ({signal_3667, signal_1978}), .a ({key_s1[59], key_s0[59]}), .c ({signal_3727, signal_1345}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1549 ( .s (reset), .b ({signal_3668, signal_1977}), .a ({key_s1[60], key_s0[60]}), .c ({signal_3729, signal_1347}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1552 ( .s (reset), .b ({signal_3669, signal_1976}), .a ({key_s1[61], key_s0[61]}), .c ({signal_3731, signal_1349}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1555 ( .s (reset), .b ({signal_3670, signal_1975}), .a ({key_s1[62], key_s0[62]}), .c ({signal_3733, signal_1351}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1558 ( .s (reset), .b ({signal_3671, signal_1974}), .a ({key_s1[63], key_s0[63]}), .c ({signal_3735, signal_1353}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1561 ( .s (reset), .b ({signal_3404, signal_1973}), .a ({key_s1[64], key_s0[64]}), .c ({signal_3441, signal_1355}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1564 ( .s (reset), .b ({signal_3405, signal_1972}), .a ({key_s1[65], key_s0[65]}), .c ({signal_3443, signal_1357}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1567 ( .s (reset), .b ({signal_3406, signal_1971}), .a ({key_s1[66], key_s0[66]}), .c ({signal_3445, signal_1359}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1570 ( .s (reset), .b ({signal_3407, signal_1970}), .a ({key_s1[67], key_s0[67]}), .c ({signal_3447, signal_1361}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1573 ( .s (reset), .b ({signal_3408, signal_1969}), .a ({key_s1[68], key_s0[68]}), .c ({signal_3449, signal_1363}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1576 ( .s (reset), .b ({signal_3409, signal_1968}), .a ({key_s1[69], key_s0[69]}), .c ({signal_3451, signal_1365}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1579 ( .s (reset), .b ({signal_3410, signal_1967}), .a ({key_s1[70], key_s0[70]}), .c ({signal_3453, signal_1367}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1582 ( .s (reset), .b ({signal_3411, signal_1966}), .a ({key_s1[71], key_s0[71]}), .c ({signal_3455, signal_1369}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1585 ( .s (reset), .b ({signal_3412, signal_1965}), .a ({key_s1[72], key_s0[72]}), .c ({signal_3457, signal_1371}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1588 ( .s (reset), .b ({signal_3413, signal_1964}), .a ({key_s1[73], key_s0[73]}), .c ({signal_3459, signal_1373}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1591 ( .s (reset), .b ({signal_3414, signal_1963}), .a ({key_s1[74], key_s0[74]}), .c ({signal_3461, signal_1375}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1594 ( .s (reset), .b ({signal_3415, signal_1962}), .a ({key_s1[75], key_s0[75]}), .c ({signal_3463, signal_1377}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1597 ( .s (reset), .b ({signal_3416, signal_1961}), .a ({key_s1[76], key_s0[76]}), .c ({signal_3465, signal_1379}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1600 ( .s (reset), .b ({signal_3417, signal_1960}), .a ({key_s1[77], key_s0[77]}), .c ({signal_3467, signal_1381}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1603 ( .s (reset), .b ({signal_3418, signal_1959}), .a ({key_s1[78], key_s0[78]}), .c ({signal_3469, signal_1383}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1606 ( .s (reset), .b ({signal_3419, signal_1958}), .a ({key_s1[79], key_s0[79]}), .c ({signal_3471, signal_1385}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1609 ( .s (reset), .b ({signal_3420, signal_1957}), .a ({key_s1[80], key_s0[80]}), .c ({signal_3473, signal_1387}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1612 ( .s (reset), .b ({signal_3421, signal_1956}), .a ({key_s1[81], key_s0[81]}), .c ({signal_3475, signal_1389}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1615 ( .s (reset), .b ({signal_3422, signal_1955}), .a ({key_s1[82], key_s0[82]}), .c ({signal_3477, signal_1391}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1618 ( .s (reset), .b ({signal_3423, signal_1954}), .a ({key_s1[83], key_s0[83]}), .c ({signal_3479, signal_1393}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1621 ( .s (reset), .b ({signal_3424, signal_1953}), .a ({key_s1[84], key_s0[84]}), .c ({signal_3481, signal_1395}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1624 ( .s (reset), .b ({signal_3425, signal_1952}), .a ({key_s1[85], key_s0[85]}), .c ({signal_3483, signal_1397}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1627 ( .s (reset), .b ({signal_3426, signal_1951}), .a ({key_s1[86], key_s0[86]}), .c ({signal_3485, signal_1399}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1630 ( .s (reset), .b ({signal_3427, signal_1950}), .a ({key_s1[87], key_s0[87]}), .c ({signal_3487, signal_1401}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1633 ( .s (reset), .b ({signal_3560, signal_1949}), .a ({key_s1[88], key_s0[88]}), .c ({signal_3617, signal_1403}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1636 ( .s (reset), .b ({signal_3561, signal_1948}), .a ({key_s1[89], key_s0[89]}), .c ({signal_3619, signal_1405}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1639 ( .s (reset), .b ({signal_3562, signal_1947}), .a ({key_s1[90], key_s0[90]}), .c ({signal_3621, signal_1407}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1642 ( .s (reset), .b ({signal_3563, signal_1946}), .a ({key_s1[91], key_s0[91]}), .c ({signal_3623, signal_1409}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1645 ( .s (reset), .b ({signal_3564, signal_1945}), .a ({key_s1[92], key_s0[92]}), .c ({signal_3625, signal_1411}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1648 ( .s (reset), .b ({signal_3565, signal_1944}), .a ({key_s1[93], key_s0[93]}), .c ({signal_3627, signal_1413}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1651 ( .s (reset), .b ({signal_3566, signal_1943}), .a ({key_s1[94], key_s0[94]}), .c ({signal_3629, signal_1415}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1654 ( .s (reset), .b ({signal_3567, signal_1942}), .a ({key_s1[95], key_s0[95]}), .c ({signal_3631, signal_1417}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1657 ( .s (reset), .b ({signal_3238, signal_1941}), .a ({key_s1[96], key_s0[96]}), .c ({signal_3325, signal_1419}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1660 ( .s (reset), .b ({signal_3239, signal_1940}), .a ({key_s1[97], key_s0[97]}), .c ({signal_3327, signal_1421}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1663 ( .s (reset), .b ({signal_3240, signal_1939}), .a ({key_s1[98], key_s0[98]}), .c ({signal_3329, signal_1423}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1666 ( .s (reset), .b ({signal_3241, signal_1938}), .a ({key_s1[99], key_s0[99]}), .c ({signal_3331, signal_1425}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1669 ( .s (reset), .b ({signal_3242, signal_1937}), .a ({key_s1[100], key_s0[100]}), .c ({signal_3333, signal_1427}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1672 ( .s (reset), .b ({signal_3243, signal_1936}), .a ({key_s1[101], key_s0[101]}), .c ({signal_3335, signal_1429}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1675 ( .s (reset), .b ({signal_3244, signal_1935}), .a ({key_s1[102], key_s0[102]}), .c ({signal_3337, signal_1431}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1678 ( .s (reset), .b ({signal_3245, signal_1934}), .a ({key_s1[103], key_s0[103]}), .c ({signal_3339, signal_1433}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1681 ( .s (reset), .b ({signal_3246, signal_1933}), .a ({key_s1[104], key_s0[104]}), .c ({signal_3341, signal_1435}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1684 ( .s (reset), .b ({signal_3247, signal_1932}), .a ({key_s1[105], key_s0[105]}), .c ({signal_3343, signal_1437}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1687 ( .s (reset), .b ({signal_3248, signal_1931}), .a ({key_s1[106], key_s0[106]}), .c ({signal_3345, signal_1439}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1690 ( .s (reset), .b ({signal_3249, signal_1930}), .a ({key_s1[107], key_s0[107]}), .c ({signal_3347, signal_1441}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1693 ( .s (reset), .b ({signal_3250, signal_1929}), .a ({key_s1[108], key_s0[108]}), .c ({signal_3349, signal_1443}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1696 ( .s (reset), .b ({signal_3251, signal_1928}), .a ({key_s1[109], key_s0[109]}), .c ({signal_3351, signal_1445}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1699 ( .s (reset), .b ({signal_3252, signal_1927}), .a ({key_s1[110], key_s0[110]}), .c ({signal_3353, signal_1447}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1702 ( .s (reset), .b ({signal_3253, signal_1926}), .a ({key_s1[111], key_s0[111]}), .c ({signal_3355, signal_1449}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1705 ( .s (reset), .b ({signal_3254, signal_1925}), .a ({key_s1[112], key_s0[112]}), .c ({signal_3357, signal_1451}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1708 ( .s (reset), .b ({signal_3255, signal_1924}), .a ({key_s1[113], key_s0[113]}), .c ({signal_3359, signal_1453}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1711 ( .s (reset), .b ({signal_3256, signal_1923}), .a ({key_s1[114], key_s0[114]}), .c ({signal_3361, signal_1455}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1714 ( .s (reset), .b ({signal_3257, signal_1922}), .a ({key_s1[115], key_s0[115]}), .c ({signal_3363, signal_1457}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1717 ( .s (reset), .b ({signal_3258, signal_1921}), .a ({key_s1[116], key_s0[116]}), .c ({signal_3365, signal_1459}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1720 ( .s (reset), .b ({signal_3259, signal_1920}), .a ({key_s1[117], key_s0[117]}), .c ({signal_3367, signal_1461}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1723 ( .s (reset), .b ({signal_3260, signal_1919}), .a ({key_s1[118], key_s0[118]}), .c ({signal_3369, signal_1463}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1726 ( .s (reset), .b ({signal_3261, signal_1918}), .a ({key_s1[119], key_s0[119]}), .c ({signal_3371, signal_1465}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1729 ( .s (reset), .b ({signal_3428, signal_1917}), .a ({key_s1[120], key_s0[120]}), .c ({signal_3489, signal_1467}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1732 ( .s (reset), .b ({signal_3429, signal_1916}), .a ({key_s1[121], key_s0[121]}), .c ({signal_3491, signal_1469}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1735 ( .s (reset), .b ({signal_3430, signal_1915}), .a ({key_s1[122], key_s0[122]}), .c ({signal_3493, signal_1471}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1738 ( .s (reset), .b ({signal_3431, signal_1914}), .a ({key_s1[123], key_s0[123]}), .c ({signal_3495, signal_1473}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1741 ( .s (reset), .b ({signal_3432, signal_1913}), .a ({key_s1[124], key_s0[124]}), .c ({signal_3497, signal_1475}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1744 ( .s (reset), .b ({signal_3433, signal_1912}), .a ({key_s1[125], key_s0[125]}), .c ({signal_3499, signal_1477}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1747 ( .s (reset), .b ({signal_3434, signal_1911}), .a ({key_s1[126], key_s0[126]}), .c ({signal_3501, signal_1479}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1750 ( .s (reset), .b ({signal_3435, signal_1910}), .a ({key_s1[127], key_s0[127]}), .c ({signal_3503, signal_1481}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1751 ( .a ({signal_2720, signal_1800}), .b ({signal_3372, signal_2228}), .c ({signal_3504, signal_2260}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1752 ( .a ({signal_2687, signal_1801}), .b ({signal_3373, signal_2229}), .c ({signal_3505, signal_2261}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1753 ( .a ({signal_2654, signal_1786}), .b ({signal_3374, signal_2230}), .c ({signal_3506, signal_2262}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1754 ( .a ({signal_2621, signal_1787}), .b ({signal_3375, signal_2231}), .c ({signal_3507, signal_2263}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1755 ( .a ({signal_2588, signal_1788}), .b ({signal_3376, signal_2232}), .c ({signal_3508, signal_2264}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1756 ( .a ({signal_2555, signal_1789}), .b ({signal_3377, signal_2233}), .c ({signal_3509, signal_2265}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1757 ( .a ({signal_2528, signal_2124}), .b ({signal_3206, signal_2196}), .c ({signal_3372, signal_2228}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1758 ( .a ({signal_2633, signal_2092}), .b ({signal_3159, signal_2164}), .c ({signal_3206, signal_2196}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1759 ( .a ({signal_2525, signal_2125}), .b ({signal_3207, signal_2197}), .c ({signal_3373, signal_2229}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1760 ( .a ({signal_2630, signal_2093}), .b ({signal_3160, signal_2165}), .c ({signal_3207, signal_2197}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1761 ( .a ({signal_2522, signal_1790}), .b ({signal_3378, signal_2234}), .c ({signal_3510, signal_2266}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1762 ( .a ({signal_2519, signal_2126}), .b ({signal_3208, signal_2198}), .c ({signal_3374, signal_2230}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1763 ( .a ({signal_2627, signal_2094}), .b ({signal_3161, signal_2166}), .c ({signal_3208, signal_2198}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1764 ( .a ({signal_2516, signal_2127}), .b ({signal_3209, signal_2199}), .c ({signal_3375, signal_2231}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1765 ( .a ({signal_2624, signal_2095}), .b ({signal_3162, signal_2167}), .c ({signal_3209, signal_2199}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1766 ( .a ({signal_2513, signal_2128}), .b ({signal_3210, signal_2200}), .c ({signal_3376, signal_2232}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1767 ( .a ({signal_2618, signal_2096}), .b ({signal_3163, signal_2168}), .c ({signal_3210, signal_2200}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1768 ( .a ({signal_2510, signal_2129}), .b ({signal_3211, signal_2201}), .c ({signal_3377, signal_2233}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1769 ( .a ({signal_2615, signal_2097}), .b ({signal_3164, signal_2169}), .c ({signal_3211, signal_2201}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1770 ( .a ({signal_2507, signal_2130}), .b ({signal_3212, signal_2202}), .c ({signal_3378, signal_2234}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1771 ( .a ({signal_2612, signal_2098}), .b ({signal_3142, signal_2170}), .c ({signal_3212, signal_2202}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1772 ( .a ({signal_2717, signal_2066}), .b ({signal_3106, signal_2334}), .c ({signal_3142, signal_2170}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1773 ( .a ({signal_2495, signal_1778}), .b ({signal_3511, signal_2206}), .c ({signal_3632, signal_2238}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1774 ( .a ({signal_2600, signal_2102}), .b ({signal_3379, signal_2174}), .c ({signal_3511, signal_2206}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1775 ( .a ({signal_2705, signal_2070}), .b ({signal_3227, signal_2142}), .c ({signal_3379, signal_2174}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1776 ( .a ({signal_2492, signal_1779}), .b ({signal_3512, signal_2207}), .c ({signal_3633, signal_2239}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1777 ( .a ({signal_2597, signal_2103}), .b ({signal_3380, signal_2175}), .c ({signal_3512, signal_2207}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1778 ( .a ({signal_2702, signal_2071}), .b ({signal_3228, signal_2143}), .c ({signal_3380, signal_2175}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1779 ( .a ({signal_2489, signal_1791}), .b ({signal_3381, signal_2235}), .c ({signal_3513, signal_2267}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1780 ( .a ({signal_2504, signal_2131}), .b ({signal_3213, signal_2203}), .c ({signal_3381, signal_2235}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1781 ( .a ({signal_2609, signal_2099}), .b ({signal_3143, signal_2171}), .c ({signal_3213, signal_2203}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1782 ( .a ({signal_2714, signal_2067}), .b ({signal_3107, signal_2335}), .c ({signal_3143, signal_2171}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1783 ( .a ({signal_2486, signal_1780}), .b ({signal_3514, signal_2208}), .c ({signal_3634, signal_2240}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1784 ( .a ({signal_2594, signal_2104}), .b ({signal_3382, signal_2176}), .c ({signal_3514, signal_2208}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1785 ( .a ({signal_2699, signal_2072}), .b ({signal_3229, signal_2144}), .c ({signal_3382, signal_2176}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1786 ( .a ({signal_2483, signal_1781}), .b ({signal_3515, signal_2209}), .c ({signal_3635, signal_2241}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1787 ( .a ({signal_2591, signal_2105}), .b ({signal_3383, signal_2177}), .c ({signal_3515, signal_2209}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1788 ( .a ({signal_2696, signal_2073}), .b ({signal_3230, signal_2145}), .c ({signal_3383, signal_2177}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1789 ( .a ({signal_2480, signal_1782}), .b ({signal_3516, signal_2210}), .c ({signal_3636, signal_2242}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1790 ( .a ({signal_2585, signal_2106}), .b ({signal_3384, signal_2178}), .c ({signal_3516, signal_2210}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1791 ( .a ({signal_2693, signal_2074}), .b ({signal_3231, signal_2146}), .c ({signal_3384, signal_2178}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1792 ( .a ({signal_2477, signal_1783}), .b ({signal_3517, signal_2211}), .c ({signal_3637, signal_2243}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1793 ( .a ({signal_2582, signal_2107}), .b ({signal_3385, signal_2179}), .c ({signal_3517, signal_2211}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1794 ( .a ({signal_2690, signal_2075}), .b ({signal_3232, signal_2147}), .c ({signal_3385, signal_2179}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1795 ( .a ({signal_2474, signal_1784}), .b ({signal_3518, signal_2212}), .c ({signal_3638, signal_2244}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1796 ( .a ({signal_2579, signal_2108}), .b ({signal_3386, signal_2180}), .c ({signal_3518, signal_2212}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1797 ( .a ({signal_2684, signal_2076}), .b ({signal_3233, signal_2148}), .c ({signal_3386, signal_2180}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1798 ( .a ({signal_2471, signal_1785}), .b ({signal_3519, signal_2213}), .c ({signal_3639, signal_2245}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1799 ( .a ({signal_2576, signal_2109}), .b ({signal_3387, signal_2181}), .c ({signal_3519, signal_2213}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1800 ( .a ({signal_2681, signal_2077}), .b ({signal_3234, signal_2149}), .c ({signal_3387, signal_2181}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1801 ( .a ({signal_2468, signal_1802}), .b ({signal_3388, signal_2214}), .c ({signal_3520, signal_2246}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1802 ( .a ({signal_2573, signal_2110}), .b ({signal_3214, signal_2182}), .c ({signal_3388, signal_2214}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1803 ( .a ({signal_2678, signal_2078}), .b ({signal_3145, signal_2150}), .c ({signal_3214, signal_2182}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1804 ( .a ({signal_2465, signal_1803}), .b ({signal_3389, signal_2215}), .c ({signal_3521, signal_2247}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1805 ( .a ({signal_2570, signal_2111}), .b ({signal_3215, signal_2183}), .c ({signal_3389, signal_2215}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1806 ( .a ({signal_2675, signal_2079}), .b ({signal_3146, signal_2151}), .c ({signal_3215, signal_2183}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1807 ( .a ({signal_2462, signal_1804}), .b ({signal_3390, signal_2216}), .c ({signal_3522, signal_2248}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1808 ( .a ({signal_2567, signal_2112}), .b ({signal_3216, signal_2184}), .c ({signal_3390, signal_2216}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1809 ( .a ({signal_2672, signal_2080}), .b ({signal_3147, signal_2152}), .c ({signal_3216, signal_2184}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1810 ( .a ({signal_2459, signal_1805}), .b ({signal_3391, signal_2217}), .c ({signal_3523, signal_2249}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1811 ( .a ({signal_2564, signal_2113}), .b ({signal_3217, signal_2185}), .c ({signal_3391, signal_2217}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1812 ( .a ({signal_2669, signal_2081}), .b ({signal_3148, signal_2153}), .c ({signal_3217, signal_2185}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1813 ( .a ({signal_2456, signal_1792}), .b ({signal_3392, signal_2236}), .c ({signal_3524, signal_2268}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1814 ( .a ({signal_2501, signal_2132}), .b ({signal_3218, signal_2204}), .c ({signal_3392, signal_2236}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1815 ( .a ({signal_2606, signal_2100}), .b ({signal_3144, signal_2172}), .c ({signal_3218, signal_2204}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1816 ( .a ({signal_2711, signal_2068}), .b ({signal_3108, signal_2336}), .c ({signal_3144, signal_2172}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1817 ( .a ({signal_2453, signal_1806}), .b ({signal_3393, signal_2218}), .c ({signal_3525, signal_2250}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1818 ( .a ({signal_2561, signal_2114}), .b ({signal_3219, signal_2186}), .c ({signal_3393, signal_2218}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1819 ( .a ({signal_2666, signal_2082}), .b ({signal_3149, signal_2154}), .c ({signal_3219, signal_2186}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1820 ( .a ({signal_2450, signal_1807}), .b ({signal_3394, signal_2219}), .c ({signal_3526, signal_2251}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1821 ( .a ({signal_2558, signal_2115}), .b ({signal_3220, signal_2187}), .c ({signal_3394, signal_2219}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1822 ( .a ({signal_2663, signal_2083}), .b ({signal_3150, signal_2155}), .c ({signal_3220, signal_2187}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1823 ( .a ({signal_2447, signal_1808}), .b ({signal_3395, signal_2220}), .c ({signal_3527, signal_2252}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1824 ( .a ({signal_2552, signal_2116}), .b ({signal_3221, signal_2188}), .c ({signal_3395, signal_2220}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1825 ( .a ({signal_2660, signal_2084}), .b ({signal_3151, signal_2156}), .c ({signal_3221, signal_2188}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1826 ( .a ({signal_2444, signal_1809}), .b ({signal_3396, signal_2221}), .c ({signal_3528, signal_2253}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1827 ( .a ({signal_2549, signal_2117}), .b ({signal_3222, signal_2189}), .c ({signal_3396, signal_2221}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1828 ( .a ({signal_2657, signal_2085}), .b ({signal_3152, signal_2157}), .c ({signal_3222, signal_2189}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1829 ( .a ({signal_2441, signal_1794}), .b ({signal_3397, signal_2222}), .c ({signal_3529, signal_2254}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1830 ( .a ({signal_2546, signal_2118}), .b ({signal_3223, signal_2190}), .c ({signal_3397, signal_2222}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1831 ( .a ({signal_2651, signal_2086}), .b ({signal_3153, signal_2158}), .c ({signal_3223, signal_2190}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1832 ( .a ({signal_2438, signal_1795}), .b ({signal_3398, signal_2223}), .c ({signal_3530, signal_2255}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1833 ( .a ({signal_2543, signal_2119}), .b ({signal_3224, signal_2191}), .c ({signal_3398, signal_2223}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1834 ( .a ({signal_2648, signal_2087}), .b ({signal_3154, signal_2159}), .c ({signal_3224, signal_2191}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1835 ( .a ({signal_2435, signal_1796}), .b ({signal_3399, signal_2224}), .c ({signal_3531, signal_2256}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1836 ( .a ({signal_2540, signal_2120}), .b ({signal_3225, signal_2192}), .c ({signal_3399, signal_2224}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1837 ( .a ({signal_2645, signal_2088}), .b ({signal_3155, signal_2160}), .c ({signal_3225, signal_2192}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1838 ( .a ({signal_2432, signal_1797}), .b ({signal_3400, signal_2225}), .c ({signal_3532, signal_2257}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1839 ( .a ({signal_2537, signal_2121}), .b ({signal_3226, signal_2193}), .c ({signal_3400, signal_2225}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1840 ( .a ({signal_2642, signal_2089}), .b ({signal_3156, signal_2161}), .c ({signal_3226, signal_2193}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1841 ( .a ({signal_2429, signal_2038}), .b ({signal_3166, signal_2306}), .c ({signal_3227, signal_2142}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1842 ( .a ({signal_2426, signal_2039}), .b ({signal_3167, signal_2307}), .c ({signal_3228, signal_2143}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1843 ( .a ({signal_2423, signal_2040}), .b ({signal_3168, signal_2308}), .c ({signal_3229, signal_2144}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1844 ( .a ({signal_2420, signal_2041}), .b ({signal_3169, signal_2309}), .c ({signal_3230, signal_2145}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1845 ( .a ({signal_2417, signal_2042}), .b ({signal_3170, signal_2310}), .c ({signal_3231, signal_2146}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1846 ( .a ({signal_2414, signal_2043}), .b ({signal_3171, signal_2311}), .c ({signal_3232, signal_2147}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1847 ( .a ({signal_2411, signal_2044}), .b ({signal_3172, signal_2312}), .c ({signal_3233, signal_2148}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1848 ( .a ({signal_2408, signal_2045}), .b ({signal_3173, signal_2313}), .c ({signal_3234, signal_2149}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1849 ( .a ({signal_2405, signal_1798}), .b ({signal_3401, signal_2226}), .c ({signal_3533, signal_2258}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1850 ( .a ({signal_2534, signal_2122}), .b ({signal_3235, signal_2194}), .c ({signal_3401, signal_2226}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1851 ( .a ({signal_2639, signal_2090}), .b ({signal_3157, signal_2162}), .c ({signal_3235, signal_2194}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1852 ( .a ({signal_2402, signal_2046}), .b ({signal_3086, signal_2314}), .c ({signal_3145, signal_2150}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1853 ( .a ({signal_2399, signal_2047}), .b ({signal_3087, signal_2315}), .c ({signal_3146, signal_2151}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1854 ( .a ({signal_2396, signal_2048}), .b ({signal_3088, signal_2316}), .c ({signal_3147, signal_2152}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1855 ( .a ({signal_2393, signal_2049}), .b ({signal_3089, signal_2317}), .c ({signal_3148, signal_2153}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1856 ( .a ({signal_2390, signal_2050}), .b ({signal_3090, signal_2318}), .c ({signal_3149, signal_2154}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1857 ( .a ({signal_2387, signal_2051}), .b ({signal_3091, signal_2319}), .c ({signal_3150, signal_2155}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1858 ( .a ({signal_2384, signal_2052}), .b ({signal_3092, signal_2320}), .c ({signal_3151, signal_2156}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1859 ( .a ({signal_2381, signal_2053}), .b ({signal_3093, signal_2321}), .c ({signal_3152, signal_2157}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1860 ( .a ({signal_2378, signal_2054}), .b ({signal_3094, signal_2322}), .c ({signal_3153, signal_2158}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1861 ( .a ({signal_2375, signal_2055}), .b ({signal_3095, signal_2323}), .c ({signal_3154, signal_2159}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1862 ( .a ({signal_2372, signal_1799}), .b ({signal_3402, signal_2227}), .c ({signal_3534, signal_2259}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1863 ( .a ({signal_2531, signal_2123}), .b ({signal_3236, signal_2195}), .c ({signal_3402, signal_2227}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1864 ( .a ({signal_2636, signal_2091}), .b ({signal_3158, signal_2163}), .c ({signal_3236, signal_2195}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1865 ( .a ({signal_2369, signal_2056}), .b ({signal_3096, signal_2324}), .c ({signal_3155, signal_2160}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1866 ( .a ({signal_2366, signal_2057}), .b ({signal_3097, signal_2325}), .c ({signal_3156, signal_2161}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1867 ( .a ({signal_2363, signal_2058}), .b ({signal_3098, signal_2326}), .c ({signal_3157, signal_2162}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1868 ( .a ({signal_2360, signal_2059}), .b ({signal_3099, signal_2327}), .c ({signal_3158, signal_2163}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1869 ( .a ({signal_2357, signal_2060}), .b ({signal_3100, signal_2328}), .c ({signal_3159, signal_2164}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1870 ( .a ({signal_2354, signal_2061}), .b ({signal_3101, signal_2329}), .c ({signal_3160, signal_2165}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1871 ( .a ({signal_2351, signal_2062}), .b ({signal_3102, signal_2330}), .c ({signal_3161, signal_2166}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1872 ( .a ({signal_2348, signal_2063}), .b ({signal_3103, signal_2331}), .c ({signal_3162, signal_2167}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1873 ( .a ({signal_2345, signal_2064}), .b ({signal_3104, signal_2332}), .c ({signal_3163, signal_2168}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1874 ( .a ({signal_2342, signal_2065}), .b ({signal_3105, signal_2333}), .c ({signal_3164, signal_2169}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1875 ( .a ({signal_2339, signal_1793}), .b ({signal_3403, signal_2237}), .c ({signal_3535, signal_2269}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1876 ( .a ({signal_2498, signal_2133}), .b ({signal_3237, signal_2205}), .c ({signal_3403, signal_2237}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1877 ( .a ({signal_2603, signal_2101}), .b ({signal_3165, signal_2173}), .c ({signal_3237, signal_2205}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1878 ( .a ({signal_2708, signal_2069}), .b ({signal_3109, signal_2337}), .c ({signal_3165, signal_2173}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1879 ( .a ({1'b0, signal_2134}), .b ({signal_3085, signal_2305}), .c ({signal_3166, signal_2306}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1880 ( .a ({1'b0, signal_2135}), .b ({signal_3081, signal_2298}), .c ({signal_3167, signal_2307}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1881 ( .a ({1'b0, signal_2136}), .b ({signal_3082, signal_2299}), .c ({signal_3168, signal_2308}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1882 ( .a ({1'b0, signal_2137}), .b ({signal_3083, signal_2300}), .c ({signal_3169, signal_2309}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1883 ( .a ({1'b0, signal_2138}), .b ({signal_3048, signal_1842}), .c ({signal_3170, signal_2310}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1884 ( .a ({1'b0, signal_2139}), .b ({signal_3049, signal_1843}), .c ({signal_3171, signal_2311}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1885 ( .a ({1'b0, signal_2140}), .b ({signal_3084, signal_2303}), .c ({signal_3172, signal_2312}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) cell_1886 ( .a ({1'b0, signal_2141}), .b ({signal_3050, signal_1845}), .c ({signal_3173, signal_2313}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1895 ( .s (signal_1489), .b ({signal_2339, signal_1793}), .a ({signal_3535, signal_2269}), .c ({signal_3640, signal_2037}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1896 ( .s (signal_1488), .b ({signal_2456, signal_1792}), .a ({signal_3524, signal_2268}), .c ({signal_3641, signal_2036}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1897 ( .s (signal_1487), .b ({signal_2489, signal_1791}), .a ({signal_3513, signal_2267}), .c ({signal_3642, signal_2035}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1898 ( .s (signal_1486), .b ({signal_2522, signal_1790}), .a ({signal_3510, signal_2266}), .c ({signal_3643, signal_2034}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1899 ( .s (signal_1485), .b ({signal_2555, signal_1789}), .a ({signal_3509, signal_2265}), .c ({signal_3644, signal_2033}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1900 ( .s (signal_1484), .b ({signal_2588, signal_1788}), .a ({signal_3508, signal_2264}), .c ({signal_3645, signal_2032}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1901 ( .s (signal_1488), .b ({signal_2621, signal_1787}), .a ({signal_3507, signal_2263}), .c ({signal_3646, signal_2031}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1902 ( .s (signal_1486), .b ({signal_2654, signal_1786}), .a ({signal_3506, signal_2262}), .c ({signal_3647, signal_2030}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1903 ( .s (signal_1489), .b ({signal_2687, signal_1801}), .a ({signal_3505, signal_2261}), .c ({signal_3648, signal_2029}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1904 ( .s (signal_1488), .b ({signal_2720, signal_1800}), .a ({signal_3504, signal_2260}), .c ({signal_3649, signal_2028}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1905 ( .s (signal_1487), .b ({signal_2372, signal_1799}), .a ({signal_3534, signal_2259}), .c ({signal_3650, signal_2027}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1906 ( .s (signal_1486), .b ({signal_2405, signal_1798}), .a ({signal_3533, signal_2258}), .c ({signal_3651, signal_2026}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1907 ( .s (signal_1485), .b ({signal_2432, signal_1797}), .a ({signal_3532, signal_2257}), .c ({signal_3652, signal_2025}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1908 ( .s (signal_1484), .b ({signal_2435, signal_1796}), .a ({signal_3531, signal_2256}), .c ({signal_3653, signal_2024}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1909 ( .s (signal_1485), .b ({signal_2438, signal_1795}), .a ({signal_3530, signal_2255}), .c ({signal_3654, signal_2023}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1910 ( .s (signal_1485), .b ({signal_2441, signal_1794}), .a ({signal_3529, signal_2254}), .c ({signal_3655, signal_2022}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1911 ( .s (signal_1489), .b ({signal_2444, signal_1809}), .a ({signal_3528, signal_2253}), .c ({signal_3656, signal_2021}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1912 ( .s (signal_1488), .b ({signal_2447, signal_1808}), .a ({signal_3527, signal_2252}), .c ({signal_3657, signal_2020}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1913 ( .s (signal_1487), .b ({signal_2450, signal_1807}), .a ({signal_3526, signal_2251}), .c ({signal_3658, signal_2019}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1914 ( .s (signal_1486), .b ({signal_2453, signal_1806}), .a ({signal_3525, signal_2250}), .c ({signal_3659, signal_2018}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1915 ( .s (signal_1484), .b ({signal_2459, signal_1805}), .a ({signal_3523, signal_2249}), .c ({signal_3660, signal_2017}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1916 ( .s (signal_1484), .b ({signal_2462, signal_1804}), .a ({signal_3522, signal_2248}), .c ({signal_3661, signal_2016}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1917 ( .s (signal_1489), .b ({signal_2465, signal_1803}), .a ({signal_3521, signal_2247}), .c ({signal_3662, signal_2015}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1918 ( .s (signal_1488), .b ({signal_2468, signal_1802}), .a ({signal_3520, signal_2246}), .c ({signal_3663, signal_2014}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1919 ( .s (signal_1487), .b ({signal_2471, signal_1785}), .a ({signal_3639, signal_2245}), .c ({signal_3736, signal_2013}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1920 ( .s (signal_1486), .b ({signal_2474, signal_1784}), .a ({signal_3638, signal_2244}), .c ({signal_3737, signal_2012}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1921 ( .s (signal_1485), .b ({signal_2477, signal_1783}), .a ({signal_3637, signal_2243}), .c ({signal_3738, signal_2011}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1922 ( .s (signal_1484), .b ({signal_2480, signal_1782}), .a ({signal_3636, signal_2242}), .c ({signal_3739, signal_2010}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1923 ( .s (signal_1489), .b ({signal_2483, signal_1781}), .a ({signal_3635, signal_2241}), .c ({signal_3740, signal_2009}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1924 ( .s (signal_1489), .b ({signal_2486, signal_1780}), .a ({signal_3634, signal_2240}), .c ({signal_3741, signal_2008}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1925 ( .s (signal_1488), .b ({signal_2492, signal_1779}), .a ({signal_3633, signal_2239}), .c ({signal_3742, signal_2007}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1926 ( .s (signal_1487), .b ({signal_2495, signal_1778}), .a ({signal_3632, signal_2238}), .c ({signal_3743, signal_2006}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1927 ( .s (signal_1488), .b ({signal_2498, signal_2133}), .a ({signal_3403, signal_2237}), .c ({signal_3536, signal_2005}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1928 ( .s (signal_1487), .b ({signal_2501, signal_2132}), .a ({signal_3392, signal_2236}), .c ({signal_3537, signal_2004}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1929 ( .s (signal_1486), .b ({signal_2504, signal_2131}), .a ({signal_3381, signal_2235}), .c ({signal_3538, signal_2003}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1930 ( .s (signal_1485), .b ({signal_2507, signal_2130}), .a ({signal_3378, signal_2234}), .c ({signal_3539, signal_2002}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1931 ( .s (signal_1484), .b ({signal_2510, signal_2129}), .a ({signal_3377, signal_2233}), .c ({signal_3540, signal_2001}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1932 ( .s (signal_1489), .b ({signal_2513, signal_2128}), .a ({signal_3376, signal_2232}), .c ({signal_3541, signal_2000}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1933 ( .s (signal_1488), .b ({signal_2516, signal_2127}), .a ({signal_3375, signal_2231}), .c ({signal_3542, signal_1999}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1934 ( .s (signal_1487), .b ({signal_2519, signal_2126}), .a ({signal_3374, signal_2230}), .c ({signal_3543, signal_1998}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1935 ( .s (signal_1486), .b ({signal_2525, signal_2125}), .a ({signal_3373, signal_2229}), .c ({signal_3544, signal_1997}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1936 ( .s (signal_1485), .b ({signal_2528, signal_2124}), .a ({signal_3372, signal_2228}), .c ({signal_3545, signal_1996}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1937 ( .s (signal_1484), .b ({signal_2531, signal_2123}), .a ({signal_3402, signal_2227}), .c ({signal_3546, signal_1995}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1938 ( .s (signal_1489), .b ({signal_2534, signal_2122}), .a ({signal_3401, signal_2226}), .c ({signal_3547, signal_1994}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1939 ( .s (signal_1484), .b ({signal_2537, signal_2121}), .a ({signal_3400, signal_2225}), .c ({signal_3548, signal_1993}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1940 ( .s (signal_1484), .b ({signal_2540, signal_2120}), .a ({signal_3399, signal_2224}), .c ({signal_3549, signal_1992}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1941 ( .s (signal_1484), .b ({signal_2543, signal_2119}), .a ({signal_3398, signal_2223}), .c ({signal_3550, signal_1991}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1942 ( .s (signal_1484), .b ({signal_2546, signal_2118}), .a ({signal_3397, signal_2222}), .c ({signal_3551, signal_1990}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1943 ( .s (signal_1484), .b ({signal_2549, signal_2117}), .a ({signal_3396, signal_2221}), .c ({signal_3552, signal_1989}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1944 ( .s (signal_1484), .b ({signal_2552, signal_2116}), .a ({signal_3395, signal_2220}), .c ({signal_3553, signal_1988}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1945 ( .s (signal_1484), .b ({signal_2558, signal_2115}), .a ({signal_3394, signal_2219}), .c ({signal_3554, signal_1987}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1946 ( .s (signal_1484), .b ({signal_2561, signal_2114}), .a ({signal_3393, signal_2218}), .c ({signal_3555, signal_1986}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1947 ( .s (signal_1484), .b ({signal_2564, signal_2113}), .a ({signal_3391, signal_2217}), .c ({signal_3556, signal_1985}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1948 ( .s (signal_1484), .b ({signal_2567, signal_2112}), .a ({signal_3390, signal_2216}), .c ({signal_3557, signal_1984}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1949 ( .s (signal_1484), .b ({signal_2570, signal_2111}), .a ({signal_3389, signal_2215}), .c ({signal_3558, signal_1983}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1950 ( .s (signal_1484), .b ({signal_2573, signal_2110}), .a ({signal_3388, signal_2214}), .c ({signal_3559, signal_1982}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1951 ( .s (signal_1485), .b ({signal_2576, signal_2109}), .a ({signal_3519, signal_2213}), .c ({signal_3664, signal_1981}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1952 ( .s (signal_1485), .b ({signal_2579, signal_2108}), .a ({signal_3518, signal_2212}), .c ({signal_3665, signal_1980}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1953 ( .s (signal_1485), .b ({signal_2582, signal_2107}), .a ({signal_3517, signal_2211}), .c ({signal_3666, signal_1979}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1954 ( .s (signal_1485), .b ({signal_2585, signal_2106}), .a ({signal_3516, signal_2210}), .c ({signal_3667, signal_1978}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1955 ( .s (signal_1485), .b ({signal_2591, signal_2105}), .a ({signal_3515, signal_2209}), .c ({signal_3668, signal_1977}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1956 ( .s (signal_1485), .b ({signal_2594, signal_2104}), .a ({signal_3514, signal_2208}), .c ({signal_3669, signal_1976}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1957 ( .s (signal_1485), .b ({signal_2597, signal_2103}), .a ({signal_3512, signal_2207}), .c ({signal_3670, signal_1975}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1958 ( .s (signal_1485), .b ({signal_2600, signal_2102}), .a ({signal_3511, signal_2206}), .c ({signal_3671, signal_1974}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1959 ( .s (signal_1485), .b ({signal_2603, signal_2101}), .a ({signal_3237, signal_2205}), .c ({signal_3404, signal_1973}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1960 ( .s (signal_1485), .b ({signal_2606, signal_2100}), .a ({signal_3218, signal_2204}), .c ({signal_3405, signal_1972}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1961 ( .s (signal_1485), .b ({signal_2609, signal_2099}), .a ({signal_3213, signal_2203}), .c ({signal_3406, signal_1971}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1962 ( .s (signal_1485), .b ({signal_2612, signal_2098}), .a ({signal_3212, signal_2202}), .c ({signal_3407, signal_1970}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1963 ( .s (signal_1486), .b ({signal_2615, signal_2097}), .a ({signal_3211, signal_2201}), .c ({signal_3408, signal_1969}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1964 ( .s (signal_1486), .b ({signal_2618, signal_2096}), .a ({signal_3210, signal_2200}), .c ({signal_3409, signal_1968}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1965 ( .s (signal_1486), .b ({signal_2624, signal_2095}), .a ({signal_3209, signal_2199}), .c ({signal_3410, signal_1967}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1966 ( .s (signal_1486), .b ({signal_2627, signal_2094}), .a ({signal_3208, signal_2198}), .c ({signal_3411, signal_1966}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1967 ( .s (signal_1486), .b ({signal_2630, signal_2093}), .a ({signal_3207, signal_2197}), .c ({signal_3412, signal_1965}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1968 ( .s (signal_1486), .b ({signal_2633, signal_2092}), .a ({signal_3206, signal_2196}), .c ({signal_3413, signal_1964}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1969 ( .s (signal_1486), .b ({signal_2636, signal_2091}), .a ({signal_3236, signal_2195}), .c ({signal_3414, signal_1963}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1970 ( .s (signal_1486), .b ({signal_2639, signal_2090}), .a ({signal_3235, signal_2194}), .c ({signal_3415, signal_1962}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1971 ( .s (signal_1486), .b ({signal_2642, signal_2089}), .a ({signal_3226, signal_2193}), .c ({signal_3416, signal_1961}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1972 ( .s (signal_1486), .b ({signal_2645, signal_2088}), .a ({signal_3225, signal_2192}), .c ({signal_3417, signal_1960}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1973 ( .s (signal_1486), .b ({signal_2648, signal_2087}), .a ({signal_3224, signal_2191}), .c ({signal_3418, signal_1959}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1974 ( .s (signal_1486), .b ({signal_2651, signal_2086}), .a ({signal_3223, signal_2190}), .c ({signal_3419, signal_1958}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1975 ( .s (signal_1487), .b ({signal_2657, signal_2085}), .a ({signal_3222, signal_2189}), .c ({signal_3420, signal_1957}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1976 ( .s (signal_1487), .b ({signal_2660, signal_2084}), .a ({signal_3221, signal_2188}), .c ({signal_3421, signal_1956}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1977 ( .s (signal_1487), .b ({signal_2663, signal_2083}), .a ({signal_3220, signal_2187}), .c ({signal_3422, signal_1955}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1978 ( .s (signal_1487), .b ({signal_2666, signal_2082}), .a ({signal_3219, signal_2186}), .c ({signal_3423, signal_1954}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1979 ( .s (signal_1487), .b ({signal_2669, signal_2081}), .a ({signal_3217, signal_2185}), .c ({signal_3424, signal_1953}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1980 ( .s (signal_1487), .b ({signal_2672, signal_2080}), .a ({signal_3216, signal_2184}), .c ({signal_3425, signal_1952}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1981 ( .s (signal_1487), .b ({signal_2675, signal_2079}), .a ({signal_3215, signal_2183}), .c ({signal_3426, signal_1951}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1982 ( .s (signal_1487), .b ({signal_2678, signal_2078}), .a ({signal_3214, signal_2182}), .c ({signal_3427, signal_1950}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1983 ( .s (signal_1487), .b ({signal_2681, signal_2077}), .a ({signal_3387, signal_2181}), .c ({signal_3560, signal_1949}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1984 ( .s (signal_1487), .b ({signal_2684, signal_2076}), .a ({signal_3386, signal_2180}), .c ({signal_3561, signal_1948}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1985 ( .s (signal_1487), .b ({signal_2690, signal_2075}), .a ({signal_3385, signal_2179}), .c ({signal_3562, signal_1947}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1986 ( .s (signal_1487), .b ({signal_2693, signal_2074}), .a ({signal_3384, signal_2178}), .c ({signal_3563, signal_1946}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1987 ( .s (signal_1488), .b ({signal_2696, signal_2073}), .a ({signal_3383, signal_2177}), .c ({signal_3564, signal_1945}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1988 ( .s (signal_1488), .b ({signal_2699, signal_2072}), .a ({signal_3382, signal_2176}), .c ({signal_3565, signal_1944}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1989 ( .s (signal_1488), .b ({signal_2702, signal_2071}), .a ({signal_3380, signal_2175}), .c ({signal_3566, signal_1943}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1990 ( .s (signal_1488), .b ({signal_2705, signal_2070}), .a ({signal_3379, signal_2174}), .c ({signal_3567, signal_1942}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1991 ( .s (signal_1488), .b ({signal_2708, signal_2069}), .a ({signal_3165, signal_2173}), .c ({signal_3238, signal_1941}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1992 ( .s (signal_1488), .b ({signal_2711, signal_2068}), .a ({signal_3144, signal_2172}), .c ({signal_3239, signal_1940}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1993 ( .s (signal_1488), .b ({signal_2714, signal_2067}), .a ({signal_3143, signal_2171}), .c ({signal_3240, signal_1939}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1994 ( .s (signal_1488), .b ({signal_2717, signal_2066}), .a ({signal_3142, signal_2170}), .c ({signal_3241, signal_1938}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1995 ( .s (signal_1488), .b ({signal_2342, signal_2065}), .a ({signal_3164, signal_2169}), .c ({signal_3242, signal_1937}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1996 ( .s (signal_1488), .b ({signal_2345, signal_2064}), .a ({signal_3163, signal_2168}), .c ({signal_3243, signal_1936}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1997 ( .s (signal_1488), .b ({signal_2348, signal_2063}), .a ({signal_3162, signal_2167}), .c ({signal_3244, signal_1935}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1998 ( .s (signal_1488), .b ({signal_2351, signal_2062}), .a ({signal_3161, signal_2166}), .c ({signal_3245, signal_1934}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1999 ( .s (signal_1489), .b ({signal_2354, signal_2061}), .a ({signal_3160, signal_2165}), .c ({signal_3246, signal_1933}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2000 ( .s (signal_1489), .b ({signal_2357, signal_2060}), .a ({signal_3159, signal_2164}), .c ({signal_3247, signal_1932}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2001 ( .s (signal_1489), .b ({signal_2360, signal_2059}), .a ({signal_3158, signal_2163}), .c ({signal_3248, signal_1931}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2002 ( .s (signal_1489), .b ({signal_2363, signal_2058}), .a ({signal_3157, signal_2162}), .c ({signal_3249, signal_1930}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2003 ( .s (signal_1489), .b ({signal_2366, signal_2057}), .a ({signal_3156, signal_2161}), .c ({signal_3250, signal_1929}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2004 ( .s (signal_1489), .b ({signal_2369, signal_2056}), .a ({signal_3155, signal_2160}), .c ({signal_3251, signal_1928}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2005 ( .s (signal_1489), .b ({signal_2375, signal_2055}), .a ({signal_3154, signal_2159}), .c ({signal_3252, signal_1927}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2006 ( .s (signal_1489), .b ({signal_2378, signal_2054}), .a ({signal_3153, signal_2158}), .c ({signal_3253, signal_1926}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2007 ( .s (signal_1489), .b ({signal_2381, signal_2053}), .a ({signal_3152, signal_2157}), .c ({signal_3254, signal_1925}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2008 ( .s (signal_1489), .b ({signal_2384, signal_2052}), .a ({signal_3151, signal_2156}), .c ({signal_3255, signal_1924}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2009 ( .s (signal_1489), .b ({signal_2387, signal_2051}), .a ({signal_3150, signal_2155}), .c ({signal_3256, signal_1923}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2010 ( .s (signal_1489), .b ({signal_2390, signal_2050}), .a ({signal_3149, signal_2154}), .c ({signal_3257, signal_1922}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2011 ( .s (signal_1490), .b ({signal_2393, signal_2049}), .a ({signal_3148, signal_2153}), .c ({signal_3258, signal_1921}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2012 ( .s (signal_1490), .b ({signal_2396, signal_2048}), .a ({signal_3147, signal_2152}), .c ({signal_3259, signal_1920}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2013 ( .s (signal_1490), .b ({signal_2399, signal_2047}), .a ({signal_3146, signal_2151}), .c ({signal_3260, signal_1919}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2014 ( .s (signal_1490), .b ({signal_2402, signal_2046}), .a ({signal_3145, signal_2150}), .c ({signal_3261, signal_1918}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2015 ( .s (signal_1490), .b ({signal_2408, signal_2045}), .a ({signal_3234, signal_2149}), .c ({signal_3428, signal_1917}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2016 ( .s (signal_1490), .b ({signal_2411, signal_2044}), .a ({signal_3233, signal_2148}), .c ({signal_3429, signal_1916}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2017 ( .s (signal_1490), .b ({signal_2414, signal_2043}), .a ({signal_3232, signal_2147}), .c ({signal_3430, signal_1915}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2018 ( .s (signal_1490), .b ({signal_2417, signal_2042}), .a ({signal_3231, signal_2146}), .c ({signal_3431, signal_1914}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2019 ( .s (signal_1490), .b ({signal_2420, signal_2041}), .a ({signal_3230, signal_2145}), .c ({signal_3432, signal_1913}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2020 ( .s (signal_1490), .b ({signal_2423, signal_2040}), .a ({signal_3229, signal_2144}), .c ({signal_3433, signal_1912}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2021 ( .s (signal_1490), .b ({signal_2426, signal_2039}), .a ({signal_3228, signal_2143}), .c ({signal_3434, signal_1911}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2022 ( .s (signal_1490), .b ({signal_2429, signal_2038}), .a ({signal_3227, signal_2142}), .c ({signal_3435, signal_1910}) ) ;
    AES_step2_ANF #(.low_latency(0), .pipeline(0)) cell_2061 ( .in0 ({signal_908, signal_788, signal_1841, signal_1840, signal_1839, signal_1837, signal_1836, signal_1835, signal_1834, signal_1833, signal_1832, signal_1831, signal_1829, signal_1828, signal_1827, signal_1826, signal_1825, signal_1824, signal_1823, signal_1821, signal_1820, signal_1819, signal_1818, signal_1817, signal_1816, signal_1815, signal_1813, signal_1812, signal_1811, signal_1810, signal_1148, signal_1028}), .in1 ({signal_3043, signal_3042, signal_2723, signal_2724, signal_2725, signal_2727, signal_2728, signal_2729, signal_2730, signal_2722, signal_2731, signal_2732, signal_2734, signal_2735, signal_2736, signal_2737, signal_2738, signal_2739, signal_2740, signal_2742, signal_2743, signal_2744, signal_2745, signal_2746, signal_2747, signal_2748, signal_2750, signal_2751, signal_2752, signal_2753, signal_3045, signal_3044}), .clk (clk), .r ({Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .out0 ({signal_2337, signal_2336, signal_2335, signal_2334, signal_2333, signal_2332, signal_2331, signal_2330, signal_2329, signal_2328, signal_2327, signal_2326, signal_2325, signal_2324, signal_2323, signal_2322, signal_2321, signal_2320, signal_2319, signal_2318, signal_2317, signal_2316, signal_2315, signal_2314, signal_2305, signal_2303, signal_2300, signal_2299, signal_2298, signal_1876, signal_1875, signal_1874, signal_1873, signal_1872, signal_1871, signal_1870, signal_1869, signal_1867, signal_1866, signal_1865, signal_1864, signal_1863, signal_1862, signal_1861, signal_1860, signal_1859, signal_1858, signal_1857, signal_1856, signal_1855, signal_1854, signal_1853, signal_1852, signal_1851, signal_1850, signal_1849, signal_1848, signal_1847, signal_1846, signal_1845, signal_1843, signal_1842, signal_1216, signal_1153}), .out1 ({signal_3109, signal_3108, signal_3107, signal_3106, signal_3105, signal_3104, signal_3103, signal_3102, signal_3101, signal_3100, signal_3099, signal_3098, signal_3097, signal_3096, signal_3095, signal_3094, signal_3093, signal_3092, signal_3091, signal_3090, signal_3089, signal_3088, signal_3087, signal_3086, signal_3085, signal_3084, signal_3083, signal_3082, signal_3081, signal_3080, signal_3079, signal_3078, signal_3077, signal_3076, signal_3075, signal_3074, signal_3073, signal_3072, signal_3071, signal_3070, signal_3069, signal_3068, signal_3067, signal_3066, signal_3065, signal_3064, signal_3063, signal_3062, signal_3061, signal_3060, signal_3059, signal_3058, signal_3057, signal_3056, signal_3055, signal_3054, signal_3053, signal_3052, signal_3051, signal_3050, signal_3049, signal_3048, signal_3047, signal_3046}) ) ;

    /* register cells */
    reg_masked #(.low_latency(0), .pipeline(0)) cell_159 ( .D ({signal_3437, signal_414}), .clk (signal_3792), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_162 ( .D ({signal_3263, signal_416}), .clk (signal_3792), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_165 ( .D ({signal_3265, signal_418}), .clk (signal_3792), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_168 ( .D ({signal_3267, signal_420}), .clk (signal_3792), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_171 ( .D ({signal_3269, signal_422}), .clk (signal_3792), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_174 ( .D ({signal_3271, signal_424}), .clk (signal_3792), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_177 ( .D ({signal_3273, signal_426}), .clk (signal_3792), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_180 ( .D ({signal_3275, signal_428}), .clk (signal_3792), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_183 ( .D ({signal_3277, signal_430}), .clk (signal_3792), .Q ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_186 ( .D ({signal_3439, signal_432}), .clk (signal_3792), .Q ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_189 ( .D ({signal_3279, signal_434}), .clk (signal_3792), .Q ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_192 ( .D ({signal_3281, signal_436}), .clk (signal_3792), .Q ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_195 ( .D ({signal_3283, signal_438}), .clk (signal_3792), .Q ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_198 ( .D ({signal_3285, signal_440}), .clk (signal_3792), .Q ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_201 ( .D ({signal_3287, signal_442}), .clk (signal_3792), .Q ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_204 ( .D ({signal_3289, signal_444}), .clk (signal_3792), .Q ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_207 ( .D ({signal_3291, signal_446}), .clk (signal_3792), .Q ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_210 ( .D ({signal_3293, signal_448}), .clk (signal_3792), .Q ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_213 ( .D ({signal_3295, signal_450}), .clk (signal_3792), .Q ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_216 ( .D ({signal_3297, signal_452}), .clk (signal_3792), .Q ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_219 ( .D ({signal_3299, signal_454}), .clk (signal_3792), .Q ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_222 ( .D ({signal_3301, signal_456}), .clk (signal_3792), .Q ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_225 ( .D ({signal_3303, signal_458}), .clk (signal_3792), .Q ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_228 ( .D ({signal_3305, signal_460}), .clk (signal_3792), .Q ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_231 ( .D ({signal_3307, signal_462}), .clk (signal_3792), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_234 ( .D ({signal_3309, signal_464}), .clk (signal_3792), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_237 ( .D ({signal_3311, signal_466}), .clk (signal_3792), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_240 ( .D ({signal_3313, signal_468}), .clk (signal_3792), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_243 ( .D ({signal_3315, signal_470}), .clk (signal_3792), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_246 ( .D ({signal_3317, signal_472}), .clk (signal_3792), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_249 ( .D ({signal_3319, signal_474}), .clk (signal_3792), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_252 ( .D ({signal_3321, signal_476}), .clk (signal_3792), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_255 ( .D ({signal_2851, signal_478}), .clk (signal_3792), .Q ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_258 ( .D ({signal_2853, signal_480}), .clk (signal_3792), .Q ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_261 ( .D ({signal_2855, signal_482}), .clk (signal_3792), .Q ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_264 ( .D ({signal_2857, signal_484}), .clk (signal_3792), .Q ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_267 ( .D ({signal_2859, signal_486}), .clk (signal_3792), .Q ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_270 ( .D ({signal_2861, signal_488}), .clk (signal_3792), .Q ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_273 ( .D ({signal_2863, signal_490}), .clk (signal_3792), .Q ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_276 ( .D ({signal_2865, signal_492}), .clk (signal_3792), .Q ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_279 ( .D ({signal_2867, signal_494}), .clk (signal_3792), .Q ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_282 ( .D ({signal_2869, signal_496}), .clk (signal_3792), .Q ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_285 ( .D ({signal_2871, signal_498}), .clk (signal_3792), .Q ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_288 ( .D ({signal_2873, signal_500}), .clk (signal_3792), .Q ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_291 ( .D ({signal_2875, signal_502}), .clk (signal_3792), .Q ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_294 ( .D ({signal_2877, signal_504}), .clk (signal_3792), .Q ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_297 ( .D ({signal_2879, signal_506}), .clk (signal_3792), .Q ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_300 ( .D ({signal_2881, signal_508}), .clk (signal_3792), .Q ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_303 ( .D ({signal_2883, signal_510}), .clk (signal_3792), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_306 ( .D ({signal_2885, signal_512}), .clk (signal_3792), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_309 ( .D ({signal_2887, signal_514}), .clk (signal_3792), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_312 ( .D ({signal_2889, signal_516}), .clk (signal_3792), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_315 ( .D ({signal_2891, signal_518}), .clk (signal_3792), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_318 ( .D ({signal_2893, signal_520}), .clk (signal_3792), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_321 ( .D ({signal_2895, signal_522}), .clk (signal_3792), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_324 ( .D ({signal_2897, signal_524}), .clk (signal_3792), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_327 ( .D ({signal_2899, signal_526}), .clk (signal_3792), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_330 ( .D ({signal_2901, signal_528}), .clk (signal_3792), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_333 ( .D ({signal_2903, signal_530}), .clk (signal_3792), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_336 ( .D ({signal_2905, signal_532}), .clk (signal_3792), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_339 ( .D ({signal_2907, signal_534}), .clk (signal_3792), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_342 ( .D ({signal_2909, signal_536}), .clk (signal_3792), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_345 ( .D ({signal_2911, signal_538}), .clk (signal_3792), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_348 ( .D ({signal_2913, signal_540}), .clk (signal_3792), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_351 ( .D ({signal_2915, signal_542}), .clk (signal_3792), .Q ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_354 ( .D ({signal_2917, signal_544}), .clk (signal_3792), .Q ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_357 ( .D ({signal_2919, signal_546}), .clk (signal_3792), .Q ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_360 ( .D ({signal_2921, signal_548}), .clk (signal_3792), .Q ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_363 ( .D ({signal_2923, signal_550}), .clk (signal_3792), .Q ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_366 ( .D ({signal_2925, signal_552}), .clk (signal_3792), .Q ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_369 ( .D ({signal_2927, signal_554}), .clk (signal_3792), .Q ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_372 ( .D ({signal_2929, signal_556}), .clk (signal_3792), .Q ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_375 ( .D ({signal_2931, signal_558}), .clk (signal_3792), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_378 ( .D ({signal_2933, signal_560}), .clk (signal_3792), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_381 ( .D ({signal_2935, signal_562}), .clk (signal_3792), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_384 ( .D ({signal_2937, signal_564}), .clk (signal_3792), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_387 ( .D ({signal_2939, signal_566}), .clk (signal_3792), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_390 ( .D ({signal_2941, signal_568}), .clk (signal_3792), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_393 ( .D ({signal_2943, signal_570}), .clk (signal_3792), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_396 ( .D ({signal_2945, signal_572}), .clk (signal_3792), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_399 ( .D ({signal_2947, signal_574}), .clk (signal_3792), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_402 ( .D ({signal_2949, signal_576}), .clk (signal_3792), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_405 ( .D ({signal_2951, signal_578}), .clk (signal_3792), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_408 ( .D ({signal_2953, signal_580}), .clk (signal_3792), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_411 ( .D ({signal_2955, signal_582}), .clk (signal_3792), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_414 ( .D ({signal_2957, signal_584}), .clk (signal_3792), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_417 ( .D ({signal_2959, signal_586}), .clk (signal_3792), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_420 ( .D ({signal_2961, signal_588}), .clk (signal_3792), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_423 ( .D ({signal_2963, signal_590}), .clk (signal_3792), .Q ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_426 ( .D ({signal_2965, signal_592}), .clk (signal_3792), .Q ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_429 ( .D ({signal_2967, signal_594}), .clk (signal_3792), .Q ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_432 ( .D ({signal_2969, signal_596}), .clk (signal_3792), .Q ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_435 ( .D ({signal_2971, signal_598}), .clk (signal_3792), .Q ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_438 ( .D ({signal_2973, signal_600}), .clk (signal_3792), .Q ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_441 ( .D ({signal_2975, signal_602}), .clk (signal_3792), .Q ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_444 ( .D ({signal_2977, signal_604}), .clk (signal_3792), .Q ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_447 ( .D ({signal_2979, signal_606}), .clk (signal_3792), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_450 ( .D ({signal_2981, signal_608}), .clk (signal_3792), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_453 ( .D ({signal_2983, signal_610}), .clk (signal_3792), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_456 ( .D ({signal_2985, signal_612}), .clk (signal_3792), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_459 ( .D ({signal_2987, signal_614}), .clk (signal_3792), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_462 ( .D ({signal_2989, signal_616}), .clk (signal_3792), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_465 ( .D ({signal_2991, signal_618}), .clk (signal_3792), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_468 ( .D ({signal_2993, signal_620}), .clk (signal_3792), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_471 ( .D ({signal_2995, signal_622}), .clk (signal_3792), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_474 ( .D ({signal_2997, signal_624}), .clk (signal_3792), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_477 ( .D ({signal_2999, signal_626}), .clk (signal_3792), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_480 ( .D ({signal_3001, signal_628}), .clk (signal_3792), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_483 ( .D ({signal_3003, signal_630}), .clk (signal_3792), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_486 ( .D ({signal_3005, signal_632}), .clk (signal_3792), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_489 ( .D ({signal_3007, signal_634}), .clk (signal_3792), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_492 ( .D ({signal_3009, signal_636}), .clk (signal_3792), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_495 ( .D ({signal_3011, signal_638}), .clk (signal_3792), .Q ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_498 ( .D ({signal_3013, signal_640}), .clk (signal_3792), .Q ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_501 ( .D ({signal_3015, signal_642}), .clk (signal_3792), .Q ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_504 ( .D ({signal_3017, signal_644}), .clk (signal_3792), .Q ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_507 ( .D ({signal_3019, signal_646}), .clk (signal_3792), .Q ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_510 ( .D ({signal_3021, signal_648}), .clk (signal_3792), .Q ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_513 ( .D ({signal_3023, signal_650}), .clk (signal_3792), .Q ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_516 ( .D ({signal_3025, signal_652}), .clk (signal_3792), .Q ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_519 ( .D ({signal_3027, signal_654}), .clk (signal_3792), .Q ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_522 ( .D ({signal_3029, signal_656}), .clk (signal_3792), .Q ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_525 ( .D ({signal_3031, signal_658}), .clk (signal_3792), .Q ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_528 ( .D ({signal_3033, signal_660}), .clk (signal_3792), .Q ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_531 ( .D ({signal_3035, signal_662}), .clk (signal_3792), .Q ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_534 ( .D ({signal_3037, signal_664}), .clk (signal_3792), .Q ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_537 ( .D ({signal_3039, signal_666}), .clk (signal_3792), .Q ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_540 ( .D ({signal_3041, signal_668}), .clk (signal_3792), .Q ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1368 ( .D ({signal_3673, signal_1227}), .clk (signal_3792), .Q ({signal_2339, signal_1793}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1371 ( .D ({signal_3675, signal_1229}), .clk (signal_3792), .Q ({signal_2456, signal_1792}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1374 ( .D ({signal_3677, signal_1231}), .clk (signal_3792), .Q ({signal_2489, signal_1791}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1377 ( .D ({signal_3679, signal_1233}), .clk (signal_3792), .Q ({signal_2522, signal_1790}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1380 ( .D ({signal_3681, signal_1235}), .clk (signal_3792), .Q ({signal_2555, signal_1789}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1383 ( .D ({signal_3683, signal_1237}), .clk (signal_3792), .Q ({signal_2588, signal_1788}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1386 ( .D ({signal_3685, signal_1239}), .clk (signal_3792), .Q ({signal_2621, signal_1787}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1389 ( .D ({signal_3687, signal_1241}), .clk (signal_3792), .Q ({signal_2654, signal_1786}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1392 ( .D ({signal_3689, signal_1243}), .clk (signal_3792), .Q ({signal_2687, signal_1801}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1395 ( .D ({signal_3691, signal_1245}), .clk (signal_3792), .Q ({signal_2720, signal_1800}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1398 ( .D ({signal_3693, signal_1247}), .clk (signal_3792), .Q ({signal_2372, signal_1799}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1401 ( .D ({signal_3695, signal_1249}), .clk (signal_3792), .Q ({signal_2405, signal_1798}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1404 ( .D ({signal_3697, signal_1251}), .clk (signal_3792), .Q ({signal_2432, signal_1797}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1407 ( .D ({signal_3699, signal_1253}), .clk (signal_3792), .Q ({signal_2435, signal_1796}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1410 ( .D ({signal_3701, signal_1255}), .clk (signal_3792), .Q ({signal_2438, signal_1795}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1413 ( .D ({signal_3703, signal_1257}), .clk (signal_3792), .Q ({signal_2441, signal_1794}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1416 ( .D ({signal_3705, signal_1259}), .clk (signal_3792), .Q ({signal_2444, signal_1809}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1419 ( .D ({signal_3707, signal_1261}), .clk (signal_3792), .Q ({signal_2447, signal_1808}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1422 ( .D ({signal_3709, signal_1263}), .clk (signal_3792), .Q ({signal_2450, signal_1807}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1425 ( .D ({signal_3711, signal_1265}), .clk (signal_3792), .Q ({signal_2453, signal_1806}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1428 ( .D ({signal_3713, signal_1267}), .clk (signal_3792), .Q ({signal_2459, signal_1805}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1431 ( .D ({signal_3715, signal_1269}), .clk (signal_3792), .Q ({signal_2462, signal_1804}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1434 ( .D ({signal_3717, signal_1271}), .clk (signal_3792), .Q ({signal_2465, signal_1803}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1437 ( .D ({signal_3719, signal_1273}), .clk (signal_3792), .Q ({signal_2468, signal_1802}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1440 ( .D ({signal_3745, signal_1275}), .clk (signal_3792), .Q ({signal_2471, signal_1785}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1443 ( .D ({signal_3747, signal_1277}), .clk (signal_3792), .Q ({signal_2474, signal_1784}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1446 ( .D ({signal_3749, signal_1279}), .clk (signal_3792), .Q ({signal_2477, signal_1783}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1449 ( .D ({signal_3751, signal_1281}), .clk (signal_3792), .Q ({signal_2480, signal_1782}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1452 ( .D ({signal_3753, signal_1283}), .clk (signal_3792), .Q ({signal_2483, signal_1781}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1455 ( .D ({signal_3755, signal_1285}), .clk (signal_3792), .Q ({signal_2486, signal_1780}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1458 ( .D ({signal_3757, signal_1287}), .clk (signal_3792), .Q ({signal_2492, signal_1779}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1461 ( .D ({signal_3759, signal_1289}), .clk (signal_3792), .Q ({signal_2495, signal_1778}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1464 ( .D ({signal_3569, signal_1291}), .clk (signal_3792), .Q ({signal_2498, signal_2133}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1467 ( .D ({signal_3571, signal_1293}), .clk (signal_3792), .Q ({signal_2501, signal_2132}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1470 ( .D ({signal_3573, signal_1295}), .clk (signal_3792), .Q ({signal_2504, signal_2131}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1473 ( .D ({signal_3575, signal_1297}), .clk (signal_3792), .Q ({signal_2507, signal_2130}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1476 ( .D ({signal_3577, signal_1299}), .clk (signal_3792), .Q ({signal_2510, signal_2129}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1479 ( .D ({signal_3579, signal_1301}), .clk (signal_3792), .Q ({signal_2513, signal_2128}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1482 ( .D ({signal_3581, signal_1303}), .clk (signal_3792), .Q ({signal_2516, signal_2127}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1485 ( .D ({signal_3583, signal_1305}), .clk (signal_3792), .Q ({signal_2519, signal_2126}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1488 ( .D ({signal_3585, signal_1307}), .clk (signal_3792), .Q ({signal_2525, signal_2125}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1491 ( .D ({signal_3587, signal_1309}), .clk (signal_3792), .Q ({signal_2528, signal_2124}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1494 ( .D ({signal_3589, signal_1311}), .clk (signal_3792), .Q ({signal_2531, signal_2123}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1497 ( .D ({signal_3591, signal_1313}), .clk (signal_3792), .Q ({signal_2534, signal_2122}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1500 ( .D ({signal_3593, signal_1315}), .clk (signal_3792), .Q ({signal_2537, signal_2121}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1503 ( .D ({signal_3595, signal_1317}), .clk (signal_3792), .Q ({signal_2540, signal_2120}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1506 ( .D ({signal_3597, signal_1319}), .clk (signal_3792), .Q ({signal_2543, signal_2119}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1509 ( .D ({signal_3599, signal_1321}), .clk (signal_3792), .Q ({signal_2546, signal_2118}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1512 ( .D ({signal_3601, signal_1323}), .clk (signal_3792), .Q ({signal_2549, signal_2117}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1515 ( .D ({signal_3603, signal_1325}), .clk (signal_3792), .Q ({signal_2552, signal_2116}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1518 ( .D ({signal_3605, signal_1327}), .clk (signal_3792), .Q ({signal_2558, signal_2115}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1521 ( .D ({signal_3607, signal_1329}), .clk (signal_3792), .Q ({signal_2561, signal_2114}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1524 ( .D ({signal_3609, signal_1331}), .clk (signal_3792), .Q ({signal_2564, signal_2113}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1527 ( .D ({signal_3611, signal_1333}), .clk (signal_3792), .Q ({signal_2567, signal_2112}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1530 ( .D ({signal_3613, signal_1335}), .clk (signal_3792), .Q ({signal_2570, signal_2111}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1533 ( .D ({signal_3615, signal_1337}), .clk (signal_3792), .Q ({signal_2573, signal_2110}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1536 ( .D ({signal_3721, signal_1339}), .clk (signal_3792), .Q ({signal_2576, signal_2109}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1539 ( .D ({signal_3723, signal_1341}), .clk (signal_3792), .Q ({signal_2579, signal_2108}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1542 ( .D ({signal_3725, signal_1343}), .clk (signal_3792), .Q ({signal_2582, signal_2107}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1545 ( .D ({signal_3727, signal_1345}), .clk (signal_3792), .Q ({signal_2585, signal_2106}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1548 ( .D ({signal_3729, signal_1347}), .clk (signal_3792), .Q ({signal_2591, signal_2105}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1551 ( .D ({signal_3731, signal_1349}), .clk (signal_3792), .Q ({signal_2594, signal_2104}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1554 ( .D ({signal_3733, signal_1351}), .clk (signal_3792), .Q ({signal_2597, signal_2103}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1557 ( .D ({signal_3735, signal_1353}), .clk (signal_3792), .Q ({signal_2600, signal_2102}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1560 ( .D ({signal_3441, signal_1355}), .clk (signal_3792), .Q ({signal_2603, signal_2101}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1563 ( .D ({signal_3443, signal_1357}), .clk (signal_3792), .Q ({signal_2606, signal_2100}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1566 ( .D ({signal_3445, signal_1359}), .clk (signal_3792), .Q ({signal_2609, signal_2099}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1569 ( .D ({signal_3447, signal_1361}), .clk (signal_3792), .Q ({signal_2612, signal_2098}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1572 ( .D ({signal_3449, signal_1363}), .clk (signal_3792), .Q ({signal_2615, signal_2097}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1575 ( .D ({signal_3451, signal_1365}), .clk (signal_3792), .Q ({signal_2618, signal_2096}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1578 ( .D ({signal_3453, signal_1367}), .clk (signal_3792), .Q ({signal_2624, signal_2095}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1581 ( .D ({signal_3455, signal_1369}), .clk (signal_3792), .Q ({signal_2627, signal_2094}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1584 ( .D ({signal_3457, signal_1371}), .clk (signal_3792), .Q ({signal_2630, signal_2093}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1587 ( .D ({signal_3459, signal_1373}), .clk (signal_3792), .Q ({signal_2633, signal_2092}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1590 ( .D ({signal_3461, signal_1375}), .clk (signal_3792), .Q ({signal_2636, signal_2091}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1593 ( .D ({signal_3463, signal_1377}), .clk (signal_3792), .Q ({signal_2639, signal_2090}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1596 ( .D ({signal_3465, signal_1379}), .clk (signal_3792), .Q ({signal_2642, signal_2089}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1599 ( .D ({signal_3467, signal_1381}), .clk (signal_3792), .Q ({signal_2645, signal_2088}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1602 ( .D ({signal_3469, signal_1383}), .clk (signal_3792), .Q ({signal_2648, signal_2087}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1605 ( .D ({signal_3471, signal_1385}), .clk (signal_3792), .Q ({signal_2651, signal_2086}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1608 ( .D ({signal_3473, signal_1387}), .clk (signal_3792), .Q ({signal_2657, signal_2085}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1611 ( .D ({signal_3475, signal_1389}), .clk (signal_3792), .Q ({signal_2660, signal_2084}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1614 ( .D ({signal_3477, signal_1391}), .clk (signal_3792), .Q ({signal_2663, signal_2083}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1617 ( .D ({signal_3479, signal_1393}), .clk (signal_3792), .Q ({signal_2666, signal_2082}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1620 ( .D ({signal_3481, signal_1395}), .clk (signal_3792), .Q ({signal_2669, signal_2081}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1623 ( .D ({signal_3483, signal_1397}), .clk (signal_3792), .Q ({signal_2672, signal_2080}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1626 ( .D ({signal_3485, signal_1399}), .clk (signal_3792), .Q ({signal_2675, signal_2079}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1629 ( .D ({signal_3487, signal_1401}), .clk (signal_3792), .Q ({signal_2678, signal_2078}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1632 ( .D ({signal_3617, signal_1403}), .clk (signal_3792), .Q ({signal_2681, signal_2077}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1635 ( .D ({signal_3619, signal_1405}), .clk (signal_3792), .Q ({signal_2684, signal_2076}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1638 ( .D ({signal_3621, signal_1407}), .clk (signal_3792), .Q ({signal_2690, signal_2075}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1641 ( .D ({signal_3623, signal_1409}), .clk (signal_3792), .Q ({signal_2693, signal_2074}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1644 ( .D ({signal_3625, signal_1411}), .clk (signal_3792), .Q ({signal_2696, signal_2073}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1647 ( .D ({signal_3627, signal_1413}), .clk (signal_3792), .Q ({signal_2699, signal_2072}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1650 ( .D ({signal_3629, signal_1415}), .clk (signal_3792), .Q ({signal_2702, signal_2071}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1653 ( .D ({signal_3631, signal_1417}), .clk (signal_3792), .Q ({signal_2705, signal_2070}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1656 ( .D ({signal_3325, signal_1419}), .clk (signal_3792), .Q ({signal_2708, signal_2069}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1659 ( .D ({signal_3327, signal_1421}), .clk (signal_3792), .Q ({signal_2711, signal_2068}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1662 ( .D ({signal_3329, signal_1423}), .clk (signal_3792), .Q ({signal_2714, signal_2067}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1665 ( .D ({signal_3331, signal_1425}), .clk (signal_3792), .Q ({signal_2717, signal_2066}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1668 ( .D ({signal_3333, signal_1427}), .clk (signal_3792), .Q ({signal_2342, signal_2065}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1671 ( .D ({signal_3335, signal_1429}), .clk (signal_3792), .Q ({signal_2345, signal_2064}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1674 ( .D ({signal_3337, signal_1431}), .clk (signal_3792), .Q ({signal_2348, signal_2063}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1677 ( .D ({signal_3339, signal_1433}), .clk (signal_3792), .Q ({signal_2351, signal_2062}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1680 ( .D ({signal_3341, signal_1435}), .clk (signal_3792), .Q ({signal_2354, signal_2061}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1683 ( .D ({signal_3343, signal_1437}), .clk (signal_3792), .Q ({signal_2357, signal_2060}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1686 ( .D ({signal_3345, signal_1439}), .clk (signal_3792), .Q ({signal_2360, signal_2059}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1689 ( .D ({signal_3347, signal_1441}), .clk (signal_3792), .Q ({signal_2363, signal_2058}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1692 ( .D ({signal_3349, signal_1443}), .clk (signal_3792), .Q ({signal_2366, signal_2057}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1695 ( .D ({signal_3351, signal_1445}), .clk (signal_3792), .Q ({signal_2369, signal_2056}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1698 ( .D ({signal_3353, signal_1447}), .clk (signal_3792), .Q ({signal_2375, signal_2055}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1701 ( .D ({signal_3355, signal_1449}), .clk (signal_3792), .Q ({signal_2378, signal_2054}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1704 ( .D ({signal_3357, signal_1451}), .clk (signal_3792), .Q ({signal_2381, signal_2053}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1707 ( .D ({signal_3359, signal_1453}), .clk (signal_3792), .Q ({signal_2384, signal_2052}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1710 ( .D ({signal_3361, signal_1455}), .clk (signal_3792), .Q ({signal_2387, signal_2051}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1713 ( .D ({signal_3363, signal_1457}), .clk (signal_3792), .Q ({signal_2390, signal_2050}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1716 ( .D ({signal_3365, signal_1459}), .clk (signal_3792), .Q ({signal_2393, signal_2049}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1719 ( .D ({signal_3367, signal_1461}), .clk (signal_3792), .Q ({signal_2396, signal_2048}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1722 ( .D ({signal_3369, signal_1463}), .clk (signal_3792), .Q ({signal_2399, signal_2047}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1725 ( .D ({signal_3371, signal_1465}), .clk (signal_3792), .Q ({signal_2402, signal_2046}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1728 ( .D ({signal_3489, signal_1467}), .clk (signal_3792), .Q ({signal_2408, signal_2045}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1731 ( .D ({signal_3491, signal_1469}), .clk (signal_3792), .Q ({signal_2411, signal_2044}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1734 ( .D ({signal_3493, signal_1471}), .clk (signal_3792), .Q ({signal_2414, signal_2043}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1737 ( .D ({signal_3495, signal_1473}), .clk (signal_3792), .Q ({signal_2417, signal_2042}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1740 ( .D ({signal_3497, signal_1475}), .clk (signal_3792), .Q ({signal_2420, signal_2041}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1743 ( .D ({signal_3499, signal_1477}), .clk (signal_3792), .Q ({signal_2423, signal_2040}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1746 ( .D ({signal_3501, signal_1479}), .clk (signal_3792), .Q ({signal_2426, signal_2039}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_1749 ( .D ({signal_3503, signal_1481}), .clk (signal_3792), .Q ({signal_2429, signal_2038}) ) ;
    DFF_X1 cell_2035 ( .D (signal_1502), .CK (signal_3792), .Q (signal_2273), .QN () ) ;
    DFF_X1 cell_2037 ( .D (signal_1501), .CK (signal_3792), .Q (signal_2272), .QN () ) ;
    DFF_X1 cell_2039 ( .D (signal_1499), .CK (signal_3792), .Q (signal_2271), .QN () ) ;
    DFF_X1 cell_2041 ( .D (signal_1498), .CK (signal_3792), .Q (signal_2270), .QN () ) ;
    DFF_X1 cell_2056 ( .D (signal_1520), .CK (signal_3792), .Q (signal_2276), .QN () ) ;
    DFF_X1 cell_2058 ( .D (signal_1519), .CK (signal_3792), .Q (signal_2275), .QN () ) ;
    DFF_X1 cell_2060 ( .D (signal_1518), .CK (signal_3792), .Q (signal_2274), .QN () ) ;
endmodule
