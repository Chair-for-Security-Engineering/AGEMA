/* modified netlist. Source: module sbox in file Designs/AESSbox//lookup/AGEMA/sbox.v */
/* 34 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 35 register stage(s) in total */

module sbox_HPC2_Pipeline_d2 (SI_s0, clk, SI_s1, SI_s2, Fresh, SO_s0, SO_s1, SO_s2);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input [7:0] SI_s2 ;
    input [2603:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    output [7:0] SO_s2 ;
    wire N169 ;
    wire N277 ;
    wire N379 ;
    wire N470 ;
    wire N563 ;
    wire N639 ;
    wire N723 ;
    wire N789 ;
    wire n1922 ;
    wire n1923 ;
    wire n1924 ;
    wire n1925 ;
    wire n1926 ;
    wire n1927 ;
    wire n1928 ;
    wire n1929 ;
    wire n1930 ;
    wire n1931 ;
    wire n1932 ;
    wire n1933 ;
    wire n1934 ;
    wire n1935 ;
    wire n1936 ;
    wire n1937 ;
    wire n1938 ;
    wire n1939 ;
    wire n1940 ;
    wire n1941 ;
    wire n1942 ;
    wire n1943 ;
    wire n1944 ;
    wire n1945 ;
    wire n1946 ;
    wire n1947 ;
    wire n1948 ;
    wire n1949 ;
    wire n1950 ;
    wire n1951 ;
    wire n1952 ;
    wire n1953 ;
    wire n1954 ;
    wire n1955 ;
    wire n1956 ;
    wire n1957 ;
    wire n1958 ;
    wire n1959 ;
    wire n1960 ;
    wire n1961 ;
    wire n1962 ;
    wire n1963 ;
    wire n1964 ;
    wire n1965 ;
    wire n1966 ;
    wire n1967 ;
    wire n1968 ;
    wire n1969 ;
    wire n1970 ;
    wire n1971 ;
    wire n1972 ;
    wire n1973 ;
    wire n1974 ;
    wire n1975 ;
    wire n1976 ;
    wire n1977 ;
    wire n1978 ;
    wire n1979 ;
    wire n1980 ;
    wire n1981 ;
    wire n1982 ;
    wire n1983 ;
    wire n1984 ;
    wire n1985 ;
    wire n1986 ;
    wire n1987 ;
    wire n1988 ;
    wire n1989 ;
    wire n1990 ;
    wire n1991 ;
    wire n1992 ;
    wire n1993 ;
    wire n1994 ;
    wire n1995 ;
    wire n1996 ;
    wire n1997 ;
    wire n1998 ;
    wire n1999 ;
    wire n2000 ;
    wire n2001 ;
    wire n2002 ;
    wire n2003 ;
    wire n2004 ;
    wire n2005 ;
    wire n2006 ;
    wire n2007 ;
    wire n2008 ;
    wire n2009 ;
    wire n2010 ;
    wire n2011 ;
    wire n2012 ;
    wire n2013 ;
    wire n2014 ;
    wire n2015 ;
    wire n2016 ;
    wire n2017 ;
    wire n2018 ;
    wire n2019 ;
    wire n2020 ;
    wire n2021 ;
    wire n2022 ;
    wire n2023 ;
    wire n2024 ;
    wire n2025 ;
    wire n2026 ;
    wire n2027 ;
    wire n2028 ;
    wire n2029 ;
    wire n2030 ;
    wire n2031 ;
    wire n2032 ;
    wire n2033 ;
    wire n2034 ;
    wire n2035 ;
    wire n2036 ;
    wire n2037 ;
    wire n2038 ;
    wire n2039 ;
    wire n2040 ;
    wire n2041 ;
    wire n2042 ;
    wire n2043 ;
    wire n2044 ;
    wire n2045 ;
    wire n2046 ;
    wire n2047 ;
    wire n2048 ;
    wire n2049 ;
    wire n2050 ;
    wire n2051 ;
    wire n2052 ;
    wire n2053 ;
    wire n2054 ;
    wire n2055 ;
    wire n2056 ;
    wire n2057 ;
    wire n2058 ;
    wire n2059 ;
    wire n2060 ;
    wire n2061 ;
    wire n2062 ;
    wire n2063 ;
    wire n2064 ;
    wire n2065 ;
    wire n2066 ;
    wire n2067 ;
    wire n2068 ;
    wire n2069 ;
    wire n2070 ;
    wire n2071 ;
    wire n2072 ;
    wire n2073 ;
    wire n2074 ;
    wire n2075 ;
    wire n2076 ;
    wire n2077 ;
    wire n2078 ;
    wire n2079 ;
    wire n2080 ;
    wire n2081 ;
    wire n2082 ;
    wire n2083 ;
    wire n2084 ;
    wire n2085 ;
    wire n2086 ;
    wire n2087 ;
    wire n2088 ;
    wire n2089 ;
    wire n2090 ;
    wire n2091 ;
    wire n2092 ;
    wire n2093 ;
    wire n2094 ;
    wire n2095 ;
    wire n2096 ;
    wire n2097 ;
    wire n2098 ;
    wire n2099 ;
    wire n2100 ;
    wire n2101 ;
    wire n2102 ;
    wire n2103 ;
    wire n2104 ;
    wire n2105 ;
    wire n2106 ;
    wire n2107 ;
    wire n2108 ;
    wire n2109 ;
    wire n2110 ;
    wire n2111 ;
    wire n2112 ;
    wire n2113 ;
    wire n2114 ;
    wire n2115 ;
    wire n2116 ;
    wire n2117 ;
    wire n2118 ;
    wire n2119 ;
    wire n2120 ;
    wire n2121 ;
    wire n2122 ;
    wire n2123 ;
    wire n2124 ;
    wire n2125 ;
    wire n2126 ;
    wire n2127 ;
    wire n2128 ;
    wire n2129 ;
    wire n2130 ;
    wire n2131 ;
    wire n2132 ;
    wire n2133 ;
    wire n2134 ;
    wire n2135 ;
    wire n2136 ;
    wire n2137 ;
    wire n2138 ;
    wire n2139 ;
    wire n2140 ;
    wire n2141 ;
    wire n2142 ;
    wire n2143 ;
    wire n2144 ;
    wire n2145 ;
    wire n2146 ;
    wire n2147 ;
    wire n2148 ;
    wire n2149 ;
    wire n2150 ;
    wire n2151 ;
    wire n2152 ;
    wire n2153 ;
    wire n2154 ;
    wire n2155 ;
    wire n2156 ;
    wire n2157 ;
    wire n2158 ;
    wire n2159 ;
    wire n2160 ;
    wire n2161 ;
    wire n2162 ;
    wire n2163 ;
    wire n2164 ;
    wire n2165 ;
    wire n2166 ;
    wire n2167 ;
    wire n2168 ;
    wire n2169 ;
    wire n2170 ;
    wire n2171 ;
    wire n2172 ;
    wire n2173 ;
    wire n2174 ;
    wire n2175 ;
    wire n2176 ;
    wire n2177 ;
    wire n2178 ;
    wire n2179 ;
    wire n2180 ;
    wire n2181 ;
    wire n2182 ;
    wire n2183 ;
    wire n2184 ;
    wire n2185 ;
    wire n2186 ;
    wire n2187 ;
    wire n2188 ;
    wire n2189 ;
    wire n2190 ;
    wire n2191 ;
    wire n2192 ;
    wire n2193 ;
    wire n2194 ;
    wire n2195 ;
    wire n2196 ;
    wire n2197 ;
    wire n2198 ;
    wire n2199 ;
    wire n2200 ;
    wire n2201 ;
    wire n2202 ;
    wire n2203 ;
    wire n2204 ;
    wire n2205 ;
    wire n2206 ;
    wire n2207 ;
    wire n2208 ;
    wire n2209 ;
    wire n2210 ;
    wire n2211 ;
    wire n2212 ;
    wire n2213 ;
    wire n2214 ;
    wire n2215 ;
    wire n2216 ;
    wire n2217 ;
    wire n2218 ;
    wire n2219 ;
    wire n2220 ;
    wire n2221 ;
    wire n2222 ;
    wire n2223 ;
    wire n2224 ;
    wire n2225 ;
    wire n2226 ;
    wire n2227 ;
    wire n2228 ;
    wire n2229 ;
    wire n2230 ;
    wire n2231 ;
    wire n2232 ;
    wire n2233 ;
    wire n2234 ;
    wire n2235 ;
    wire n2236 ;
    wire n2237 ;
    wire n2238 ;
    wire n2239 ;
    wire n2240 ;
    wire n2241 ;
    wire n2242 ;
    wire n2243 ;
    wire n2244 ;
    wire n2245 ;
    wire n2246 ;
    wire n2247 ;
    wire n2248 ;
    wire n2249 ;
    wire n2250 ;
    wire n2251 ;
    wire n2252 ;
    wire n2253 ;
    wire n2254 ;
    wire n2255 ;
    wire n2256 ;
    wire n2257 ;
    wire n2258 ;
    wire n2259 ;
    wire n2260 ;
    wire n2261 ;
    wire n2262 ;
    wire n2263 ;
    wire n2264 ;
    wire n2265 ;
    wire n2266 ;
    wire n2267 ;
    wire n2268 ;
    wire n2269 ;
    wire n2270 ;
    wire n2271 ;
    wire n2272 ;
    wire n2273 ;
    wire n2274 ;
    wire n2275 ;
    wire n2276 ;
    wire n2277 ;
    wire n2278 ;
    wire n2279 ;
    wire n2280 ;
    wire n2281 ;
    wire n2282 ;
    wire n2283 ;
    wire n2284 ;
    wire n2285 ;
    wire n2286 ;
    wire n2287 ;
    wire n2288 ;
    wire n2289 ;
    wire n2290 ;
    wire n2291 ;
    wire n2292 ;
    wire n2293 ;
    wire n2294 ;
    wire n2295 ;
    wire n2296 ;
    wire n2297 ;
    wire n2298 ;
    wire n2299 ;
    wire n2300 ;
    wire n2301 ;
    wire n2302 ;
    wire n2303 ;
    wire n2304 ;
    wire n2305 ;
    wire n2306 ;
    wire n2307 ;
    wire n2308 ;
    wire n2309 ;
    wire n2310 ;
    wire n2311 ;
    wire n2312 ;
    wire n2313 ;
    wire n2314 ;
    wire n2315 ;
    wire n2316 ;
    wire n2317 ;
    wire n2318 ;
    wire n2319 ;
    wire n2320 ;
    wire n2321 ;
    wire n2322 ;
    wire n2323 ;
    wire n2324 ;
    wire n2325 ;
    wire n2326 ;
    wire n2327 ;
    wire n2328 ;
    wire n2329 ;
    wire n2330 ;
    wire n2331 ;
    wire n2332 ;
    wire n2333 ;
    wire n2334 ;
    wire n2335 ;
    wire n2336 ;
    wire n2337 ;
    wire n2338 ;
    wire n2339 ;
    wire n2340 ;
    wire n2341 ;
    wire n2342 ;
    wire n2343 ;
    wire n2344 ;
    wire n2345 ;
    wire n2346 ;
    wire n2347 ;
    wire n2348 ;
    wire n2349 ;
    wire n2350 ;
    wire n2351 ;
    wire n2352 ;
    wire n2353 ;
    wire n2354 ;
    wire n2355 ;
    wire n2356 ;
    wire n2357 ;
    wire n2358 ;
    wire n2359 ;
    wire n2360 ;
    wire n2361 ;
    wire n2362 ;
    wire n2363 ;
    wire n2364 ;
    wire n2365 ;
    wire n2366 ;
    wire n2367 ;
    wire n2368 ;
    wire n2369 ;
    wire n2370 ;
    wire n2371 ;
    wire n2372 ;
    wire n2373 ;
    wire n2374 ;
    wire n2375 ;
    wire n2376 ;
    wire n2377 ;
    wire n2378 ;
    wire n2379 ;
    wire n2380 ;
    wire n2381 ;
    wire n2382 ;
    wire n2383 ;
    wire n2384 ;
    wire n2385 ;
    wire n2386 ;
    wire n2387 ;
    wire n2388 ;
    wire n2389 ;
    wire n2390 ;
    wire n2391 ;
    wire n2392 ;
    wire n2393 ;
    wire n2394 ;
    wire n2395 ;
    wire n2396 ;
    wire n2397 ;
    wire n2398 ;
    wire n2399 ;
    wire n2400 ;
    wire n2401 ;
    wire n2402 ;
    wire n2403 ;
    wire n2404 ;
    wire n2405 ;
    wire n2406 ;
    wire n2407 ;
    wire n2408 ;
    wire n2409 ;
    wire n2410 ;
    wire n2411 ;
    wire n2412 ;
    wire n2413 ;
    wire n2414 ;
    wire n2415 ;
    wire n2416 ;
    wire n2417 ;
    wire n2418 ;
    wire n2419 ;
    wire n2420 ;
    wire n2421 ;
    wire n2422 ;
    wire n2423 ;
    wire n2424 ;
    wire n2425 ;
    wire n2426 ;
    wire n2427 ;
    wire n2428 ;
    wire n2429 ;
    wire n2430 ;
    wire n2431 ;
    wire n2432 ;
    wire n2433 ;
    wire n2434 ;
    wire n2435 ;
    wire n2436 ;
    wire n2437 ;
    wire n2438 ;
    wire n2439 ;
    wire n2440 ;
    wire n2441 ;
    wire n2442 ;
    wire n2443 ;
    wire n2444 ;
    wire n2445 ;
    wire n2446 ;
    wire n2447 ;
    wire n2448 ;
    wire n2449 ;
    wire n2450 ;
    wire n2451 ;
    wire n2452 ;
    wire n2453 ;
    wire n2454 ;
    wire n2455 ;
    wire n2456 ;
    wire n2457 ;
    wire n2458 ;
    wire n2459 ;
    wire n2460 ;
    wire n2461 ;
    wire n2462 ;
    wire n2463 ;
    wire n2464 ;
    wire n2465 ;
    wire n2466 ;
    wire n2467 ;
    wire n2468 ;
    wire n2469 ;
    wire n2470 ;
    wire n2471 ;
    wire n2472 ;
    wire n2473 ;
    wire n2474 ;
    wire n2475 ;
    wire n2476 ;
    wire n2477 ;
    wire n2478 ;
    wire n2479 ;
    wire n2480 ;
    wire n2481 ;
    wire n2482 ;
    wire n2483 ;
    wire n2484 ;
    wire n2485 ;
    wire n2486 ;
    wire n2487 ;
    wire n2488 ;
    wire n2489 ;
    wire n2490 ;
    wire n2491 ;
    wire n2492 ;
    wire n2493 ;
    wire n2494 ;
    wire n2495 ;
    wire n2496 ;
    wire n2497 ;
    wire n2498 ;
    wire n2499 ;
    wire n2500 ;
    wire n2501 ;
    wire n2502 ;
    wire n2503 ;
    wire n2504 ;
    wire n2505 ;
    wire n2506 ;
    wire n2507 ;
    wire n2508 ;
    wire n2509 ;
    wire n2510 ;
    wire n2511 ;
    wire n2512 ;
    wire n2513 ;
    wire n2514 ;
    wire n2515 ;
    wire n2516 ;
    wire n2517 ;
    wire n2518 ;
    wire n2519 ;
    wire n2520 ;
    wire n2521 ;
    wire n2522 ;
    wire n2523 ;
    wire n2524 ;
    wire n2525 ;
    wire n2526 ;
    wire n2527 ;
    wire n2528 ;
    wire n2529 ;
    wire n2530 ;
    wire n2531 ;
    wire n2532 ;
    wire n2533 ;
    wire n2534 ;
    wire n2535 ;
    wire n2536 ;
    wire n2537 ;
    wire n2538 ;
    wire n2539 ;
    wire n2540 ;
    wire n2541 ;
    wire n2542 ;
    wire n2543 ;
    wire n2544 ;
    wire n2545 ;
    wire n2546 ;
    wire n2547 ;
    wire n2548 ;
    wire n2549 ;
    wire n2550 ;
    wire n2551 ;
    wire n2552 ;
    wire n2553 ;
    wire n2554 ;
    wire n2555 ;
    wire n2556 ;
    wire n2557 ;
    wire n2558 ;
    wire n2559 ;
    wire n2560 ;
    wire n2561 ;
    wire n2562 ;
    wire n2563 ;
    wire n2564 ;
    wire n2565 ;
    wire n2566 ;
    wire n2567 ;
    wire n2568 ;
    wire n2569 ;
    wire n2570 ;
    wire n2571 ;
    wire n2572 ;
    wire n2573 ;
    wire n2574 ;
    wire n2575 ;
    wire n2576 ;
    wire n2577 ;
    wire n2578 ;
    wire n2579 ;
    wire n2580 ;
    wire n2581 ;
    wire n2582 ;
    wire n2583 ;
    wire n2584 ;
    wire n2585 ;
    wire n2586 ;
    wire n2587 ;
    wire n2588 ;
    wire n2589 ;
    wire n2590 ;
    wire n2591 ;
    wire n2592 ;
    wire n2593 ;
    wire n2594 ;
    wire n2595 ;
    wire n2596 ;
    wire n2597 ;
    wire n2598 ;
    wire n2599 ;
    wire n2600 ;
    wire n2601 ;
    wire n2602 ;
    wire n2603 ;
    wire n2604 ;
    wire n2605 ;
    wire n2606 ;
    wire n2607 ;
    wire n2608 ;
    wire n2609 ;
    wire n2610 ;
    wire n2611 ;
    wire n2612 ;
    wire n2613 ;
    wire n2614 ;
    wire n2615 ;
    wire n2616 ;
    wire n2617 ;
    wire n2618 ;
    wire n2619 ;
    wire n2620 ;
    wire n2621 ;
    wire n2622 ;
    wire n2623 ;
    wire n2624 ;
    wire n2625 ;
    wire n2626 ;
    wire n2627 ;
    wire n2628 ;
    wire n2629 ;
    wire n2630 ;
    wire n2631 ;
    wire n2632 ;
    wire n2633 ;
    wire n2634 ;
    wire n2635 ;
    wire n2636 ;
    wire n2637 ;
    wire n2638 ;
    wire n2639 ;
    wire n2640 ;
    wire n2641 ;
    wire n2642 ;
    wire n2643 ;
    wire n2644 ;
    wire n2645 ;
    wire n2646 ;
    wire n2647 ;
    wire n2648 ;
    wire n2649 ;
    wire n2650 ;
    wire n2651 ;
    wire n2652 ;
    wire n2653 ;
    wire n2654 ;
    wire n2655 ;
    wire n2656 ;
    wire n2657 ;
    wire n2658 ;
    wire n2659 ;
    wire n2660 ;
    wire n2661 ;
    wire n2662 ;
    wire n2663 ;
    wire n2664 ;
    wire n2665 ;
    wire n2666 ;
    wire n2667 ;
    wire n2668 ;
    wire n2669 ;
    wire n2670 ;
    wire n2671 ;
    wire n2672 ;
    wire n2673 ;
    wire n2674 ;
    wire n2675 ;
    wire n2676 ;
    wire n2677 ;
    wire n2678 ;
    wire n2679 ;
    wire n2680 ;
    wire n2681 ;
    wire n2682 ;
    wire n2683 ;
    wire n2684 ;
    wire n2685 ;
    wire n2686 ;
    wire n2687 ;
    wire n2688 ;
    wire n2689 ;
    wire n2690 ;
    wire n2691 ;
    wire n2692 ;
    wire n2693 ;
    wire n2694 ;
    wire n2695 ;
    wire n2696 ;
    wire n2697 ;
    wire n2698 ;
    wire n2699 ;
    wire n2700 ;
    wire n2701 ;
    wire n2702 ;
    wire n2703 ;
    wire n2704 ;
    wire n2705 ;
    wire n2706 ;
    wire n2707 ;
    wire n2708 ;
    wire n2709 ;
    wire n2710 ;
    wire n2711 ;
    wire n2712 ;
    wire n2713 ;
    wire n2714 ;
    wire n2715 ;
    wire n2716 ;
    wire n2717 ;
    wire n2718 ;
    wire n2719 ;
    wire n2720 ;
    wire n2721 ;
    wire n2722 ;
    wire n2723 ;
    wire n2724 ;
    wire n2725 ;
    wire n2726 ;
    wire n2727 ;
    wire n2728 ;
    wire n2729 ;
    wire n2730 ;
    wire n2731 ;
    wire n2732 ;
    wire n2733 ;
    wire n2734 ;
    wire n2735 ;
    wire n2736 ;
    wire n2737 ;
    wire n2738 ;
    wire n2739 ;
    wire n2740 ;
    wire n2741 ;
    wire n2742 ;
    wire n2743 ;
    wire n2744 ;
    wire n2745 ;
    wire n2746 ;
    wire n2747 ;
    wire n2748 ;
    wire n2749 ;
    wire n2750 ;
    wire n2751 ;
    wire n2752 ;
    wire n2753 ;
    wire n2754 ;
    wire n2755 ;
    wire n2756 ;
    wire n2757 ;
    wire n2758 ;
    wire n2759 ;
    wire n2760 ;
    wire n2761 ;
    wire n2762 ;
    wire n2763 ;
    wire n2764 ;
    wire n2765 ;
    wire n2766 ;
    wire n2767 ;
    wire n2768 ;
    wire n2769 ;
    wire n2770 ;
    wire n2771 ;
    wire n2772 ;
    wire n2773 ;
    wire n2774 ;
    wire n2775 ;
    wire n2776 ;
    wire n2777 ;
    wire n2778 ;
    wire n2779 ;
    wire n2780 ;
    wire n2781 ;
    wire n2782 ;
    wire n2783 ;
    wire n2784 ;
    wire n2785 ;
    wire n2786 ;
    wire n2787 ;
    wire n2788 ;
    wire n2789 ;
    wire n2790 ;
    wire n2791 ;
    wire n2792 ;
    wire n2793 ;
    wire n2794 ;
    wire n2795 ;
    wire n2796 ;
    wire n2797 ;
    wire n2798 ;
    wire n2799 ;
    wire n2800 ;
    wire n2801 ;
    wire n2802 ;
    wire n2803 ;
    wire n2804 ;
    wire n2805 ;
    wire n2806 ;
    wire n2807 ;
    wire n2808 ;
    wire n2809 ;
    wire n2810 ;
    wire n2811 ;
    wire n2812 ;
    wire n2813 ;
    wire n2814 ;
    wire n2815 ;
    wire n2816 ;
    wire n2817 ;
    wire n2818 ;
    wire n2819 ;
    wire n2820 ;
    wire n2821 ;
    wire n2822 ;
    wire n2823 ;
    wire n2824 ;
    wire n2825 ;
    wire n2826 ;
    wire n2827 ;
    wire n2828 ;
    wire n2829 ;
    wire n2830 ;
    wire n2831 ;
    wire n2832 ;
    wire new_AGEMA_signal_944 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_948 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_952 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_956 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_960 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_968 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_974 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_980 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_984 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_986 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_992 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7663 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7665 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7669 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7671 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7675 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7677 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7873 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7875 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7879 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7881 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7885 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7887 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7891 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7893 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7897 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7899 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7903 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7905 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8097 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8099 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8101 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8103 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8105 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8107 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8109 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8111 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8113 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8115 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8117 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8119 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8121 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8123 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8125 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8127 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8129 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8131 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8133 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8135 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8137 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8139 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8141 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8143 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8145 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8147 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8149 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8151 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8153 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8155 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8157 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8159 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8194 ;
    wire new_AGEMA_signal_8195 ;
    wire new_AGEMA_signal_8196 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8200 ;
    wire new_AGEMA_signal_8201 ;
    wire new_AGEMA_signal_8202 ;
    wire new_AGEMA_signal_8203 ;
    wire new_AGEMA_signal_8204 ;
    wire new_AGEMA_signal_8205 ;
    wire new_AGEMA_signal_8206 ;
    wire new_AGEMA_signal_8207 ;
    wire new_AGEMA_signal_8208 ;
    wire new_AGEMA_signal_8209 ;
    wire new_AGEMA_signal_8210 ;
    wire new_AGEMA_signal_8211 ;
    wire new_AGEMA_signal_8212 ;
    wire new_AGEMA_signal_8213 ;
    wire new_AGEMA_signal_8214 ;
    wire new_AGEMA_signal_8215 ;
    wire new_AGEMA_signal_8216 ;
    wire new_AGEMA_signal_8217 ;
    wire new_AGEMA_signal_8218 ;
    wire new_AGEMA_signal_8219 ;
    wire new_AGEMA_signal_8220 ;
    wire new_AGEMA_signal_8221 ;
    wire new_AGEMA_signal_8222 ;
    wire new_AGEMA_signal_8223 ;
    wire new_AGEMA_signal_8224 ;
    wire new_AGEMA_signal_8225 ;
    wire new_AGEMA_signal_8226 ;
    wire new_AGEMA_signal_8227 ;
    wire new_AGEMA_signal_8228 ;
    wire new_AGEMA_signal_8229 ;
    wire new_AGEMA_signal_8230 ;
    wire new_AGEMA_signal_8231 ;
    wire new_AGEMA_signal_8232 ;
    wire new_AGEMA_signal_8233 ;
    wire new_AGEMA_signal_8234 ;
    wire new_AGEMA_signal_8235 ;
    wire new_AGEMA_signal_8236 ;
    wire new_AGEMA_signal_8237 ;
    wire new_AGEMA_signal_8238 ;
    wire new_AGEMA_signal_8239 ;
    wire new_AGEMA_signal_8240 ;
    wire new_AGEMA_signal_8241 ;
    wire new_AGEMA_signal_8242 ;
    wire new_AGEMA_signal_8243 ;
    wire new_AGEMA_signal_8244 ;
    wire new_AGEMA_signal_8245 ;
    wire new_AGEMA_signal_8246 ;
    wire new_AGEMA_signal_8247 ;
    wire new_AGEMA_signal_8248 ;
    wire new_AGEMA_signal_8249 ;
    wire new_AGEMA_signal_8250 ;
    wire new_AGEMA_signal_8251 ;
    wire new_AGEMA_signal_8252 ;
    wire new_AGEMA_signal_8253 ;
    wire new_AGEMA_signal_8254 ;
    wire new_AGEMA_signal_8255 ;
    wire new_AGEMA_signal_8256 ;
    wire new_AGEMA_signal_8257 ;
    wire new_AGEMA_signal_8258 ;
    wire new_AGEMA_signal_8259 ;
    wire new_AGEMA_signal_8260 ;
    wire new_AGEMA_signal_8261 ;
    wire new_AGEMA_signal_8262 ;
    wire new_AGEMA_signal_8263 ;
    wire new_AGEMA_signal_8264 ;
    wire new_AGEMA_signal_8265 ;
    wire new_AGEMA_signal_8266 ;
    wire new_AGEMA_signal_8267 ;
    wire new_AGEMA_signal_8268 ;
    wire new_AGEMA_signal_8269 ;
    wire new_AGEMA_signal_8270 ;
    wire new_AGEMA_signal_8271 ;
    wire new_AGEMA_signal_8272 ;
    wire new_AGEMA_signal_8273 ;
    wire new_AGEMA_signal_8274 ;
    wire new_AGEMA_signal_8275 ;
    wire new_AGEMA_signal_8276 ;
    wire new_AGEMA_signal_8277 ;
    wire new_AGEMA_signal_8278 ;
    wire new_AGEMA_signal_8279 ;
    wire new_AGEMA_signal_8280 ;
    wire new_AGEMA_signal_8281 ;
    wire new_AGEMA_signal_8282 ;
    wire new_AGEMA_signal_8283 ;
    wire new_AGEMA_signal_8284 ;
    wire new_AGEMA_signal_8285 ;
    wire new_AGEMA_signal_8286 ;
    wire new_AGEMA_signal_8287 ;
    wire new_AGEMA_signal_8288 ;
    wire new_AGEMA_signal_8289 ;
    wire new_AGEMA_signal_8290 ;
    wire new_AGEMA_signal_8291 ;
    wire new_AGEMA_signal_8292 ;
    wire new_AGEMA_signal_8293 ;
    wire new_AGEMA_signal_8294 ;
    wire new_AGEMA_signal_8295 ;
    wire new_AGEMA_signal_8296 ;
    wire new_AGEMA_signal_8297 ;
    wire new_AGEMA_signal_8298 ;
    wire new_AGEMA_signal_8299 ;
    wire new_AGEMA_signal_8300 ;
    wire new_AGEMA_signal_8301 ;
    wire new_AGEMA_signal_8302 ;
    wire new_AGEMA_signal_8303 ;
    wire new_AGEMA_signal_8304 ;
    wire new_AGEMA_signal_8305 ;
    wire new_AGEMA_signal_8306 ;
    wire new_AGEMA_signal_8307 ;
    wire new_AGEMA_signal_8308 ;
    wire new_AGEMA_signal_8309 ;
    wire new_AGEMA_signal_8310 ;
    wire new_AGEMA_signal_8311 ;
    wire new_AGEMA_signal_8312 ;
    wire new_AGEMA_signal_8313 ;
    wire new_AGEMA_signal_8314 ;
    wire new_AGEMA_signal_8315 ;
    wire new_AGEMA_signal_8316 ;
    wire new_AGEMA_signal_8317 ;
    wire new_AGEMA_signal_8318 ;
    wire new_AGEMA_signal_8319 ;
    wire new_AGEMA_signal_8320 ;
    wire new_AGEMA_signal_8321 ;
    wire new_AGEMA_signal_8322 ;
    wire new_AGEMA_signal_8323 ;
    wire new_AGEMA_signal_8324 ;
    wire new_AGEMA_signal_8325 ;
    wire new_AGEMA_signal_8326 ;
    wire new_AGEMA_signal_8327 ;
    wire new_AGEMA_signal_8328 ;
    wire new_AGEMA_signal_8329 ;
    wire new_AGEMA_signal_8330 ;
    wire new_AGEMA_signal_8331 ;
    wire new_AGEMA_signal_8332 ;
    wire new_AGEMA_signal_8333 ;
    wire new_AGEMA_signal_8334 ;
    wire new_AGEMA_signal_8335 ;
    wire new_AGEMA_signal_8336 ;
    wire new_AGEMA_signal_8337 ;
    wire new_AGEMA_signal_8338 ;
    wire new_AGEMA_signal_8339 ;
    wire new_AGEMA_signal_8340 ;
    wire new_AGEMA_signal_8341 ;
    wire new_AGEMA_signal_8342 ;
    wire new_AGEMA_signal_8343 ;
    wire new_AGEMA_signal_8344 ;
    wire new_AGEMA_signal_8345 ;
    wire new_AGEMA_signal_8346 ;
    wire new_AGEMA_signal_8347 ;
    wire new_AGEMA_signal_8348 ;
    wire new_AGEMA_signal_8349 ;
    wire new_AGEMA_signal_8350 ;
    wire new_AGEMA_signal_8351 ;
    wire new_AGEMA_signal_8352 ;
    wire new_AGEMA_signal_8353 ;
    wire new_AGEMA_signal_8354 ;
    wire new_AGEMA_signal_8355 ;
    wire new_AGEMA_signal_8356 ;
    wire new_AGEMA_signal_8357 ;
    wire new_AGEMA_signal_8358 ;
    wire new_AGEMA_signal_8359 ;
    wire new_AGEMA_signal_8360 ;
    wire new_AGEMA_signal_8361 ;
    wire new_AGEMA_signal_8362 ;
    wire new_AGEMA_signal_8363 ;
    wire new_AGEMA_signal_8364 ;
    wire new_AGEMA_signal_8365 ;
    wire new_AGEMA_signal_8366 ;
    wire new_AGEMA_signal_8367 ;
    wire new_AGEMA_signal_8368 ;
    wire new_AGEMA_signal_8369 ;
    wire new_AGEMA_signal_8370 ;
    wire new_AGEMA_signal_8371 ;
    wire new_AGEMA_signal_8372 ;
    wire new_AGEMA_signal_8373 ;
    wire new_AGEMA_signal_8374 ;
    wire new_AGEMA_signal_8375 ;
    wire new_AGEMA_signal_8376 ;
    wire new_AGEMA_signal_8377 ;
    wire new_AGEMA_signal_8378 ;
    wire new_AGEMA_signal_8379 ;
    wire new_AGEMA_signal_8380 ;
    wire new_AGEMA_signal_8381 ;
    wire new_AGEMA_signal_8382 ;
    wire new_AGEMA_signal_8383 ;
    wire new_AGEMA_signal_8384 ;
    wire new_AGEMA_signal_8385 ;
    wire new_AGEMA_signal_8386 ;
    wire new_AGEMA_signal_8387 ;
    wire new_AGEMA_signal_8388 ;
    wire new_AGEMA_signal_8389 ;
    wire new_AGEMA_signal_8390 ;
    wire new_AGEMA_signal_8391 ;
    wire new_AGEMA_signal_8392 ;
    wire new_AGEMA_signal_8393 ;
    wire new_AGEMA_signal_8394 ;
    wire new_AGEMA_signal_8395 ;
    wire new_AGEMA_signal_8396 ;
    wire new_AGEMA_signal_8397 ;
    wire new_AGEMA_signal_8398 ;
    wire new_AGEMA_signal_8399 ;
    wire new_AGEMA_signal_8400 ;
    wire new_AGEMA_signal_8401 ;
    wire new_AGEMA_signal_8402 ;
    wire new_AGEMA_signal_8403 ;
    wire new_AGEMA_signal_8404 ;
    wire new_AGEMA_signal_8405 ;
    wire new_AGEMA_signal_8406 ;
    wire new_AGEMA_signal_8407 ;
    wire new_AGEMA_signal_8408 ;
    wire new_AGEMA_signal_8409 ;
    wire new_AGEMA_signal_8410 ;
    wire new_AGEMA_signal_8411 ;
    wire new_AGEMA_signal_8412 ;
    wire new_AGEMA_signal_8413 ;
    wire new_AGEMA_signal_8414 ;
    wire new_AGEMA_signal_8415 ;
    wire new_AGEMA_signal_8416 ;
    wire new_AGEMA_signal_8417 ;
    wire new_AGEMA_signal_8418 ;
    wire new_AGEMA_signal_8419 ;
    wire new_AGEMA_signal_8420 ;
    wire new_AGEMA_signal_8421 ;
    wire new_AGEMA_signal_8422 ;
    wire new_AGEMA_signal_8423 ;
    wire new_AGEMA_signal_8424 ;
    wire new_AGEMA_signal_8425 ;
    wire new_AGEMA_signal_8426 ;
    wire new_AGEMA_signal_8427 ;
    wire new_AGEMA_signal_8428 ;
    wire new_AGEMA_signal_8429 ;
    wire new_AGEMA_signal_8430 ;
    wire new_AGEMA_signal_8431 ;
    wire new_AGEMA_signal_8432 ;
    wire new_AGEMA_signal_8433 ;
    wire new_AGEMA_signal_8434 ;
    wire new_AGEMA_signal_8435 ;
    wire new_AGEMA_signal_8436 ;
    wire new_AGEMA_signal_8437 ;
    wire new_AGEMA_signal_8438 ;
    wire new_AGEMA_signal_8439 ;
    wire new_AGEMA_signal_8440 ;
    wire new_AGEMA_signal_8441 ;
    wire new_AGEMA_signal_8442 ;
    wire new_AGEMA_signal_8443 ;
    wire new_AGEMA_signal_8444 ;
    wire new_AGEMA_signal_8445 ;
    wire new_AGEMA_signal_8446 ;
    wire new_AGEMA_signal_8447 ;
    wire new_AGEMA_signal_8448 ;
    wire new_AGEMA_signal_8449 ;
    wire new_AGEMA_signal_8450 ;
    wire new_AGEMA_signal_8451 ;
    wire new_AGEMA_signal_8452 ;
    wire new_AGEMA_signal_8453 ;
    wire new_AGEMA_signal_8454 ;
    wire new_AGEMA_signal_8455 ;
    wire new_AGEMA_signal_8456 ;
    wire new_AGEMA_signal_8457 ;
    wire new_AGEMA_signal_8458 ;
    wire new_AGEMA_signal_8459 ;
    wire new_AGEMA_signal_8460 ;
    wire new_AGEMA_signal_8461 ;
    wire new_AGEMA_signal_8462 ;
    wire new_AGEMA_signal_8463 ;
    wire new_AGEMA_signal_8464 ;
    wire new_AGEMA_signal_8465 ;
    wire new_AGEMA_signal_8466 ;
    wire new_AGEMA_signal_8467 ;
    wire new_AGEMA_signal_8468 ;
    wire new_AGEMA_signal_8469 ;
    wire new_AGEMA_signal_8470 ;
    wire new_AGEMA_signal_8471 ;
    wire new_AGEMA_signal_8472 ;
    wire new_AGEMA_signal_8473 ;
    wire new_AGEMA_signal_8474 ;
    wire new_AGEMA_signal_8475 ;
    wire new_AGEMA_signal_8476 ;
    wire new_AGEMA_signal_8477 ;
    wire new_AGEMA_signal_8478 ;
    wire new_AGEMA_signal_8479 ;
    wire new_AGEMA_signal_8480 ;
    wire new_AGEMA_signal_8481 ;
    wire new_AGEMA_signal_8482 ;
    wire new_AGEMA_signal_8483 ;
    wire new_AGEMA_signal_8484 ;
    wire new_AGEMA_signal_8485 ;
    wire new_AGEMA_signal_8486 ;
    wire new_AGEMA_signal_8487 ;
    wire new_AGEMA_signal_8488 ;
    wire new_AGEMA_signal_8489 ;
    wire new_AGEMA_signal_8490 ;
    wire new_AGEMA_signal_8491 ;
    wire new_AGEMA_signal_8492 ;
    wire new_AGEMA_signal_8493 ;
    wire new_AGEMA_signal_8494 ;
    wire new_AGEMA_signal_8495 ;
    wire new_AGEMA_signal_8496 ;
    wire new_AGEMA_signal_8497 ;
    wire new_AGEMA_signal_8498 ;
    wire new_AGEMA_signal_8499 ;
    wire new_AGEMA_signal_8500 ;
    wire new_AGEMA_signal_8501 ;
    wire new_AGEMA_signal_8502 ;
    wire new_AGEMA_signal_8503 ;
    wire new_AGEMA_signal_8504 ;
    wire new_AGEMA_signal_8505 ;
    wire new_AGEMA_signal_8506 ;
    wire new_AGEMA_signal_8507 ;
    wire new_AGEMA_signal_8508 ;
    wire new_AGEMA_signal_8509 ;
    wire new_AGEMA_signal_8510 ;
    wire new_AGEMA_signal_8511 ;
    wire new_AGEMA_signal_8512 ;
    wire new_AGEMA_signal_8513 ;
    wire new_AGEMA_signal_8514 ;
    wire new_AGEMA_signal_8515 ;
    wire new_AGEMA_signal_8516 ;
    wire new_AGEMA_signal_8517 ;
    wire new_AGEMA_signal_8518 ;
    wire new_AGEMA_signal_8519 ;
    wire new_AGEMA_signal_8520 ;
    wire new_AGEMA_signal_8521 ;
    wire new_AGEMA_signal_8522 ;
    wire new_AGEMA_signal_8523 ;
    wire new_AGEMA_signal_8524 ;
    wire new_AGEMA_signal_8525 ;
    wire new_AGEMA_signal_8526 ;
    wire new_AGEMA_signal_8527 ;
    wire new_AGEMA_signal_8528 ;
    wire new_AGEMA_signal_8529 ;
    wire new_AGEMA_signal_8530 ;
    wire new_AGEMA_signal_8531 ;
    wire new_AGEMA_signal_8532 ;
    wire new_AGEMA_signal_8533 ;
    wire new_AGEMA_signal_8534 ;
    wire new_AGEMA_signal_8535 ;
    wire new_AGEMA_signal_8536 ;
    wire new_AGEMA_signal_8537 ;
    wire new_AGEMA_signal_8538 ;
    wire new_AGEMA_signal_8539 ;
    wire new_AGEMA_signal_8540 ;
    wire new_AGEMA_signal_8541 ;
    wire new_AGEMA_signal_8542 ;
    wire new_AGEMA_signal_8543 ;
    wire new_AGEMA_signal_8544 ;
    wire new_AGEMA_signal_8545 ;
    wire new_AGEMA_signal_8546 ;
    wire new_AGEMA_signal_8547 ;
    wire new_AGEMA_signal_8548 ;
    wire new_AGEMA_signal_8549 ;
    wire new_AGEMA_signal_8550 ;
    wire new_AGEMA_signal_8551 ;
    wire new_AGEMA_signal_8552 ;
    wire new_AGEMA_signal_8553 ;
    wire new_AGEMA_signal_8554 ;
    wire new_AGEMA_signal_8555 ;
    wire new_AGEMA_signal_8556 ;
    wire new_AGEMA_signal_8557 ;
    wire new_AGEMA_signal_8558 ;
    wire new_AGEMA_signal_8559 ;
    wire new_AGEMA_signal_8560 ;
    wire new_AGEMA_signal_8561 ;
    wire new_AGEMA_signal_8562 ;
    wire new_AGEMA_signal_8563 ;
    wire new_AGEMA_signal_8564 ;
    wire new_AGEMA_signal_8565 ;
    wire new_AGEMA_signal_8566 ;
    wire new_AGEMA_signal_8567 ;
    wire new_AGEMA_signal_8568 ;
    wire new_AGEMA_signal_8569 ;
    wire new_AGEMA_signal_8570 ;
    wire new_AGEMA_signal_8571 ;
    wire new_AGEMA_signal_8572 ;
    wire new_AGEMA_signal_8573 ;
    wire new_AGEMA_signal_8574 ;
    wire new_AGEMA_signal_8575 ;
    wire new_AGEMA_signal_8576 ;
    wire new_AGEMA_signal_8577 ;
    wire new_AGEMA_signal_8578 ;
    wire new_AGEMA_signal_8579 ;
    wire new_AGEMA_signal_8580 ;
    wire new_AGEMA_signal_8581 ;
    wire new_AGEMA_signal_8582 ;
    wire new_AGEMA_signal_8583 ;
    wire new_AGEMA_signal_8584 ;
    wire new_AGEMA_signal_8585 ;
    wire new_AGEMA_signal_8586 ;
    wire new_AGEMA_signal_8587 ;
    wire new_AGEMA_signal_8588 ;
    wire new_AGEMA_signal_8589 ;
    wire new_AGEMA_signal_8590 ;
    wire new_AGEMA_signal_8591 ;
    wire new_AGEMA_signal_8592 ;
    wire new_AGEMA_signal_8593 ;
    wire new_AGEMA_signal_8594 ;
    wire new_AGEMA_signal_8595 ;
    wire new_AGEMA_signal_8596 ;
    wire new_AGEMA_signal_8597 ;
    wire new_AGEMA_signal_8598 ;
    wire new_AGEMA_signal_8599 ;
    wire new_AGEMA_signal_8600 ;
    wire new_AGEMA_signal_8601 ;
    wire new_AGEMA_signal_8602 ;
    wire new_AGEMA_signal_8603 ;
    wire new_AGEMA_signal_8604 ;
    wire new_AGEMA_signal_8605 ;
    wire new_AGEMA_signal_8606 ;
    wire new_AGEMA_signal_8607 ;
    wire new_AGEMA_signal_8608 ;
    wire new_AGEMA_signal_8609 ;
    wire new_AGEMA_signal_8610 ;
    wire new_AGEMA_signal_8611 ;
    wire new_AGEMA_signal_8612 ;
    wire new_AGEMA_signal_8613 ;
    wire new_AGEMA_signal_8614 ;
    wire new_AGEMA_signal_8615 ;
    wire new_AGEMA_signal_8616 ;
    wire new_AGEMA_signal_8617 ;
    wire new_AGEMA_signal_8618 ;
    wire new_AGEMA_signal_8619 ;
    wire new_AGEMA_signal_8620 ;
    wire new_AGEMA_signal_8621 ;
    wire new_AGEMA_signal_8622 ;
    wire new_AGEMA_signal_8623 ;
    wire new_AGEMA_signal_8624 ;
    wire new_AGEMA_signal_8625 ;
    wire new_AGEMA_signal_8626 ;
    wire new_AGEMA_signal_8627 ;
    wire new_AGEMA_signal_8628 ;
    wire new_AGEMA_signal_8629 ;
    wire new_AGEMA_signal_8630 ;
    wire new_AGEMA_signal_8631 ;
    wire new_AGEMA_signal_8632 ;
    wire new_AGEMA_signal_8633 ;
    wire new_AGEMA_signal_8634 ;
    wire new_AGEMA_signal_8635 ;
    wire new_AGEMA_signal_8636 ;
    wire new_AGEMA_signal_8637 ;
    wire new_AGEMA_signal_8638 ;
    wire new_AGEMA_signal_8639 ;
    wire new_AGEMA_signal_8640 ;
    wire new_AGEMA_signal_8641 ;
    wire new_AGEMA_signal_8642 ;
    wire new_AGEMA_signal_8643 ;
    wire new_AGEMA_signal_8644 ;
    wire new_AGEMA_signal_8645 ;
    wire new_AGEMA_signal_8646 ;
    wire new_AGEMA_signal_8647 ;
    wire new_AGEMA_signal_8648 ;
    wire new_AGEMA_signal_8649 ;
    wire new_AGEMA_signal_8650 ;
    wire new_AGEMA_signal_8651 ;
    wire new_AGEMA_signal_8652 ;
    wire new_AGEMA_signal_8653 ;
    wire new_AGEMA_signal_8654 ;
    wire new_AGEMA_signal_8655 ;
    wire new_AGEMA_signal_8656 ;
    wire new_AGEMA_signal_8657 ;
    wire new_AGEMA_signal_8658 ;
    wire new_AGEMA_signal_8659 ;
    wire new_AGEMA_signal_8660 ;
    wire new_AGEMA_signal_8661 ;
    wire new_AGEMA_signal_8662 ;
    wire new_AGEMA_signal_8663 ;
    wire new_AGEMA_signal_8664 ;
    wire new_AGEMA_signal_8665 ;
    wire new_AGEMA_signal_8666 ;
    wire new_AGEMA_signal_8667 ;
    wire new_AGEMA_signal_8668 ;
    wire new_AGEMA_signal_8669 ;
    wire new_AGEMA_signal_8670 ;
    wire new_AGEMA_signal_8671 ;
    wire new_AGEMA_signal_8672 ;
    wire new_AGEMA_signal_8673 ;
    wire new_AGEMA_signal_8674 ;
    wire new_AGEMA_signal_8675 ;
    wire new_AGEMA_signal_8676 ;
    wire new_AGEMA_signal_8677 ;
    wire new_AGEMA_signal_8678 ;
    wire new_AGEMA_signal_8679 ;
    wire new_AGEMA_signal_8680 ;
    wire new_AGEMA_signal_8681 ;
    wire new_AGEMA_signal_8682 ;
    wire new_AGEMA_signal_8683 ;
    wire new_AGEMA_signal_8684 ;
    wire new_AGEMA_signal_8685 ;
    wire new_AGEMA_signal_8686 ;
    wire new_AGEMA_signal_8687 ;
    wire new_AGEMA_signal_8688 ;
    wire new_AGEMA_signal_8689 ;
    wire new_AGEMA_signal_8690 ;
    wire new_AGEMA_signal_8691 ;
    wire new_AGEMA_signal_8692 ;
    wire new_AGEMA_signal_8693 ;
    wire new_AGEMA_signal_8694 ;
    wire new_AGEMA_signal_8695 ;
    wire new_AGEMA_signal_8696 ;
    wire new_AGEMA_signal_8697 ;
    wire new_AGEMA_signal_8698 ;
    wire new_AGEMA_signal_8699 ;
    wire new_AGEMA_signal_8700 ;
    wire new_AGEMA_signal_8701 ;
    wire new_AGEMA_signal_8702 ;
    wire new_AGEMA_signal_8703 ;
    wire new_AGEMA_signal_8704 ;
    wire new_AGEMA_signal_8705 ;
    wire new_AGEMA_signal_8706 ;
    wire new_AGEMA_signal_8707 ;
    wire new_AGEMA_signal_8708 ;
    wire new_AGEMA_signal_8709 ;
    wire new_AGEMA_signal_8710 ;
    wire new_AGEMA_signal_8711 ;
    wire new_AGEMA_signal_8712 ;
    wire new_AGEMA_signal_8713 ;
    wire new_AGEMA_signal_8714 ;
    wire new_AGEMA_signal_8715 ;
    wire new_AGEMA_signal_8716 ;
    wire new_AGEMA_signal_8717 ;
    wire new_AGEMA_signal_8718 ;
    wire new_AGEMA_signal_8719 ;
    wire new_AGEMA_signal_8720 ;
    wire new_AGEMA_signal_8721 ;
    wire new_AGEMA_signal_8722 ;
    wire new_AGEMA_signal_8723 ;
    wire new_AGEMA_signal_8724 ;
    wire new_AGEMA_signal_8725 ;
    wire new_AGEMA_signal_8726 ;
    wire new_AGEMA_signal_8727 ;
    wire new_AGEMA_signal_8728 ;
    wire new_AGEMA_signal_8729 ;
    wire new_AGEMA_signal_8730 ;
    wire new_AGEMA_signal_8731 ;
    wire new_AGEMA_signal_8732 ;
    wire new_AGEMA_signal_8733 ;
    wire new_AGEMA_signal_8734 ;
    wire new_AGEMA_signal_8735 ;
    wire new_AGEMA_signal_8736 ;
    wire new_AGEMA_signal_8737 ;
    wire new_AGEMA_signal_8738 ;
    wire new_AGEMA_signal_8739 ;
    wire new_AGEMA_signal_8740 ;
    wire new_AGEMA_signal_8741 ;
    wire new_AGEMA_signal_8742 ;
    wire new_AGEMA_signal_8743 ;
    wire new_AGEMA_signal_8744 ;
    wire new_AGEMA_signal_8745 ;
    wire new_AGEMA_signal_8746 ;
    wire new_AGEMA_signal_8747 ;
    wire new_AGEMA_signal_8748 ;
    wire new_AGEMA_signal_8749 ;
    wire new_AGEMA_signal_8750 ;
    wire new_AGEMA_signal_8751 ;
    wire new_AGEMA_signal_8752 ;
    wire new_AGEMA_signal_8753 ;
    wire new_AGEMA_signal_8754 ;
    wire new_AGEMA_signal_8755 ;
    wire new_AGEMA_signal_8756 ;
    wire new_AGEMA_signal_8757 ;
    wire new_AGEMA_signal_8758 ;
    wire new_AGEMA_signal_8759 ;
    wire new_AGEMA_signal_8760 ;
    wire new_AGEMA_signal_8761 ;
    wire new_AGEMA_signal_8762 ;
    wire new_AGEMA_signal_8763 ;
    wire new_AGEMA_signal_8764 ;
    wire new_AGEMA_signal_8765 ;
    wire new_AGEMA_signal_8766 ;
    wire new_AGEMA_signal_8767 ;
    wire new_AGEMA_signal_8768 ;
    wire new_AGEMA_signal_8769 ;
    wire new_AGEMA_signal_8770 ;
    wire new_AGEMA_signal_8771 ;
    wire new_AGEMA_signal_8772 ;
    wire new_AGEMA_signal_8773 ;
    wire new_AGEMA_signal_8774 ;
    wire new_AGEMA_signal_8775 ;
    wire new_AGEMA_signal_8776 ;
    wire new_AGEMA_signal_8777 ;
    wire new_AGEMA_signal_8778 ;
    wire new_AGEMA_signal_8779 ;
    wire new_AGEMA_signal_8780 ;
    wire new_AGEMA_signal_8781 ;
    wire new_AGEMA_signal_8782 ;
    wire new_AGEMA_signal_8783 ;
    wire new_AGEMA_signal_8784 ;
    wire new_AGEMA_signal_8785 ;
    wire new_AGEMA_signal_8786 ;
    wire new_AGEMA_signal_8787 ;
    wire new_AGEMA_signal_8788 ;
    wire new_AGEMA_signal_8789 ;
    wire new_AGEMA_signal_8790 ;
    wire new_AGEMA_signal_8791 ;
    wire new_AGEMA_signal_8792 ;
    wire new_AGEMA_signal_8793 ;
    wire new_AGEMA_signal_8794 ;
    wire new_AGEMA_signal_8795 ;
    wire new_AGEMA_signal_8796 ;
    wire new_AGEMA_signal_8797 ;
    wire new_AGEMA_signal_8798 ;
    wire new_AGEMA_signal_8799 ;
    wire new_AGEMA_signal_8800 ;
    wire new_AGEMA_signal_8801 ;
    wire new_AGEMA_signal_8802 ;
    wire new_AGEMA_signal_8803 ;
    wire new_AGEMA_signal_8804 ;
    wire new_AGEMA_signal_8805 ;
    wire new_AGEMA_signal_8806 ;
    wire new_AGEMA_signal_8807 ;
    wire new_AGEMA_signal_8808 ;
    wire new_AGEMA_signal_8809 ;
    wire new_AGEMA_signal_8810 ;
    wire new_AGEMA_signal_8811 ;
    wire new_AGEMA_signal_8812 ;
    wire new_AGEMA_signal_8813 ;
    wire new_AGEMA_signal_8814 ;
    wire new_AGEMA_signal_8815 ;
    wire new_AGEMA_signal_8816 ;
    wire new_AGEMA_signal_8817 ;
    wire new_AGEMA_signal_8818 ;
    wire new_AGEMA_signal_8819 ;
    wire new_AGEMA_signal_8820 ;
    wire new_AGEMA_signal_8821 ;
    wire new_AGEMA_signal_8822 ;
    wire new_AGEMA_signal_8823 ;
    wire new_AGEMA_signal_8824 ;
    wire new_AGEMA_signal_8825 ;
    wire new_AGEMA_signal_8826 ;
    wire new_AGEMA_signal_8827 ;
    wire new_AGEMA_signal_8828 ;
    wire new_AGEMA_signal_8829 ;
    wire new_AGEMA_signal_8830 ;
    wire new_AGEMA_signal_8831 ;
    wire new_AGEMA_signal_8832 ;
    wire new_AGEMA_signal_8833 ;
    wire new_AGEMA_signal_8834 ;
    wire new_AGEMA_signal_8835 ;
    wire new_AGEMA_signal_8836 ;
    wire new_AGEMA_signal_8837 ;
    wire new_AGEMA_signal_8838 ;
    wire new_AGEMA_signal_8839 ;
    wire new_AGEMA_signal_8840 ;
    wire new_AGEMA_signal_8841 ;
    wire new_AGEMA_signal_8842 ;
    wire new_AGEMA_signal_8843 ;
    wire new_AGEMA_signal_8844 ;
    wire new_AGEMA_signal_8845 ;
    wire new_AGEMA_signal_8846 ;
    wire new_AGEMA_signal_8847 ;
    wire new_AGEMA_signal_8848 ;
    wire new_AGEMA_signal_8849 ;
    wire new_AGEMA_signal_8850 ;
    wire new_AGEMA_signal_8851 ;
    wire new_AGEMA_signal_8852 ;
    wire new_AGEMA_signal_8853 ;
    wire new_AGEMA_signal_8854 ;
    wire new_AGEMA_signal_8855 ;
    wire new_AGEMA_signal_8856 ;
    wire new_AGEMA_signal_8857 ;
    wire new_AGEMA_signal_8858 ;
    wire new_AGEMA_signal_8859 ;
    wire new_AGEMA_signal_8860 ;
    wire new_AGEMA_signal_8861 ;
    wire new_AGEMA_signal_8862 ;
    wire new_AGEMA_signal_8863 ;
    wire new_AGEMA_signal_8864 ;
    wire new_AGEMA_signal_8865 ;
    wire new_AGEMA_signal_8866 ;
    wire new_AGEMA_signal_8867 ;
    wire new_AGEMA_signal_8868 ;
    wire new_AGEMA_signal_8869 ;
    wire new_AGEMA_signal_8870 ;
    wire new_AGEMA_signal_8871 ;
    wire new_AGEMA_signal_8872 ;
    wire new_AGEMA_signal_8873 ;
    wire new_AGEMA_signal_8874 ;
    wire new_AGEMA_signal_8875 ;
    wire new_AGEMA_signal_8876 ;
    wire new_AGEMA_signal_8877 ;
    wire new_AGEMA_signal_8878 ;
    wire new_AGEMA_signal_8879 ;
    wire new_AGEMA_signal_8880 ;
    wire new_AGEMA_signal_8881 ;
    wire new_AGEMA_signal_8882 ;
    wire new_AGEMA_signal_8883 ;
    wire new_AGEMA_signal_8884 ;
    wire new_AGEMA_signal_8885 ;
    wire new_AGEMA_signal_8886 ;
    wire new_AGEMA_signal_8887 ;
    wire new_AGEMA_signal_8888 ;
    wire new_AGEMA_signal_8889 ;
    wire new_AGEMA_signal_8890 ;
    wire new_AGEMA_signal_8891 ;
    wire new_AGEMA_signal_8892 ;
    wire new_AGEMA_signal_8893 ;
    wire new_AGEMA_signal_8894 ;
    wire new_AGEMA_signal_8895 ;
    wire new_AGEMA_signal_8896 ;
    wire new_AGEMA_signal_8897 ;
    wire new_AGEMA_signal_8898 ;
    wire new_AGEMA_signal_8899 ;
    wire new_AGEMA_signal_8900 ;
    wire new_AGEMA_signal_8901 ;
    wire new_AGEMA_signal_8902 ;
    wire new_AGEMA_signal_8903 ;
    wire new_AGEMA_signal_8904 ;
    wire new_AGEMA_signal_8905 ;
    wire new_AGEMA_signal_8906 ;
    wire new_AGEMA_signal_8907 ;
    wire new_AGEMA_signal_8908 ;
    wire new_AGEMA_signal_8909 ;
    wire new_AGEMA_signal_8910 ;
    wire new_AGEMA_signal_8911 ;
    wire new_AGEMA_signal_8912 ;
    wire new_AGEMA_signal_8913 ;
    wire new_AGEMA_signal_8914 ;
    wire new_AGEMA_signal_8915 ;
    wire new_AGEMA_signal_8916 ;
    wire new_AGEMA_signal_8917 ;
    wire new_AGEMA_signal_8918 ;
    wire new_AGEMA_signal_8919 ;
    wire new_AGEMA_signal_8920 ;
    wire new_AGEMA_signal_8921 ;
    wire new_AGEMA_signal_8922 ;
    wire new_AGEMA_signal_8923 ;
    wire new_AGEMA_signal_8924 ;
    wire new_AGEMA_signal_8925 ;
    wire new_AGEMA_signal_8926 ;
    wire new_AGEMA_signal_8927 ;
    wire new_AGEMA_signal_8928 ;
    wire new_AGEMA_signal_8929 ;
    wire new_AGEMA_signal_8930 ;
    wire new_AGEMA_signal_8931 ;
    wire new_AGEMA_signal_8932 ;
    wire new_AGEMA_signal_8933 ;
    wire new_AGEMA_signal_8934 ;
    wire new_AGEMA_signal_8935 ;
    wire new_AGEMA_signal_8936 ;
    wire new_AGEMA_signal_8937 ;
    wire new_AGEMA_signal_8938 ;
    wire new_AGEMA_signal_8939 ;
    wire new_AGEMA_signal_8940 ;
    wire new_AGEMA_signal_8941 ;
    wire new_AGEMA_signal_8942 ;
    wire new_AGEMA_signal_8943 ;
    wire new_AGEMA_signal_8944 ;
    wire new_AGEMA_signal_8945 ;
    wire new_AGEMA_signal_8946 ;
    wire new_AGEMA_signal_8947 ;
    wire new_AGEMA_signal_8948 ;
    wire new_AGEMA_signal_8949 ;
    wire new_AGEMA_signal_8950 ;
    wire new_AGEMA_signal_8951 ;
    wire new_AGEMA_signal_8952 ;
    wire new_AGEMA_signal_8953 ;
    wire new_AGEMA_signal_8954 ;
    wire new_AGEMA_signal_8955 ;
    wire new_AGEMA_signal_8956 ;
    wire new_AGEMA_signal_8957 ;
    wire new_AGEMA_signal_8958 ;
    wire new_AGEMA_signal_8959 ;
    wire new_AGEMA_signal_8960 ;
    wire new_AGEMA_signal_8961 ;
    wire new_AGEMA_signal_8962 ;
    wire new_AGEMA_signal_8963 ;
    wire new_AGEMA_signal_8964 ;
    wire new_AGEMA_signal_8965 ;
    wire new_AGEMA_signal_8966 ;
    wire new_AGEMA_signal_8967 ;
    wire new_AGEMA_signal_8968 ;
    wire new_AGEMA_signal_8969 ;
    wire new_AGEMA_signal_8970 ;
    wire new_AGEMA_signal_8971 ;
    wire new_AGEMA_signal_8972 ;
    wire new_AGEMA_signal_8973 ;
    wire new_AGEMA_signal_8974 ;
    wire new_AGEMA_signal_8975 ;
    wire new_AGEMA_signal_8976 ;
    wire new_AGEMA_signal_8977 ;
    wire new_AGEMA_signal_8978 ;
    wire new_AGEMA_signal_8979 ;
    wire new_AGEMA_signal_8980 ;
    wire new_AGEMA_signal_8981 ;
    wire new_AGEMA_signal_8982 ;
    wire new_AGEMA_signal_8983 ;
    wire new_AGEMA_signal_8984 ;
    wire new_AGEMA_signal_8985 ;
    wire new_AGEMA_signal_8986 ;
    wire new_AGEMA_signal_8987 ;
    wire new_AGEMA_signal_8988 ;
    wire new_AGEMA_signal_8989 ;
    wire new_AGEMA_signal_8990 ;
    wire new_AGEMA_signal_8991 ;
    wire new_AGEMA_signal_8992 ;
    wire new_AGEMA_signal_8993 ;
    wire new_AGEMA_signal_8994 ;
    wire new_AGEMA_signal_8995 ;
    wire new_AGEMA_signal_8996 ;
    wire new_AGEMA_signal_8997 ;
    wire new_AGEMA_signal_8998 ;
    wire new_AGEMA_signal_8999 ;
    wire new_AGEMA_signal_9000 ;
    wire new_AGEMA_signal_9001 ;
    wire new_AGEMA_signal_9002 ;
    wire new_AGEMA_signal_9003 ;
    wire new_AGEMA_signal_9004 ;
    wire new_AGEMA_signal_9005 ;
    wire new_AGEMA_signal_9006 ;
    wire new_AGEMA_signal_9007 ;
    wire new_AGEMA_signal_9008 ;
    wire new_AGEMA_signal_9009 ;
    wire new_AGEMA_signal_9010 ;
    wire new_AGEMA_signal_9011 ;
    wire new_AGEMA_signal_9012 ;
    wire new_AGEMA_signal_9013 ;
    wire new_AGEMA_signal_9014 ;
    wire new_AGEMA_signal_9015 ;
    wire new_AGEMA_signal_9016 ;
    wire new_AGEMA_signal_9017 ;
    wire new_AGEMA_signal_9018 ;
    wire new_AGEMA_signal_9019 ;
    wire new_AGEMA_signal_9020 ;
    wire new_AGEMA_signal_9021 ;
    wire new_AGEMA_signal_9022 ;
    wire new_AGEMA_signal_9023 ;
    wire new_AGEMA_signal_9024 ;
    wire new_AGEMA_signal_9025 ;
    wire new_AGEMA_signal_9026 ;
    wire new_AGEMA_signal_9027 ;
    wire new_AGEMA_signal_9028 ;
    wire new_AGEMA_signal_9029 ;
    wire new_AGEMA_signal_9030 ;
    wire new_AGEMA_signal_9031 ;
    wire new_AGEMA_signal_9032 ;
    wire new_AGEMA_signal_9033 ;
    wire new_AGEMA_signal_9034 ;
    wire new_AGEMA_signal_9035 ;
    wire new_AGEMA_signal_9036 ;
    wire new_AGEMA_signal_9037 ;
    wire new_AGEMA_signal_9038 ;
    wire new_AGEMA_signal_9039 ;
    wire new_AGEMA_signal_9040 ;
    wire new_AGEMA_signal_9041 ;
    wire new_AGEMA_signal_9042 ;
    wire new_AGEMA_signal_9043 ;
    wire new_AGEMA_signal_9044 ;
    wire new_AGEMA_signal_9045 ;
    wire new_AGEMA_signal_9046 ;
    wire new_AGEMA_signal_9047 ;
    wire new_AGEMA_signal_9048 ;
    wire new_AGEMA_signal_9049 ;
    wire new_AGEMA_signal_9050 ;
    wire new_AGEMA_signal_9051 ;
    wire new_AGEMA_signal_9052 ;
    wire new_AGEMA_signal_9053 ;
    wire new_AGEMA_signal_9054 ;
    wire new_AGEMA_signal_9055 ;
    wire new_AGEMA_signal_9056 ;
    wire new_AGEMA_signal_9057 ;
    wire new_AGEMA_signal_9058 ;
    wire new_AGEMA_signal_9059 ;
    wire new_AGEMA_signal_9060 ;
    wire new_AGEMA_signal_9061 ;
    wire new_AGEMA_signal_9062 ;
    wire new_AGEMA_signal_9063 ;
    wire new_AGEMA_signal_9064 ;
    wire new_AGEMA_signal_9065 ;
    wire new_AGEMA_signal_9066 ;
    wire new_AGEMA_signal_9067 ;
    wire new_AGEMA_signal_9068 ;
    wire new_AGEMA_signal_9069 ;
    wire new_AGEMA_signal_9070 ;
    wire new_AGEMA_signal_9071 ;
    wire new_AGEMA_signal_9072 ;
    wire new_AGEMA_signal_9073 ;
    wire new_AGEMA_signal_9074 ;
    wire new_AGEMA_signal_9075 ;
    wire new_AGEMA_signal_9076 ;
    wire new_AGEMA_signal_9077 ;
    wire new_AGEMA_signal_9078 ;
    wire new_AGEMA_signal_9079 ;
    wire new_AGEMA_signal_9080 ;
    wire new_AGEMA_signal_9081 ;
    wire new_AGEMA_signal_9082 ;
    wire new_AGEMA_signal_9083 ;
    wire new_AGEMA_signal_9084 ;
    wire new_AGEMA_signal_9085 ;
    wire new_AGEMA_signal_9086 ;
    wire new_AGEMA_signal_9087 ;
    wire new_AGEMA_signal_9088 ;
    wire new_AGEMA_signal_9089 ;
    wire new_AGEMA_signal_9090 ;
    wire new_AGEMA_signal_9091 ;
    wire new_AGEMA_signal_9092 ;
    wire new_AGEMA_signal_9093 ;
    wire new_AGEMA_signal_9094 ;
    wire new_AGEMA_signal_9095 ;
    wire new_AGEMA_signal_9096 ;
    wire new_AGEMA_signal_9097 ;
    wire new_AGEMA_signal_9098 ;
    wire new_AGEMA_signal_9099 ;
    wire new_AGEMA_signal_9100 ;
    wire new_AGEMA_signal_9101 ;
    wire new_AGEMA_signal_9102 ;
    wire new_AGEMA_signal_9103 ;
    wire new_AGEMA_signal_9104 ;
    wire new_AGEMA_signal_9105 ;
    wire new_AGEMA_signal_9106 ;
    wire new_AGEMA_signal_9107 ;
    wire new_AGEMA_signal_9108 ;
    wire new_AGEMA_signal_9109 ;
    wire new_AGEMA_signal_9110 ;
    wire new_AGEMA_signal_9111 ;
    wire new_AGEMA_signal_9112 ;
    wire new_AGEMA_signal_9113 ;
    wire new_AGEMA_signal_9114 ;
    wire new_AGEMA_signal_9115 ;
    wire new_AGEMA_signal_9116 ;
    wire new_AGEMA_signal_9117 ;
    wire new_AGEMA_signal_9118 ;
    wire new_AGEMA_signal_9119 ;
    wire new_AGEMA_signal_9120 ;
    wire new_AGEMA_signal_9121 ;
    wire new_AGEMA_signal_9122 ;
    wire new_AGEMA_signal_9123 ;
    wire new_AGEMA_signal_9124 ;
    wire new_AGEMA_signal_9125 ;
    wire new_AGEMA_signal_9126 ;
    wire new_AGEMA_signal_9127 ;
    wire new_AGEMA_signal_9128 ;
    wire new_AGEMA_signal_9129 ;
    wire new_AGEMA_signal_9130 ;
    wire new_AGEMA_signal_9131 ;
    wire new_AGEMA_signal_9132 ;
    wire new_AGEMA_signal_9133 ;
    wire new_AGEMA_signal_9134 ;
    wire new_AGEMA_signal_9135 ;
    wire new_AGEMA_signal_9136 ;
    wire new_AGEMA_signal_9137 ;
    wire new_AGEMA_signal_9138 ;
    wire new_AGEMA_signal_9139 ;
    wire new_AGEMA_signal_9140 ;
    wire new_AGEMA_signal_9141 ;
    wire new_AGEMA_signal_9142 ;
    wire new_AGEMA_signal_9143 ;
    wire new_AGEMA_signal_9144 ;
    wire new_AGEMA_signal_9145 ;
    wire new_AGEMA_signal_9146 ;
    wire new_AGEMA_signal_9147 ;
    wire new_AGEMA_signal_9148 ;
    wire new_AGEMA_signal_9149 ;
    wire new_AGEMA_signal_9150 ;
    wire new_AGEMA_signal_9151 ;
    wire new_AGEMA_signal_9152 ;
    wire new_AGEMA_signal_9153 ;
    wire new_AGEMA_signal_9154 ;
    wire new_AGEMA_signal_9155 ;
    wire new_AGEMA_signal_9156 ;
    wire new_AGEMA_signal_9157 ;
    wire new_AGEMA_signal_9158 ;
    wire new_AGEMA_signal_9159 ;
    wire new_AGEMA_signal_9160 ;
    wire new_AGEMA_signal_9161 ;
    wire new_AGEMA_signal_9162 ;
    wire new_AGEMA_signal_9163 ;
    wire new_AGEMA_signal_9164 ;
    wire new_AGEMA_signal_9165 ;
    wire new_AGEMA_signal_9166 ;
    wire new_AGEMA_signal_9167 ;
    wire new_AGEMA_signal_9168 ;
    wire new_AGEMA_signal_9169 ;
    wire new_AGEMA_signal_9170 ;
    wire new_AGEMA_signal_9171 ;
    wire new_AGEMA_signal_9172 ;
    wire new_AGEMA_signal_9173 ;
    wire new_AGEMA_signal_9174 ;
    wire new_AGEMA_signal_9175 ;
    wire new_AGEMA_signal_9176 ;
    wire new_AGEMA_signal_9177 ;
    wire new_AGEMA_signal_9178 ;
    wire new_AGEMA_signal_9179 ;
    wire new_AGEMA_signal_9180 ;
    wire new_AGEMA_signal_9181 ;
    wire new_AGEMA_signal_9182 ;
    wire new_AGEMA_signal_9183 ;
    wire new_AGEMA_signal_9184 ;
    wire new_AGEMA_signal_9185 ;
    wire new_AGEMA_signal_9186 ;
    wire new_AGEMA_signal_9187 ;
    wire new_AGEMA_signal_9188 ;
    wire new_AGEMA_signal_9189 ;
    wire new_AGEMA_signal_9190 ;
    wire new_AGEMA_signal_9191 ;
    wire new_AGEMA_signal_9192 ;
    wire new_AGEMA_signal_9193 ;
    wire new_AGEMA_signal_9194 ;
    wire new_AGEMA_signal_9195 ;
    wire new_AGEMA_signal_9196 ;
    wire new_AGEMA_signal_9197 ;
    wire new_AGEMA_signal_9198 ;
    wire new_AGEMA_signal_9199 ;
    wire new_AGEMA_signal_9200 ;
    wire new_AGEMA_signal_9201 ;
    wire new_AGEMA_signal_9202 ;
    wire new_AGEMA_signal_9203 ;
    wire new_AGEMA_signal_9204 ;
    wire new_AGEMA_signal_9205 ;
    wire new_AGEMA_signal_9206 ;
    wire new_AGEMA_signal_9207 ;
    wire new_AGEMA_signal_9208 ;
    wire new_AGEMA_signal_9209 ;
    wire new_AGEMA_signal_9210 ;
    wire new_AGEMA_signal_9211 ;
    wire new_AGEMA_signal_9212 ;
    wire new_AGEMA_signal_9213 ;
    wire new_AGEMA_signal_9214 ;
    wire new_AGEMA_signal_9215 ;
    wire new_AGEMA_signal_9216 ;
    wire new_AGEMA_signal_9217 ;
    wire new_AGEMA_signal_9218 ;
    wire new_AGEMA_signal_9219 ;
    wire new_AGEMA_signal_9220 ;
    wire new_AGEMA_signal_9221 ;
    wire new_AGEMA_signal_9222 ;
    wire new_AGEMA_signal_9223 ;
    wire new_AGEMA_signal_9224 ;
    wire new_AGEMA_signal_9225 ;
    wire new_AGEMA_signal_9226 ;
    wire new_AGEMA_signal_9227 ;
    wire new_AGEMA_signal_9228 ;
    wire new_AGEMA_signal_9229 ;
    wire new_AGEMA_signal_9230 ;
    wire new_AGEMA_signal_9231 ;
    wire new_AGEMA_signal_9232 ;
    wire new_AGEMA_signal_9233 ;
    wire new_AGEMA_signal_9234 ;
    wire new_AGEMA_signal_9235 ;
    wire new_AGEMA_signal_9236 ;
    wire new_AGEMA_signal_9237 ;
    wire new_AGEMA_signal_9238 ;
    wire new_AGEMA_signal_9239 ;
    wire new_AGEMA_signal_9240 ;
    wire new_AGEMA_signal_9241 ;
    wire new_AGEMA_signal_9242 ;
    wire new_AGEMA_signal_9243 ;
    wire new_AGEMA_signal_9244 ;
    wire new_AGEMA_signal_9245 ;
    wire new_AGEMA_signal_9246 ;
    wire new_AGEMA_signal_9247 ;
    wire new_AGEMA_signal_9248 ;
    wire new_AGEMA_signal_9249 ;
    wire new_AGEMA_signal_9250 ;
    wire new_AGEMA_signal_9251 ;
    wire new_AGEMA_signal_9252 ;
    wire new_AGEMA_signal_9253 ;
    wire new_AGEMA_signal_9254 ;
    wire new_AGEMA_signal_9255 ;
    wire new_AGEMA_signal_9256 ;
    wire new_AGEMA_signal_9257 ;
    wire new_AGEMA_signal_9258 ;
    wire new_AGEMA_signal_9259 ;
    wire new_AGEMA_signal_9260 ;
    wire new_AGEMA_signal_9261 ;
    wire new_AGEMA_signal_9262 ;
    wire new_AGEMA_signal_9263 ;
    wire new_AGEMA_signal_9264 ;
    wire new_AGEMA_signal_9265 ;
    wire new_AGEMA_signal_9266 ;
    wire new_AGEMA_signal_9267 ;
    wire new_AGEMA_signal_9268 ;
    wire new_AGEMA_signal_9269 ;
    wire new_AGEMA_signal_9270 ;
    wire new_AGEMA_signal_9271 ;
    wire new_AGEMA_signal_9272 ;
    wire new_AGEMA_signal_9273 ;
    wire new_AGEMA_signal_9274 ;
    wire new_AGEMA_signal_9275 ;
    wire new_AGEMA_signal_9276 ;
    wire new_AGEMA_signal_9277 ;
    wire new_AGEMA_signal_9278 ;
    wire new_AGEMA_signal_9279 ;
    wire new_AGEMA_signal_9280 ;
    wire new_AGEMA_signal_9281 ;
    wire new_AGEMA_signal_9282 ;
    wire new_AGEMA_signal_9283 ;
    wire new_AGEMA_signal_9284 ;
    wire new_AGEMA_signal_9285 ;
    wire new_AGEMA_signal_9286 ;
    wire new_AGEMA_signal_9287 ;
    wire new_AGEMA_signal_9288 ;
    wire new_AGEMA_signal_9289 ;
    wire new_AGEMA_signal_9290 ;
    wire new_AGEMA_signal_9291 ;
    wire new_AGEMA_signal_9292 ;
    wire new_AGEMA_signal_9293 ;
    wire new_AGEMA_signal_9294 ;
    wire new_AGEMA_signal_9295 ;
    wire new_AGEMA_signal_9296 ;
    wire new_AGEMA_signal_9297 ;
    wire new_AGEMA_signal_9298 ;
    wire new_AGEMA_signal_9299 ;
    wire new_AGEMA_signal_9300 ;
    wire new_AGEMA_signal_9301 ;
    wire new_AGEMA_signal_9302 ;
    wire new_AGEMA_signal_9303 ;
    wire new_AGEMA_signal_9304 ;
    wire new_AGEMA_signal_9305 ;
    wire new_AGEMA_signal_9306 ;
    wire new_AGEMA_signal_9307 ;
    wire new_AGEMA_signal_9308 ;
    wire new_AGEMA_signal_9309 ;
    wire new_AGEMA_signal_9310 ;
    wire new_AGEMA_signal_9311 ;
    wire new_AGEMA_signal_9312 ;
    wire new_AGEMA_signal_9313 ;
    wire new_AGEMA_signal_9314 ;
    wire new_AGEMA_signal_9315 ;
    wire new_AGEMA_signal_9316 ;
    wire new_AGEMA_signal_9317 ;
    wire new_AGEMA_signal_9318 ;
    wire new_AGEMA_signal_9319 ;
    wire new_AGEMA_signal_9320 ;
    wire new_AGEMA_signal_9321 ;
    wire new_AGEMA_signal_9322 ;
    wire new_AGEMA_signal_9323 ;
    wire new_AGEMA_signal_9324 ;
    wire new_AGEMA_signal_9325 ;
    wire new_AGEMA_signal_9326 ;
    wire new_AGEMA_signal_9327 ;
    wire new_AGEMA_signal_9328 ;
    wire new_AGEMA_signal_9329 ;
    wire new_AGEMA_signal_9330 ;
    wire new_AGEMA_signal_9331 ;
    wire new_AGEMA_signal_9332 ;
    wire new_AGEMA_signal_9333 ;
    wire new_AGEMA_signal_9334 ;
    wire new_AGEMA_signal_9335 ;
    wire new_AGEMA_signal_9336 ;
    wire new_AGEMA_signal_9337 ;
    wire new_AGEMA_signal_9338 ;
    wire new_AGEMA_signal_9339 ;
    wire new_AGEMA_signal_9340 ;
    wire new_AGEMA_signal_9341 ;
    wire new_AGEMA_signal_9342 ;
    wire new_AGEMA_signal_9343 ;
    wire new_AGEMA_signal_9344 ;
    wire new_AGEMA_signal_9345 ;
    wire new_AGEMA_signal_9346 ;
    wire new_AGEMA_signal_9347 ;
    wire new_AGEMA_signal_9348 ;
    wire new_AGEMA_signal_9349 ;
    wire new_AGEMA_signal_9350 ;
    wire new_AGEMA_signal_9351 ;
    wire new_AGEMA_signal_9352 ;
    wire new_AGEMA_signal_9353 ;
    wire new_AGEMA_signal_9354 ;
    wire new_AGEMA_signal_9355 ;
    wire new_AGEMA_signal_9356 ;
    wire new_AGEMA_signal_9357 ;
    wire new_AGEMA_signal_9358 ;
    wire new_AGEMA_signal_9359 ;
    wire new_AGEMA_signal_9360 ;
    wire new_AGEMA_signal_9361 ;
    wire new_AGEMA_signal_9362 ;
    wire new_AGEMA_signal_9363 ;
    wire new_AGEMA_signal_9364 ;
    wire new_AGEMA_signal_9365 ;
    wire new_AGEMA_signal_9366 ;
    wire new_AGEMA_signal_9367 ;
    wire new_AGEMA_signal_9368 ;
    wire new_AGEMA_signal_9369 ;
    wire new_AGEMA_signal_9370 ;
    wire new_AGEMA_signal_9371 ;
    wire new_AGEMA_signal_9372 ;
    wire new_AGEMA_signal_9373 ;
    wire new_AGEMA_signal_9374 ;
    wire new_AGEMA_signal_9375 ;
    wire new_AGEMA_signal_9376 ;
    wire new_AGEMA_signal_9377 ;
    wire new_AGEMA_signal_9378 ;
    wire new_AGEMA_signal_9379 ;
    wire new_AGEMA_signal_9380 ;
    wire new_AGEMA_signal_9381 ;
    wire new_AGEMA_signal_9382 ;
    wire new_AGEMA_signal_9383 ;
    wire new_AGEMA_signal_9384 ;
    wire new_AGEMA_signal_9385 ;
    wire new_AGEMA_signal_9386 ;
    wire new_AGEMA_signal_9387 ;
    wire new_AGEMA_signal_9388 ;
    wire new_AGEMA_signal_9389 ;
    wire new_AGEMA_signal_9390 ;
    wire new_AGEMA_signal_9391 ;
    wire new_AGEMA_signal_9392 ;
    wire new_AGEMA_signal_9393 ;
    wire new_AGEMA_signal_9394 ;
    wire new_AGEMA_signal_9395 ;
    wire new_AGEMA_signal_9396 ;
    wire new_AGEMA_signal_9397 ;
    wire new_AGEMA_signal_9398 ;
    wire new_AGEMA_signal_9399 ;
    wire new_AGEMA_signal_9400 ;
    wire new_AGEMA_signal_9401 ;
    wire new_AGEMA_signal_9402 ;
    wire new_AGEMA_signal_9403 ;
    wire new_AGEMA_signal_9404 ;
    wire new_AGEMA_signal_9405 ;
    wire new_AGEMA_signal_9406 ;
    wire new_AGEMA_signal_9407 ;
    wire new_AGEMA_signal_9408 ;
    wire new_AGEMA_signal_9409 ;
    wire new_AGEMA_signal_9410 ;
    wire new_AGEMA_signal_9411 ;
    wire new_AGEMA_signal_9412 ;
    wire new_AGEMA_signal_9413 ;
    wire new_AGEMA_signal_9414 ;
    wire new_AGEMA_signal_9415 ;
    wire new_AGEMA_signal_9416 ;
    wire new_AGEMA_signal_9417 ;
    wire new_AGEMA_signal_9418 ;
    wire new_AGEMA_signal_9419 ;
    wire new_AGEMA_signal_9420 ;
    wire new_AGEMA_signal_9421 ;
    wire new_AGEMA_signal_9422 ;
    wire new_AGEMA_signal_9423 ;
    wire new_AGEMA_signal_9424 ;
    wire new_AGEMA_signal_9425 ;
    wire new_AGEMA_signal_9426 ;
    wire new_AGEMA_signal_9427 ;
    wire new_AGEMA_signal_9428 ;
    wire new_AGEMA_signal_9429 ;
    wire new_AGEMA_signal_9430 ;
    wire new_AGEMA_signal_9431 ;
    wire new_AGEMA_signal_9432 ;
    wire new_AGEMA_signal_9433 ;
    wire new_AGEMA_signal_9434 ;
    wire new_AGEMA_signal_9435 ;
    wire new_AGEMA_signal_9436 ;
    wire new_AGEMA_signal_9437 ;
    wire new_AGEMA_signal_9438 ;
    wire new_AGEMA_signal_9439 ;
    wire new_AGEMA_signal_9440 ;
    wire new_AGEMA_signal_9441 ;
    wire new_AGEMA_signal_9442 ;
    wire new_AGEMA_signal_9443 ;
    wire new_AGEMA_signal_9444 ;
    wire new_AGEMA_signal_9445 ;
    wire new_AGEMA_signal_9446 ;
    wire new_AGEMA_signal_9447 ;
    wire new_AGEMA_signal_9448 ;
    wire new_AGEMA_signal_9449 ;
    wire new_AGEMA_signal_9450 ;
    wire new_AGEMA_signal_9451 ;
    wire new_AGEMA_signal_9452 ;
    wire new_AGEMA_signal_9453 ;
    wire new_AGEMA_signal_9454 ;
    wire new_AGEMA_signal_9455 ;
    wire new_AGEMA_signal_9456 ;
    wire new_AGEMA_signal_9457 ;
    wire new_AGEMA_signal_9458 ;
    wire new_AGEMA_signal_9459 ;
    wire new_AGEMA_signal_9460 ;
    wire new_AGEMA_signal_9461 ;
    wire new_AGEMA_signal_9462 ;
    wire new_AGEMA_signal_9463 ;
    wire new_AGEMA_signal_9464 ;
    wire new_AGEMA_signal_9465 ;
    wire new_AGEMA_signal_9466 ;
    wire new_AGEMA_signal_9467 ;
    wire new_AGEMA_signal_9468 ;
    wire new_AGEMA_signal_9469 ;
    wire new_AGEMA_signal_9470 ;
    wire new_AGEMA_signal_9471 ;
    wire new_AGEMA_signal_9472 ;
    wire new_AGEMA_signal_9473 ;
    wire new_AGEMA_signal_9474 ;
    wire new_AGEMA_signal_9475 ;
    wire new_AGEMA_signal_9476 ;
    wire new_AGEMA_signal_9477 ;
    wire new_AGEMA_signal_9478 ;
    wire new_AGEMA_signal_9479 ;
    wire new_AGEMA_signal_9480 ;
    wire new_AGEMA_signal_9481 ;
    wire new_AGEMA_signal_9482 ;
    wire new_AGEMA_signal_9483 ;
    wire new_AGEMA_signal_9484 ;
    wire new_AGEMA_signal_9485 ;
    wire new_AGEMA_signal_9486 ;
    wire new_AGEMA_signal_9487 ;
    wire new_AGEMA_signal_9488 ;
    wire new_AGEMA_signal_9489 ;
    wire new_AGEMA_signal_9490 ;
    wire new_AGEMA_signal_9491 ;
    wire new_AGEMA_signal_9492 ;
    wire new_AGEMA_signal_9493 ;
    wire new_AGEMA_signal_9494 ;
    wire new_AGEMA_signal_9495 ;
    wire new_AGEMA_signal_9496 ;
    wire new_AGEMA_signal_9497 ;
    wire new_AGEMA_signal_9498 ;
    wire new_AGEMA_signal_9499 ;
    wire new_AGEMA_signal_9500 ;
    wire new_AGEMA_signal_9501 ;
    wire new_AGEMA_signal_9502 ;
    wire new_AGEMA_signal_9503 ;
    wire new_AGEMA_signal_9504 ;
    wire new_AGEMA_signal_9505 ;
    wire new_AGEMA_signal_9506 ;
    wire new_AGEMA_signal_9507 ;
    wire new_AGEMA_signal_9508 ;
    wire new_AGEMA_signal_9509 ;
    wire new_AGEMA_signal_9510 ;
    wire new_AGEMA_signal_9511 ;
    wire new_AGEMA_signal_9512 ;
    wire new_AGEMA_signal_9513 ;
    wire new_AGEMA_signal_9514 ;
    wire new_AGEMA_signal_9515 ;
    wire new_AGEMA_signal_9516 ;
    wire new_AGEMA_signal_9517 ;
    wire new_AGEMA_signal_9518 ;
    wire new_AGEMA_signal_9519 ;
    wire new_AGEMA_signal_9520 ;
    wire new_AGEMA_signal_9521 ;
    wire new_AGEMA_signal_9522 ;
    wire new_AGEMA_signal_9523 ;
    wire new_AGEMA_signal_9524 ;
    wire new_AGEMA_signal_9525 ;
    wire new_AGEMA_signal_9526 ;
    wire new_AGEMA_signal_9527 ;
    wire new_AGEMA_signal_9528 ;
    wire new_AGEMA_signal_9529 ;
    wire new_AGEMA_signal_9530 ;
    wire new_AGEMA_signal_9531 ;
    wire new_AGEMA_signal_9532 ;
    wire new_AGEMA_signal_9533 ;
    wire new_AGEMA_signal_9534 ;
    wire new_AGEMA_signal_9535 ;
    wire new_AGEMA_signal_9536 ;
    wire new_AGEMA_signal_9537 ;
    wire new_AGEMA_signal_9538 ;
    wire new_AGEMA_signal_9539 ;
    wire new_AGEMA_signal_9540 ;
    wire new_AGEMA_signal_9541 ;
    wire new_AGEMA_signal_9542 ;
    wire new_AGEMA_signal_9543 ;
    wire new_AGEMA_signal_9544 ;
    wire new_AGEMA_signal_9545 ;
    wire new_AGEMA_signal_9546 ;
    wire new_AGEMA_signal_9547 ;
    wire new_AGEMA_signal_9548 ;
    wire new_AGEMA_signal_9549 ;
    wire new_AGEMA_signal_9550 ;
    wire new_AGEMA_signal_9551 ;
    wire new_AGEMA_signal_9552 ;
    wire new_AGEMA_signal_9553 ;
    wire new_AGEMA_signal_9554 ;
    wire new_AGEMA_signal_9555 ;
    wire new_AGEMA_signal_9556 ;
    wire new_AGEMA_signal_9557 ;
    wire new_AGEMA_signal_9558 ;
    wire new_AGEMA_signal_9559 ;
    wire new_AGEMA_signal_9560 ;
    wire new_AGEMA_signal_9561 ;
    wire new_AGEMA_signal_9562 ;
    wire new_AGEMA_signal_9563 ;
    wire new_AGEMA_signal_9564 ;
    wire new_AGEMA_signal_9565 ;
    wire new_AGEMA_signal_9566 ;
    wire new_AGEMA_signal_9567 ;
    wire new_AGEMA_signal_9568 ;
    wire new_AGEMA_signal_9569 ;
    wire new_AGEMA_signal_9570 ;
    wire new_AGEMA_signal_9571 ;
    wire new_AGEMA_signal_9572 ;
    wire new_AGEMA_signal_9573 ;
    wire new_AGEMA_signal_9574 ;
    wire new_AGEMA_signal_9575 ;
    wire new_AGEMA_signal_9576 ;
    wire new_AGEMA_signal_9577 ;
    wire new_AGEMA_signal_9578 ;
    wire new_AGEMA_signal_9579 ;
    wire new_AGEMA_signal_9580 ;
    wire new_AGEMA_signal_9581 ;
    wire new_AGEMA_signal_9582 ;
    wire new_AGEMA_signal_9583 ;
    wire new_AGEMA_signal_9584 ;
    wire new_AGEMA_signal_9585 ;
    wire new_AGEMA_signal_9586 ;
    wire new_AGEMA_signal_9587 ;
    wire new_AGEMA_signal_9588 ;
    wire new_AGEMA_signal_9589 ;
    wire new_AGEMA_signal_9590 ;
    wire new_AGEMA_signal_9591 ;
    wire new_AGEMA_signal_9592 ;
    wire new_AGEMA_signal_9593 ;
    wire new_AGEMA_signal_9594 ;
    wire new_AGEMA_signal_9595 ;
    wire new_AGEMA_signal_9596 ;
    wire new_AGEMA_signal_9597 ;
    wire new_AGEMA_signal_9598 ;
    wire new_AGEMA_signal_9599 ;
    wire new_AGEMA_signal_9600 ;
    wire new_AGEMA_signal_9601 ;
    wire new_AGEMA_signal_9602 ;
    wire new_AGEMA_signal_9603 ;
    wire new_AGEMA_signal_9604 ;
    wire new_AGEMA_signal_9605 ;
    wire new_AGEMA_signal_9606 ;
    wire new_AGEMA_signal_9607 ;
    wire new_AGEMA_signal_9608 ;
    wire new_AGEMA_signal_9609 ;
    wire new_AGEMA_signal_9610 ;
    wire new_AGEMA_signal_9611 ;
    wire new_AGEMA_signal_9612 ;
    wire new_AGEMA_signal_9613 ;
    wire new_AGEMA_signal_9614 ;
    wire new_AGEMA_signal_9615 ;
    wire new_AGEMA_signal_9616 ;
    wire new_AGEMA_signal_9617 ;
    wire new_AGEMA_signal_9618 ;
    wire new_AGEMA_signal_9619 ;
    wire new_AGEMA_signal_9620 ;
    wire new_AGEMA_signal_9621 ;
    wire new_AGEMA_signal_9622 ;
    wire new_AGEMA_signal_9623 ;
    wire new_AGEMA_signal_9624 ;
    wire new_AGEMA_signal_9625 ;
    wire new_AGEMA_signal_9626 ;
    wire new_AGEMA_signal_9627 ;
    wire new_AGEMA_signal_9628 ;
    wire new_AGEMA_signal_9629 ;
    wire new_AGEMA_signal_9630 ;
    wire new_AGEMA_signal_9631 ;
    wire new_AGEMA_signal_9632 ;
    wire new_AGEMA_signal_9633 ;
    wire new_AGEMA_signal_9634 ;
    wire new_AGEMA_signal_9635 ;
    wire new_AGEMA_signal_9636 ;
    wire new_AGEMA_signal_9637 ;
    wire new_AGEMA_signal_9638 ;
    wire new_AGEMA_signal_9639 ;
    wire new_AGEMA_signal_9640 ;
    wire new_AGEMA_signal_9641 ;
    wire new_AGEMA_signal_9642 ;
    wire new_AGEMA_signal_9643 ;
    wire new_AGEMA_signal_9644 ;
    wire new_AGEMA_signal_9645 ;
    wire new_AGEMA_signal_9646 ;
    wire new_AGEMA_signal_9647 ;
    wire new_AGEMA_signal_9648 ;
    wire new_AGEMA_signal_9649 ;
    wire new_AGEMA_signal_9650 ;
    wire new_AGEMA_signal_9651 ;
    wire new_AGEMA_signal_9652 ;
    wire new_AGEMA_signal_9653 ;
    wire new_AGEMA_signal_9654 ;
    wire new_AGEMA_signal_9655 ;
    wire new_AGEMA_signal_9656 ;
    wire new_AGEMA_signal_9657 ;
    wire new_AGEMA_signal_9658 ;
    wire new_AGEMA_signal_9659 ;
    wire new_AGEMA_signal_9660 ;
    wire new_AGEMA_signal_9661 ;
    wire new_AGEMA_signal_9662 ;
    wire new_AGEMA_signal_9663 ;
    wire new_AGEMA_signal_9664 ;
    wire new_AGEMA_signal_9665 ;
    wire new_AGEMA_signal_9666 ;
    wire new_AGEMA_signal_9667 ;
    wire new_AGEMA_signal_9668 ;
    wire new_AGEMA_signal_9669 ;
    wire new_AGEMA_signal_9670 ;
    wire new_AGEMA_signal_9671 ;
    wire new_AGEMA_signal_9672 ;
    wire new_AGEMA_signal_9673 ;
    wire new_AGEMA_signal_9674 ;
    wire new_AGEMA_signal_9675 ;
    wire new_AGEMA_signal_9676 ;
    wire new_AGEMA_signal_9677 ;
    wire new_AGEMA_signal_9678 ;
    wire new_AGEMA_signal_9679 ;
    wire new_AGEMA_signal_9680 ;
    wire new_AGEMA_signal_9681 ;
    wire new_AGEMA_signal_9682 ;
    wire new_AGEMA_signal_9683 ;
    wire new_AGEMA_signal_9684 ;
    wire new_AGEMA_signal_9685 ;
    wire new_AGEMA_signal_9686 ;
    wire new_AGEMA_signal_9687 ;
    wire new_AGEMA_signal_9688 ;
    wire new_AGEMA_signal_9689 ;
    wire new_AGEMA_signal_9690 ;
    wire new_AGEMA_signal_9691 ;
    wire new_AGEMA_signal_9692 ;
    wire new_AGEMA_signal_9693 ;
    wire new_AGEMA_signal_9694 ;
    wire new_AGEMA_signal_9695 ;
    wire new_AGEMA_signal_9696 ;
    wire new_AGEMA_signal_9697 ;
    wire new_AGEMA_signal_9698 ;
    wire new_AGEMA_signal_9699 ;
    wire new_AGEMA_signal_9700 ;
    wire new_AGEMA_signal_9701 ;
    wire new_AGEMA_signal_9702 ;
    wire new_AGEMA_signal_9703 ;
    wire new_AGEMA_signal_9704 ;
    wire new_AGEMA_signal_9705 ;
    wire new_AGEMA_signal_9706 ;
    wire new_AGEMA_signal_9707 ;
    wire new_AGEMA_signal_9708 ;
    wire new_AGEMA_signal_9709 ;
    wire new_AGEMA_signal_9710 ;
    wire new_AGEMA_signal_9711 ;
    wire new_AGEMA_signal_9712 ;
    wire new_AGEMA_signal_9713 ;
    wire new_AGEMA_signal_9714 ;
    wire new_AGEMA_signal_9715 ;
    wire new_AGEMA_signal_9716 ;
    wire new_AGEMA_signal_9717 ;
    wire new_AGEMA_signal_9718 ;
    wire new_AGEMA_signal_9719 ;
    wire new_AGEMA_signal_9720 ;
    wire new_AGEMA_signal_9721 ;
    wire new_AGEMA_signal_9722 ;
    wire new_AGEMA_signal_9723 ;
    wire new_AGEMA_signal_9724 ;
    wire new_AGEMA_signal_9725 ;
    wire new_AGEMA_signal_9726 ;
    wire new_AGEMA_signal_9727 ;
    wire new_AGEMA_signal_9728 ;
    wire new_AGEMA_signal_9729 ;
    wire new_AGEMA_signal_9730 ;
    wire new_AGEMA_signal_9731 ;
    wire new_AGEMA_signal_9732 ;
    wire new_AGEMA_signal_9733 ;
    wire new_AGEMA_signal_9734 ;
    wire new_AGEMA_signal_9735 ;
    wire new_AGEMA_signal_9736 ;
    wire new_AGEMA_signal_9737 ;
    wire new_AGEMA_signal_9738 ;
    wire new_AGEMA_signal_9739 ;
    wire new_AGEMA_signal_9740 ;
    wire new_AGEMA_signal_9741 ;
    wire new_AGEMA_signal_9742 ;
    wire new_AGEMA_signal_9743 ;
    wire new_AGEMA_signal_9744 ;
    wire new_AGEMA_signal_9745 ;
    wire new_AGEMA_signal_9746 ;
    wire new_AGEMA_signal_9747 ;
    wire new_AGEMA_signal_9748 ;
    wire new_AGEMA_signal_9749 ;
    wire new_AGEMA_signal_9750 ;
    wire new_AGEMA_signal_9751 ;
    wire new_AGEMA_signal_9752 ;
    wire new_AGEMA_signal_9753 ;
    wire new_AGEMA_signal_9754 ;
    wire new_AGEMA_signal_9755 ;
    wire new_AGEMA_signal_9756 ;
    wire new_AGEMA_signal_9757 ;
    wire new_AGEMA_signal_9758 ;
    wire new_AGEMA_signal_9759 ;
    wire new_AGEMA_signal_9760 ;
    wire new_AGEMA_signal_9761 ;
    wire new_AGEMA_signal_9762 ;
    wire new_AGEMA_signal_9763 ;
    wire new_AGEMA_signal_9764 ;
    wire new_AGEMA_signal_9765 ;
    wire new_AGEMA_signal_9766 ;
    wire new_AGEMA_signal_9767 ;
    wire new_AGEMA_signal_9768 ;
    wire new_AGEMA_signal_9769 ;
    wire new_AGEMA_signal_9770 ;
    wire new_AGEMA_signal_9771 ;
    wire new_AGEMA_signal_9772 ;
    wire new_AGEMA_signal_9773 ;
    wire new_AGEMA_signal_9774 ;
    wire new_AGEMA_signal_9775 ;
    wire new_AGEMA_signal_9776 ;
    wire new_AGEMA_signal_9777 ;
    wire new_AGEMA_signal_9778 ;
    wire new_AGEMA_signal_9779 ;
    wire new_AGEMA_signal_9780 ;
    wire new_AGEMA_signal_9781 ;
    wire new_AGEMA_signal_9782 ;
    wire new_AGEMA_signal_9783 ;
    wire new_AGEMA_signal_9784 ;
    wire new_AGEMA_signal_9785 ;
    wire new_AGEMA_signal_9786 ;
    wire new_AGEMA_signal_9787 ;
    wire new_AGEMA_signal_9788 ;
    wire new_AGEMA_signal_9789 ;
    wire new_AGEMA_signal_9790 ;
    wire new_AGEMA_signal_9791 ;
    wire new_AGEMA_signal_9792 ;
    wire new_AGEMA_signal_9793 ;
    wire new_AGEMA_signal_9794 ;
    wire new_AGEMA_signal_9795 ;
    wire new_AGEMA_signal_9796 ;
    wire new_AGEMA_signal_9797 ;
    wire new_AGEMA_signal_9798 ;
    wire new_AGEMA_signal_9799 ;
    wire new_AGEMA_signal_9800 ;
    wire new_AGEMA_signal_9801 ;
    wire new_AGEMA_signal_9802 ;
    wire new_AGEMA_signal_9803 ;
    wire new_AGEMA_signal_9804 ;
    wire new_AGEMA_signal_9805 ;
    wire new_AGEMA_signal_9806 ;
    wire new_AGEMA_signal_9807 ;
    wire new_AGEMA_signal_9808 ;
    wire new_AGEMA_signal_9809 ;
    wire new_AGEMA_signal_9810 ;
    wire new_AGEMA_signal_9811 ;
    wire new_AGEMA_signal_9812 ;
    wire new_AGEMA_signal_9813 ;
    wire new_AGEMA_signal_9814 ;
    wire new_AGEMA_signal_9815 ;
    wire new_AGEMA_signal_9816 ;
    wire new_AGEMA_signal_9817 ;
    wire new_AGEMA_signal_9818 ;
    wire new_AGEMA_signal_9819 ;
    wire new_AGEMA_signal_9820 ;
    wire new_AGEMA_signal_9821 ;
    wire new_AGEMA_signal_9822 ;
    wire new_AGEMA_signal_9823 ;
    wire new_AGEMA_signal_9824 ;
    wire new_AGEMA_signal_9825 ;
    wire new_AGEMA_signal_9826 ;
    wire new_AGEMA_signal_9827 ;
    wire new_AGEMA_signal_9828 ;
    wire new_AGEMA_signal_9829 ;
    wire new_AGEMA_signal_9830 ;
    wire new_AGEMA_signal_9831 ;
    wire new_AGEMA_signal_9832 ;
    wire new_AGEMA_signal_9833 ;
    wire new_AGEMA_signal_9834 ;
    wire new_AGEMA_signal_9835 ;
    wire new_AGEMA_signal_9836 ;
    wire new_AGEMA_signal_9837 ;
    wire new_AGEMA_signal_9838 ;
    wire new_AGEMA_signal_9839 ;
    wire new_AGEMA_signal_9840 ;
    wire new_AGEMA_signal_9841 ;
    wire new_AGEMA_signal_9842 ;
    wire new_AGEMA_signal_9843 ;
    wire new_AGEMA_signal_9844 ;
    wire new_AGEMA_signal_9845 ;
    wire new_AGEMA_signal_9846 ;
    wire new_AGEMA_signal_9847 ;
    wire new_AGEMA_signal_9848 ;
    wire new_AGEMA_signal_9849 ;
    wire new_AGEMA_signal_9850 ;
    wire new_AGEMA_signal_9851 ;
    wire new_AGEMA_signal_9852 ;
    wire new_AGEMA_signal_9853 ;
    wire new_AGEMA_signal_9854 ;
    wire new_AGEMA_signal_9855 ;
    wire new_AGEMA_signal_9856 ;
    wire new_AGEMA_signal_9857 ;
    wire new_AGEMA_signal_9858 ;
    wire new_AGEMA_signal_9859 ;
    wire new_AGEMA_signal_9860 ;
    wire new_AGEMA_signal_9861 ;
    wire new_AGEMA_signal_9862 ;
    wire new_AGEMA_signal_9863 ;
    wire new_AGEMA_signal_9864 ;
    wire new_AGEMA_signal_9865 ;
    wire new_AGEMA_signal_9866 ;
    wire new_AGEMA_signal_9867 ;
    wire new_AGEMA_signal_9868 ;
    wire new_AGEMA_signal_9869 ;
    wire new_AGEMA_signal_9870 ;
    wire new_AGEMA_signal_9871 ;
    wire new_AGEMA_signal_9872 ;
    wire new_AGEMA_signal_9873 ;
    wire new_AGEMA_signal_9874 ;
    wire new_AGEMA_signal_9875 ;
    wire new_AGEMA_signal_9876 ;
    wire new_AGEMA_signal_9877 ;
    wire new_AGEMA_signal_9878 ;
    wire new_AGEMA_signal_9879 ;
    wire new_AGEMA_signal_9880 ;
    wire new_AGEMA_signal_9881 ;
    wire new_AGEMA_signal_9882 ;
    wire new_AGEMA_signal_9883 ;
    wire new_AGEMA_signal_9884 ;
    wire new_AGEMA_signal_9885 ;
    wire new_AGEMA_signal_9886 ;
    wire new_AGEMA_signal_9887 ;
    wire new_AGEMA_signal_9888 ;
    wire new_AGEMA_signal_9889 ;
    wire new_AGEMA_signal_9890 ;
    wire new_AGEMA_signal_9891 ;
    wire new_AGEMA_signal_9892 ;
    wire new_AGEMA_signal_9893 ;
    wire new_AGEMA_signal_9894 ;
    wire new_AGEMA_signal_9895 ;
    wire new_AGEMA_signal_9896 ;
    wire new_AGEMA_signal_9897 ;
    wire new_AGEMA_signal_9898 ;
    wire new_AGEMA_signal_9899 ;
    wire new_AGEMA_signal_9900 ;
    wire new_AGEMA_signal_9901 ;
    wire new_AGEMA_signal_9902 ;
    wire new_AGEMA_signal_9903 ;
    wire new_AGEMA_signal_9904 ;
    wire new_AGEMA_signal_9905 ;
    wire new_AGEMA_signal_9906 ;
    wire new_AGEMA_signal_9907 ;
    wire new_AGEMA_signal_9908 ;
    wire new_AGEMA_signal_9909 ;
    wire new_AGEMA_signal_9910 ;
    wire new_AGEMA_signal_9911 ;
    wire new_AGEMA_signal_9912 ;
    wire new_AGEMA_signal_9913 ;
    wire new_AGEMA_signal_9914 ;
    wire new_AGEMA_signal_9915 ;
    wire new_AGEMA_signal_9916 ;
    wire new_AGEMA_signal_9917 ;
    wire new_AGEMA_signal_9918 ;
    wire new_AGEMA_signal_9919 ;
    wire new_AGEMA_signal_9920 ;
    wire new_AGEMA_signal_9921 ;
    wire new_AGEMA_signal_9922 ;
    wire new_AGEMA_signal_9923 ;
    wire new_AGEMA_signal_9924 ;
    wire new_AGEMA_signal_9925 ;
    wire new_AGEMA_signal_9926 ;
    wire new_AGEMA_signal_9927 ;
    wire new_AGEMA_signal_9928 ;
    wire new_AGEMA_signal_9929 ;
    wire new_AGEMA_signal_9930 ;
    wire new_AGEMA_signal_9931 ;
    wire new_AGEMA_signal_9932 ;
    wire new_AGEMA_signal_9933 ;
    wire new_AGEMA_signal_9934 ;
    wire new_AGEMA_signal_9935 ;
    wire new_AGEMA_signal_9936 ;
    wire new_AGEMA_signal_9937 ;
    wire new_AGEMA_signal_9938 ;
    wire new_AGEMA_signal_9939 ;
    wire new_AGEMA_signal_9940 ;
    wire new_AGEMA_signal_9941 ;
    wire new_AGEMA_signal_9942 ;
    wire new_AGEMA_signal_9943 ;
    wire new_AGEMA_signal_9944 ;
    wire new_AGEMA_signal_9945 ;
    wire new_AGEMA_signal_9946 ;
    wire new_AGEMA_signal_9947 ;
    wire new_AGEMA_signal_9948 ;
    wire new_AGEMA_signal_9949 ;
    wire new_AGEMA_signal_9950 ;
    wire new_AGEMA_signal_9951 ;
    wire new_AGEMA_signal_9952 ;
    wire new_AGEMA_signal_9953 ;
    wire new_AGEMA_signal_9954 ;
    wire new_AGEMA_signal_9955 ;
    wire new_AGEMA_signal_9956 ;
    wire new_AGEMA_signal_9957 ;
    wire new_AGEMA_signal_9958 ;
    wire new_AGEMA_signal_9959 ;
    wire new_AGEMA_signal_9960 ;
    wire new_AGEMA_signal_9961 ;
    wire new_AGEMA_signal_9962 ;
    wire new_AGEMA_signal_9963 ;
    wire new_AGEMA_signal_9964 ;
    wire new_AGEMA_signal_9965 ;
    wire new_AGEMA_signal_9966 ;
    wire new_AGEMA_signal_9967 ;
    wire new_AGEMA_signal_9968 ;
    wire new_AGEMA_signal_9969 ;
    wire new_AGEMA_signal_9970 ;
    wire new_AGEMA_signal_9971 ;
    wire new_AGEMA_signal_9972 ;
    wire new_AGEMA_signal_9973 ;
    wire new_AGEMA_signal_9974 ;
    wire new_AGEMA_signal_9975 ;
    wire new_AGEMA_signal_9976 ;
    wire new_AGEMA_signal_9977 ;
    wire new_AGEMA_signal_9978 ;
    wire new_AGEMA_signal_9979 ;
    wire new_AGEMA_signal_9980 ;
    wire new_AGEMA_signal_9981 ;
    wire new_AGEMA_signal_9982 ;
    wire new_AGEMA_signal_9983 ;
    wire new_AGEMA_signal_9984 ;
    wire new_AGEMA_signal_9985 ;
    wire new_AGEMA_signal_9986 ;
    wire new_AGEMA_signal_9987 ;
    wire new_AGEMA_signal_9988 ;
    wire new_AGEMA_signal_9989 ;
    wire new_AGEMA_signal_9990 ;
    wire new_AGEMA_signal_9991 ;
    wire new_AGEMA_signal_9992 ;
    wire new_AGEMA_signal_9993 ;
    wire new_AGEMA_signal_9994 ;
    wire new_AGEMA_signal_9995 ;
    wire new_AGEMA_signal_9996 ;
    wire new_AGEMA_signal_9997 ;
    wire new_AGEMA_signal_9998 ;
    wire new_AGEMA_signal_9999 ;
    wire new_AGEMA_signal_10000 ;
    wire new_AGEMA_signal_10001 ;
    wire new_AGEMA_signal_10002 ;
    wire new_AGEMA_signal_10003 ;
    wire new_AGEMA_signal_10004 ;
    wire new_AGEMA_signal_10005 ;
    wire new_AGEMA_signal_10006 ;
    wire new_AGEMA_signal_10007 ;
    wire new_AGEMA_signal_10008 ;
    wire new_AGEMA_signal_10009 ;
    wire new_AGEMA_signal_10010 ;
    wire new_AGEMA_signal_10011 ;
    wire new_AGEMA_signal_10012 ;
    wire new_AGEMA_signal_10013 ;
    wire new_AGEMA_signal_10014 ;
    wire new_AGEMA_signal_10015 ;
    wire new_AGEMA_signal_10016 ;
    wire new_AGEMA_signal_10017 ;
    wire new_AGEMA_signal_10018 ;
    wire new_AGEMA_signal_10019 ;
    wire new_AGEMA_signal_10020 ;
    wire new_AGEMA_signal_10021 ;
    wire new_AGEMA_signal_10022 ;
    wire new_AGEMA_signal_10023 ;
    wire new_AGEMA_signal_10024 ;
    wire new_AGEMA_signal_10025 ;
    wire new_AGEMA_signal_10026 ;
    wire new_AGEMA_signal_10027 ;
    wire new_AGEMA_signal_10028 ;
    wire new_AGEMA_signal_10029 ;
    wire new_AGEMA_signal_10030 ;
    wire new_AGEMA_signal_10031 ;
    wire new_AGEMA_signal_10032 ;
    wire new_AGEMA_signal_10033 ;
    wire new_AGEMA_signal_10034 ;
    wire new_AGEMA_signal_10035 ;
    wire new_AGEMA_signal_10036 ;
    wire new_AGEMA_signal_10037 ;
    wire new_AGEMA_signal_10038 ;
    wire new_AGEMA_signal_10039 ;
    wire new_AGEMA_signal_10040 ;
    wire new_AGEMA_signal_10041 ;
    wire new_AGEMA_signal_10042 ;
    wire new_AGEMA_signal_10043 ;
    wire new_AGEMA_signal_10044 ;
    wire new_AGEMA_signal_10045 ;
    wire new_AGEMA_signal_10046 ;
    wire new_AGEMA_signal_10047 ;
    wire new_AGEMA_signal_10048 ;
    wire new_AGEMA_signal_10049 ;
    wire new_AGEMA_signal_10050 ;
    wire new_AGEMA_signal_10051 ;
    wire new_AGEMA_signal_10052 ;
    wire new_AGEMA_signal_10053 ;
    wire new_AGEMA_signal_10054 ;
    wire new_AGEMA_signal_10055 ;
    wire new_AGEMA_signal_10056 ;
    wire new_AGEMA_signal_10057 ;
    wire new_AGEMA_signal_10058 ;
    wire new_AGEMA_signal_10059 ;
    wire new_AGEMA_signal_10060 ;
    wire new_AGEMA_signal_10061 ;
    wire new_AGEMA_signal_10062 ;
    wire new_AGEMA_signal_10063 ;
    wire new_AGEMA_signal_10064 ;
    wire new_AGEMA_signal_10065 ;
    wire new_AGEMA_signal_10066 ;
    wire new_AGEMA_signal_10067 ;
    wire new_AGEMA_signal_10068 ;
    wire new_AGEMA_signal_10069 ;
    wire new_AGEMA_signal_10070 ;
    wire new_AGEMA_signal_10071 ;
    wire new_AGEMA_signal_10072 ;
    wire new_AGEMA_signal_10073 ;
    wire new_AGEMA_signal_10074 ;
    wire new_AGEMA_signal_10075 ;
    wire new_AGEMA_signal_10076 ;
    wire new_AGEMA_signal_10077 ;
    wire new_AGEMA_signal_10078 ;
    wire new_AGEMA_signal_10079 ;
    wire new_AGEMA_signal_10080 ;
    wire new_AGEMA_signal_10081 ;
    wire new_AGEMA_signal_10082 ;
    wire new_AGEMA_signal_10083 ;
    wire new_AGEMA_signal_10084 ;
    wire new_AGEMA_signal_10085 ;
    wire new_AGEMA_signal_10086 ;
    wire new_AGEMA_signal_10087 ;
    wire new_AGEMA_signal_10088 ;
    wire new_AGEMA_signal_10089 ;
    wire new_AGEMA_signal_10090 ;
    wire new_AGEMA_signal_10091 ;
    wire new_AGEMA_signal_10092 ;
    wire new_AGEMA_signal_10093 ;
    wire new_AGEMA_signal_10094 ;
    wire new_AGEMA_signal_10095 ;
    wire new_AGEMA_signal_10096 ;
    wire new_AGEMA_signal_10097 ;
    wire new_AGEMA_signal_10098 ;
    wire new_AGEMA_signal_10099 ;
    wire new_AGEMA_signal_10100 ;
    wire new_AGEMA_signal_10101 ;
    wire new_AGEMA_signal_10102 ;
    wire new_AGEMA_signal_10103 ;
    wire new_AGEMA_signal_10104 ;
    wire new_AGEMA_signal_10105 ;
    wire new_AGEMA_signal_10106 ;
    wire new_AGEMA_signal_10107 ;
    wire new_AGEMA_signal_10108 ;
    wire new_AGEMA_signal_10109 ;
    wire new_AGEMA_signal_10110 ;
    wire new_AGEMA_signal_10111 ;
    wire new_AGEMA_signal_10112 ;
    wire new_AGEMA_signal_10113 ;
    wire new_AGEMA_signal_10114 ;
    wire new_AGEMA_signal_10115 ;
    wire new_AGEMA_signal_10116 ;
    wire new_AGEMA_signal_10117 ;
    wire new_AGEMA_signal_10118 ;
    wire new_AGEMA_signal_10119 ;
    wire new_AGEMA_signal_10120 ;
    wire new_AGEMA_signal_10121 ;
    wire new_AGEMA_signal_10122 ;
    wire new_AGEMA_signal_10123 ;
    wire new_AGEMA_signal_10124 ;
    wire new_AGEMA_signal_10125 ;
    wire new_AGEMA_signal_10126 ;
    wire new_AGEMA_signal_10127 ;
    wire new_AGEMA_signal_10128 ;
    wire new_AGEMA_signal_10129 ;
    wire new_AGEMA_signal_10130 ;
    wire new_AGEMA_signal_10131 ;
    wire new_AGEMA_signal_10132 ;
    wire new_AGEMA_signal_10133 ;
    wire new_AGEMA_signal_10134 ;
    wire new_AGEMA_signal_10135 ;
    wire new_AGEMA_signal_10136 ;
    wire new_AGEMA_signal_10137 ;
    wire new_AGEMA_signal_10138 ;
    wire new_AGEMA_signal_10139 ;
    wire new_AGEMA_signal_10140 ;
    wire new_AGEMA_signal_10141 ;
    wire new_AGEMA_signal_10142 ;
    wire new_AGEMA_signal_10143 ;
    wire new_AGEMA_signal_10144 ;
    wire new_AGEMA_signal_10145 ;
    wire new_AGEMA_signal_10146 ;
    wire new_AGEMA_signal_10147 ;
    wire new_AGEMA_signal_10148 ;
    wire new_AGEMA_signal_10149 ;
    wire new_AGEMA_signal_10150 ;
    wire new_AGEMA_signal_10151 ;
    wire new_AGEMA_signal_10152 ;
    wire new_AGEMA_signal_10153 ;
    wire new_AGEMA_signal_10154 ;
    wire new_AGEMA_signal_10155 ;
    wire new_AGEMA_signal_10156 ;
    wire new_AGEMA_signal_10157 ;
    wire new_AGEMA_signal_10158 ;
    wire new_AGEMA_signal_10159 ;
    wire new_AGEMA_signal_10160 ;
    wire new_AGEMA_signal_10161 ;
    wire new_AGEMA_signal_10162 ;
    wire new_AGEMA_signal_10163 ;
    wire new_AGEMA_signal_10164 ;
    wire new_AGEMA_signal_10165 ;
    wire new_AGEMA_signal_10166 ;
    wire new_AGEMA_signal_10167 ;
    wire new_AGEMA_signal_10168 ;
    wire new_AGEMA_signal_10169 ;
    wire new_AGEMA_signal_10170 ;
    wire new_AGEMA_signal_10171 ;
    wire new_AGEMA_signal_10172 ;
    wire new_AGEMA_signal_10173 ;
    wire new_AGEMA_signal_10174 ;
    wire new_AGEMA_signal_10175 ;
    wire new_AGEMA_signal_10176 ;
    wire new_AGEMA_signal_10177 ;
    wire new_AGEMA_signal_10178 ;
    wire new_AGEMA_signal_10179 ;
    wire new_AGEMA_signal_10180 ;
    wire new_AGEMA_signal_10181 ;
    wire new_AGEMA_signal_10182 ;
    wire new_AGEMA_signal_10183 ;
    wire new_AGEMA_signal_10184 ;
    wire new_AGEMA_signal_10185 ;
    wire new_AGEMA_signal_10186 ;
    wire new_AGEMA_signal_10187 ;
    wire new_AGEMA_signal_10188 ;
    wire new_AGEMA_signal_10189 ;
    wire new_AGEMA_signal_10190 ;
    wire new_AGEMA_signal_10191 ;
    wire new_AGEMA_signal_10192 ;
    wire new_AGEMA_signal_10193 ;
    wire new_AGEMA_signal_10194 ;
    wire new_AGEMA_signal_10195 ;
    wire new_AGEMA_signal_10196 ;
    wire new_AGEMA_signal_10197 ;
    wire new_AGEMA_signal_10198 ;
    wire new_AGEMA_signal_10199 ;
    wire new_AGEMA_signal_10200 ;
    wire new_AGEMA_signal_10201 ;
    wire new_AGEMA_signal_10202 ;
    wire new_AGEMA_signal_10203 ;
    wire new_AGEMA_signal_10204 ;
    wire new_AGEMA_signal_10205 ;
    wire new_AGEMA_signal_10206 ;
    wire new_AGEMA_signal_10207 ;
    wire new_AGEMA_signal_10208 ;
    wire new_AGEMA_signal_10209 ;
    wire new_AGEMA_signal_10210 ;
    wire new_AGEMA_signal_10211 ;
    wire new_AGEMA_signal_10212 ;
    wire new_AGEMA_signal_10213 ;
    wire new_AGEMA_signal_10214 ;
    wire new_AGEMA_signal_10215 ;
    wire new_AGEMA_signal_10216 ;
    wire new_AGEMA_signal_10217 ;
    wire new_AGEMA_signal_10218 ;
    wire new_AGEMA_signal_10219 ;
    wire new_AGEMA_signal_10220 ;
    wire new_AGEMA_signal_10221 ;
    wire new_AGEMA_signal_10222 ;
    wire new_AGEMA_signal_10223 ;
    wire new_AGEMA_signal_10224 ;
    wire new_AGEMA_signal_10225 ;
    wire new_AGEMA_signal_10226 ;
    wire new_AGEMA_signal_10227 ;
    wire new_AGEMA_signal_10228 ;
    wire new_AGEMA_signal_10229 ;
    wire new_AGEMA_signal_10230 ;
    wire new_AGEMA_signal_10231 ;
    wire new_AGEMA_signal_10232 ;
    wire new_AGEMA_signal_10233 ;
    wire new_AGEMA_signal_10234 ;
    wire new_AGEMA_signal_10235 ;
    wire new_AGEMA_signal_10236 ;
    wire new_AGEMA_signal_10237 ;
    wire new_AGEMA_signal_10238 ;
    wire new_AGEMA_signal_10239 ;
    wire new_AGEMA_signal_10240 ;
    wire new_AGEMA_signal_10241 ;
    wire new_AGEMA_signal_10242 ;
    wire new_AGEMA_signal_10243 ;
    wire new_AGEMA_signal_10244 ;
    wire new_AGEMA_signal_10245 ;
    wire new_AGEMA_signal_10246 ;
    wire new_AGEMA_signal_10247 ;
    wire new_AGEMA_signal_10248 ;
    wire new_AGEMA_signal_10249 ;
    wire new_AGEMA_signal_10250 ;
    wire new_AGEMA_signal_10251 ;
    wire new_AGEMA_signal_10252 ;
    wire new_AGEMA_signal_10253 ;
    wire new_AGEMA_signal_10254 ;
    wire new_AGEMA_signal_10255 ;
    wire new_AGEMA_signal_10256 ;
    wire new_AGEMA_signal_10257 ;
    wire new_AGEMA_signal_10258 ;
    wire new_AGEMA_signal_10259 ;
    wire new_AGEMA_signal_10260 ;
    wire new_AGEMA_signal_10261 ;
    wire new_AGEMA_signal_10262 ;
    wire new_AGEMA_signal_10263 ;
    wire new_AGEMA_signal_10264 ;
    wire new_AGEMA_signal_10265 ;
    wire new_AGEMA_signal_10266 ;
    wire new_AGEMA_signal_10267 ;
    wire new_AGEMA_signal_10268 ;
    wire new_AGEMA_signal_10269 ;
    wire new_AGEMA_signal_10270 ;
    wire new_AGEMA_signal_10271 ;
    wire new_AGEMA_signal_10272 ;
    wire new_AGEMA_signal_10273 ;
    wire new_AGEMA_signal_10274 ;
    wire new_AGEMA_signal_10275 ;
    wire new_AGEMA_signal_10276 ;
    wire new_AGEMA_signal_10277 ;
    wire new_AGEMA_signal_10278 ;
    wire new_AGEMA_signal_10279 ;
    wire new_AGEMA_signal_10280 ;
    wire new_AGEMA_signal_10281 ;
    wire new_AGEMA_signal_10282 ;
    wire new_AGEMA_signal_10283 ;
    wire new_AGEMA_signal_10284 ;
    wire new_AGEMA_signal_10285 ;
    wire new_AGEMA_signal_10286 ;
    wire new_AGEMA_signal_10287 ;
    wire new_AGEMA_signal_10288 ;
    wire new_AGEMA_signal_10289 ;
    wire new_AGEMA_signal_10290 ;
    wire new_AGEMA_signal_10291 ;
    wire new_AGEMA_signal_10292 ;
    wire new_AGEMA_signal_10293 ;
    wire new_AGEMA_signal_10294 ;
    wire new_AGEMA_signal_10295 ;
    wire new_AGEMA_signal_10296 ;
    wire new_AGEMA_signal_10297 ;
    wire new_AGEMA_signal_10298 ;
    wire new_AGEMA_signal_10299 ;
    wire new_AGEMA_signal_10300 ;
    wire new_AGEMA_signal_10301 ;
    wire new_AGEMA_signal_10302 ;
    wire new_AGEMA_signal_10303 ;
    wire new_AGEMA_signal_10304 ;
    wire new_AGEMA_signal_10305 ;
    wire new_AGEMA_signal_10306 ;
    wire new_AGEMA_signal_10307 ;
    wire new_AGEMA_signal_10308 ;
    wire new_AGEMA_signal_10309 ;
    wire new_AGEMA_signal_10310 ;
    wire new_AGEMA_signal_10311 ;
    wire new_AGEMA_signal_10312 ;
    wire new_AGEMA_signal_10313 ;
    wire new_AGEMA_signal_10314 ;
    wire new_AGEMA_signal_10315 ;
    wire new_AGEMA_signal_10316 ;
    wire new_AGEMA_signal_10317 ;
    wire new_AGEMA_signal_10318 ;
    wire new_AGEMA_signal_10319 ;
    wire new_AGEMA_signal_10320 ;
    wire new_AGEMA_signal_10321 ;
    wire new_AGEMA_signal_10322 ;
    wire new_AGEMA_signal_10323 ;
    wire new_AGEMA_signal_10324 ;
    wire new_AGEMA_signal_10325 ;
    wire new_AGEMA_signal_10326 ;
    wire new_AGEMA_signal_10327 ;
    wire new_AGEMA_signal_10328 ;
    wire new_AGEMA_signal_10329 ;
    wire new_AGEMA_signal_10330 ;
    wire new_AGEMA_signal_10331 ;
    wire new_AGEMA_signal_10332 ;
    wire new_AGEMA_signal_10333 ;
    wire new_AGEMA_signal_10334 ;
    wire new_AGEMA_signal_10335 ;
    wire new_AGEMA_signal_10336 ;
    wire new_AGEMA_signal_10337 ;
    wire new_AGEMA_signal_10338 ;
    wire new_AGEMA_signal_10339 ;
    wire new_AGEMA_signal_10340 ;
    wire new_AGEMA_signal_10341 ;
    wire new_AGEMA_signal_10342 ;
    wire new_AGEMA_signal_10343 ;
    wire new_AGEMA_signal_10344 ;
    wire new_AGEMA_signal_10345 ;
    wire new_AGEMA_signal_10346 ;
    wire new_AGEMA_signal_10347 ;
    wire new_AGEMA_signal_10348 ;
    wire new_AGEMA_signal_10349 ;
    wire new_AGEMA_signal_10350 ;
    wire new_AGEMA_signal_10351 ;
    wire new_AGEMA_signal_10352 ;
    wire new_AGEMA_signal_10353 ;
    wire new_AGEMA_signal_10354 ;
    wire new_AGEMA_signal_10355 ;
    wire new_AGEMA_signal_10356 ;
    wire new_AGEMA_signal_10357 ;
    wire new_AGEMA_signal_10358 ;
    wire new_AGEMA_signal_10359 ;
    wire new_AGEMA_signal_10360 ;
    wire new_AGEMA_signal_10361 ;
    wire new_AGEMA_signal_10362 ;
    wire new_AGEMA_signal_10363 ;
    wire new_AGEMA_signal_10364 ;
    wire new_AGEMA_signal_10365 ;
    wire new_AGEMA_signal_10366 ;
    wire new_AGEMA_signal_10367 ;
    wire new_AGEMA_signal_10368 ;
    wire new_AGEMA_signal_10369 ;
    wire new_AGEMA_signal_10370 ;
    wire new_AGEMA_signal_10371 ;
    wire new_AGEMA_signal_10372 ;
    wire new_AGEMA_signal_10373 ;
    wire new_AGEMA_signal_10374 ;
    wire new_AGEMA_signal_10375 ;
    wire new_AGEMA_signal_10376 ;
    wire new_AGEMA_signal_10377 ;
    wire new_AGEMA_signal_10378 ;
    wire new_AGEMA_signal_10379 ;
    wire new_AGEMA_signal_10380 ;
    wire new_AGEMA_signal_10381 ;
    wire new_AGEMA_signal_10382 ;
    wire new_AGEMA_signal_10383 ;
    wire new_AGEMA_signal_10384 ;
    wire new_AGEMA_signal_10385 ;
    wire new_AGEMA_signal_10386 ;
    wire new_AGEMA_signal_10387 ;
    wire new_AGEMA_signal_10388 ;
    wire new_AGEMA_signal_10389 ;
    wire new_AGEMA_signal_10390 ;
    wire new_AGEMA_signal_10391 ;
    wire new_AGEMA_signal_10392 ;
    wire new_AGEMA_signal_10393 ;
    wire new_AGEMA_signal_10394 ;
    wire new_AGEMA_signal_10395 ;
    wire new_AGEMA_signal_10396 ;
    wire new_AGEMA_signal_10397 ;
    wire new_AGEMA_signal_10398 ;
    wire new_AGEMA_signal_10399 ;
    wire new_AGEMA_signal_10400 ;
    wire new_AGEMA_signal_10401 ;
    wire new_AGEMA_signal_10402 ;
    wire new_AGEMA_signal_10403 ;
    wire new_AGEMA_signal_10404 ;
    wire new_AGEMA_signal_10405 ;
    wire new_AGEMA_signal_10406 ;
    wire new_AGEMA_signal_10407 ;
    wire new_AGEMA_signal_10408 ;
    wire new_AGEMA_signal_10409 ;
    wire new_AGEMA_signal_10410 ;
    wire new_AGEMA_signal_10411 ;
    wire new_AGEMA_signal_10412 ;
    wire new_AGEMA_signal_10413 ;
    wire new_AGEMA_signal_10414 ;
    wire new_AGEMA_signal_10415 ;
    wire new_AGEMA_signal_10416 ;
    wire new_AGEMA_signal_10417 ;
    wire new_AGEMA_signal_10418 ;
    wire new_AGEMA_signal_10419 ;
    wire new_AGEMA_signal_10420 ;
    wire new_AGEMA_signal_10421 ;
    wire new_AGEMA_signal_10422 ;
    wire new_AGEMA_signal_10423 ;
    wire new_AGEMA_signal_10424 ;
    wire new_AGEMA_signal_10425 ;
    wire new_AGEMA_signal_10426 ;
    wire new_AGEMA_signal_10427 ;
    wire new_AGEMA_signal_10428 ;
    wire new_AGEMA_signal_10429 ;
    wire new_AGEMA_signal_10430 ;
    wire new_AGEMA_signal_10431 ;
    wire new_AGEMA_signal_10432 ;
    wire new_AGEMA_signal_10433 ;
    wire new_AGEMA_signal_10434 ;
    wire new_AGEMA_signal_10435 ;
    wire new_AGEMA_signal_10436 ;
    wire new_AGEMA_signal_10437 ;
    wire new_AGEMA_signal_10438 ;
    wire new_AGEMA_signal_10439 ;
    wire new_AGEMA_signal_10440 ;
    wire new_AGEMA_signal_10441 ;
    wire new_AGEMA_signal_10442 ;
    wire new_AGEMA_signal_10443 ;
    wire new_AGEMA_signal_10444 ;
    wire new_AGEMA_signal_10445 ;
    wire new_AGEMA_signal_10446 ;
    wire new_AGEMA_signal_10447 ;
    wire new_AGEMA_signal_10448 ;
    wire new_AGEMA_signal_10449 ;
    wire new_AGEMA_signal_10450 ;
    wire new_AGEMA_signal_10451 ;
    wire new_AGEMA_signal_10452 ;
    wire new_AGEMA_signal_10453 ;
    wire new_AGEMA_signal_10454 ;
    wire new_AGEMA_signal_10455 ;
    wire new_AGEMA_signal_10456 ;
    wire new_AGEMA_signal_10457 ;
    wire new_AGEMA_signal_10458 ;
    wire new_AGEMA_signal_10459 ;
    wire new_AGEMA_signal_10460 ;
    wire new_AGEMA_signal_10461 ;
    wire new_AGEMA_signal_10462 ;
    wire new_AGEMA_signal_10463 ;
    wire new_AGEMA_signal_10464 ;
    wire new_AGEMA_signal_10465 ;
    wire new_AGEMA_signal_10466 ;
    wire new_AGEMA_signal_10467 ;

    /* cells in depth 0 */
    not_masked #(.security_order(2), .pipeline(1)) U1938 ( .a ({SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({new_AGEMA_signal_945, new_AGEMA_signal_944, n2796}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1939 ( .a ({SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({new_AGEMA_signal_949, new_AGEMA_signal_948, n2810}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1940 ( .a ({SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_953, new_AGEMA_signal_952, n2462}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1941 ( .a ({SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_957, new_AGEMA_signal_956, n2760}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1942 ( .a ({SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_961, new_AGEMA_signal_960, n2791}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1944 ( .a ({SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({new_AGEMA_signal_965, new_AGEMA_signal_964, n2813}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1945 ( .a ({SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_969, new_AGEMA_signal_968, n2630}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1946 ( .a ({SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_973, new_AGEMA_signal_972, n2765}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_927 ( .C ( clk ), .D ( SI_s0[4] ), .Q ( new_AGEMA_signal_5416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_929 ( .C ( clk ), .D ( SI_s1[4] ), .Q ( new_AGEMA_signal_5418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_931 ( .C ( clk ), .D ( SI_s2[4] ), .Q ( new_AGEMA_signal_5420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_933 ( .C ( clk ), .D ( SI_s0[6] ), .Q ( new_AGEMA_signal_5422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_935 ( .C ( clk ), .D ( SI_s1[6] ), .Q ( new_AGEMA_signal_5424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_937 ( .C ( clk ), .D ( SI_s2[6] ), .Q ( new_AGEMA_signal_5426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_939 ( .C ( clk ), .D ( SI_s0[7] ), .Q ( new_AGEMA_signal_5428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_941 ( .C ( clk ), .D ( SI_s1[7] ), .Q ( new_AGEMA_signal_5430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_943 ( .C ( clk ), .D ( SI_s2[7] ), .Q ( new_AGEMA_signal_5432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_945 ( .C ( clk ), .D ( SI_s0[0] ), .Q ( new_AGEMA_signal_5434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_947 ( .C ( clk ), .D ( SI_s1[0] ), .Q ( new_AGEMA_signal_5436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_949 ( .C ( clk ), .D ( SI_s2[0] ), .Q ( new_AGEMA_signal_5438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_951 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( new_AGEMA_signal_5440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_953 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( new_AGEMA_signal_5442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_955 ( .C ( clk ), .D ( SI_s2[1] ), .Q ( new_AGEMA_signal_5444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_957 ( .C ( clk ), .D ( n2630 ), .Q ( new_AGEMA_signal_5446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_959 ( .C ( clk ), .D ( new_AGEMA_signal_968 ), .Q ( new_AGEMA_signal_5448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_961 ( .C ( clk ), .D ( new_AGEMA_signal_969 ), .Q ( new_AGEMA_signal_5450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_963 ( .C ( clk ), .D ( SI_s0[5] ), .Q ( new_AGEMA_signal_5452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_965 ( .C ( clk ), .D ( SI_s1[5] ), .Q ( new_AGEMA_signal_5454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_967 ( .C ( clk ), .D ( SI_s2[5] ), .Q ( new_AGEMA_signal_5456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_969 ( .C ( clk ), .D ( n2462 ), .Q ( new_AGEMA_signal_5458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_971 ( .C ( clk ), .D ( new_AGEMA_signal_952 ), .Q ( new_AGEMA_signal_5460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_973 ( .C ( clk ), .D ( new_AGEMA_signal_953 ), .Q ( new_AGEMA_signal_5462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_975 ( .C ( clk ), .D ( n2760 ), .Q ( new_AGEMA_signal_5464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_977 ( .C ( clk ), .D ( new_AGEMA_signal_956 ), .Q ( new_AGEMA_signal_5466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_979 ( .C ( clk ), .D ( new_AGEMA_signal_957 ), .Q ( new_AGEMA_signal_5468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_981 ( .C ( clk ), .D ( n2796 ), .Q ( new_AGEMA_signal_5470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_983 ( .C ( clk ), .D ( new_AGEMA_signal_944 ), .Q ( new_AGEMA_signal_5472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_985 ( .C ( clk ), .D ( new_AGEMA_signal_945 ), .Q ( new_AGEMA_signal_5474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_987 ( .C ( clk ), .D ( n2765 ), .Q ( new_AGEMA_signal_5476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_989 ( .C ( clk ), .D ( new_AGEMA_signal_972 ), .Q ( new_AGEMA_signal_5478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_991 ( .C ( clk ), .D ( new_AGEMA_signal_973 ), .Q ( new_AGEMA_signal_5480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_993 ( .C ( clk ), .D ( n2791 ), .Q ( new_AGEMA_signal_5482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_995 ( .C ( clk ), .D ( new_AGEMA_signal_960 ), .Q ( new_AGEMA_signal_5484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_997 ( .C ( clk ), .D ( new_AGEMA_signal_961 ), .Q ( new_AGEMA_signal_5486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_999 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( new_AGEMA_signal_5488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1001 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( new_AGEMA_signal_5490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1003 ( .C ( clk ), .D ( SI_s2[3] ), .Q ( new_AGEMA_signal_5492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1005 ( .C ( clk ), .D ( n2813 ), .Q ( new_AGEMA_signal_5494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1007 ( .C ( clk ), .D ( new_AGEMA_signal_964 ), .Q ( new_AGEMA_signal_5496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1009 ( .C ( clk ), .D ( new_AGEMA_signal_965 ), .Q ( new_AGEMA_signal_5498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1011 ( .C ( clk ), .D ( n2810 ), .Q ( new_AGEMA_signal_5500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1013 ( .C ( clk ), .D ( new_AGEMA_signal_948 ), .Q ( new_AGEMA_signal_5502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1015 ( .C ( clk ), .D ( new_AGEMA_signal_949 ), .Q ( new_AGEMA_signal_5504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( new_AGEMA_signal_6274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( new_AGEMA_signal_6280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C ( clk ), .D ( SI_s2[2] ), .Q ( new_AGEMA_signal_6286 ) ) ;

    /* cells in depth 2 */
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1937 ( .a ({new_AGEMA_signal_945, new_AGEMA_signal_944, n2796}), .b ({SI_s2[6], SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_999, new_AGEMA_signal_998, n2719}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1943 ( .a ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, n2624}), .b ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2672}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1947 ( .a ({SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({new_AGEMA_signal_975, new_AGEMA_signal_974, n2635}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1948 ( .a ({new_AGEMA_signal_953, new_AGEMA_signal_952, n2462}), .b ({SI_s2[7], SI_s1[7], SI_s0[7]}), .clk ( clk ), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, n2641}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1949 ( .a ({SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({new_AGEMA_signal_977, new_AGEMA_signal_976, n2790}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1950 ( .a ({SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({SI_s2[7], SI_s1[7], SI_s0[7]}), .clk ( clk ), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_979, new_AGEMA_signal_978, n2519}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1951 ( .a ({new_AGEMA_signal_979, new_AGEMA_signal_978, n2519}), .b ({new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2750}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1952 ( .a ({new_AGEMA_signal_957, new_AGEMA_signal_956, n2760}), .b ({SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, n2615}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1953 ( .a ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, n2615}), .b ({new_AGEMA_signal_1107, new_AGEMA_signal_1106, n2640}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1955 ( .a ({new_AGEMA_signal_973, new_AGEMA_signal_972, n2765}), .b ({new_AGEMA_signal_969, new_AGEMA_signal_968, n2630}), .clk ( clk ), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, n2699}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1956 ( .a ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, n2699}), .b ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, n2737}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1957 ( .a ({new_AGEMA_signal_973, new_AGEMA_signal_972, n2765}), .b ({new_AGEMA_signal_965, new_AGEMA_signal_964, n2813}), .clk ( clk ), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2816}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1958 ( .a ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2816}), .b ({new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2767}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1961 ( .a ({new_AGEMA_signal_973, new_AGEMA_signal_972, n2765}), .b ({SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_1011, new_AGEMA_signal_1010, n2780}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1962 ( .a ({new_AGEMA_signal_1011, new_AGEMA_signal_1010, n2780}), .b ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, n2789}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1963 ( .a ({SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_949, new_AGEMA_signal_948, n2810}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, n2317}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1965 ( .a ({new_AGEMA_signal_961, new_AGEMA_signal_960, n2791}), .b ({new_AGEMA_signal_957, new_AGEMA_signal_956, n2760}), .clk ( clk ), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2694}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1966 ( .a ({new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2694}), .b ({new_AGEMA_signal_1115, new_AGEMA_signal_1114, n2769}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1969 ( .a ({new_AGEMA_signal_957, new_AGEMA_signal_956, n2760}), .b ({SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, n2073}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1970 ( .a ({new_AGEMA_signal_1017, new_AGEMA_signal_1016, n2073}), .b ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2707}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1971 ( .a ({SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_981, new_AGEMA_signal_980, n2315}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1972 ( .a ({SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({new_AGEMA_signal_983, new_AGEMA_signal_982, n2682}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1973 ( .a ({new_AGEMA_signal_983, new_AGEMA_signal_982, n2682}), .b ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2713}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1975 ( .a ({new_AGEMA_signal_965, new_AGEMA_signal_964, n2813}), .b ({SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2723}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1976 ( .a ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2723}), .b ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, n2688}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1978 ( .a ({new_AGEMA_signal_949, new_AGEMA_signal_948, n2810}), .b ({SI_s2[7], SI_s1[7], SI_s0[7]}), .clk ( clk ), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({new_AGEMA_signal_1023, new_AGEMA_signal_1022, n2725}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1979 ( .a ({new_AGEMA_signal_1023, new_AGEMA_signal_1022, n2725}), .b ({new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2541}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1984 ( .a ({new_AGEMA_signal_957, new_AGEMA_signal_956, n2760}), .b ({SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, n2815}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1985 ( .a ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, n2815}), .b ({new_AGEMA_signal_1125, new_AGEMA_signal_1124, n2086}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1987 ( .a ({new_AGEMA_signal_949, new_AGEMA_signal_948, n2810}), .b ({new_AGEMA_signal_961, new_AGEMA_signal_960, n2791}), .clk ( clk ), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2600}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1990 ( .a ({new_AGEMA_signal_953, new_AGEMA_signal_952, n2462}), .b ({SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_1029, new_AGEMA_signal_1028, n2538}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1991 ( .a ({new_AGEMA_signal_1029, new_AGEMA_signal_1028, n2538}), .b ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2786}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1995 ( .a ({SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({new_AGEMA_signal_985, new_AGEMA_signal_984, n2595}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1996 ( .a ({new_AGEMA_signal_985, new_AGEMA_signal_984, n2595}), .b ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, n2742}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1999 ( .a ({new_AGEMA_signal_973, new_AGEMA_signal_972, n2765}), .b ({new_AGEMA_signal_969, new_AGEMA_signal_968, n2630}), .clk ( clk ), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2753}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2000 ( .a ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2753}), .b ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, n2577}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2004 ( .a ({new_AGEMA_signal_949, new_AGEMA_signal_948, n2810}), .b ({SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({new_AGEMA_signal_1035, new_AGEMA_signal_1034, n2400}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2008 ( .a ({new_AGEMA_signal_973, new_AGEMA_signal_972, n2765}), .b ({SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, n2785}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2009 ( .a ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, n2785}), .b ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, n2792}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2013 ( .a ({new_AGEMA_signal_965, new_AGEMA_signal_964, n2813}), .b ({SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2609}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2014 ( .a ({new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2609}), .b ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, n2724}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2017 ( .a ({new_AGEMA_signal_957, new_AGEMA_signal_956, n2760}), .b ({new_AGEMA_signal_965, new_AGEMA_signal_964, n2813}), .clk ( clk ), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_1041, new_AGEMA_signal_1040, n2661}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2018 ( .a ({new_AGEMA_signal_1041, new_AGEMA_signal_1040, n2661}), .b ({new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2174}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2020 ( .a ({SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({new_AGEMA_signal_987, new_AGEMA_signal_986, n2708}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2021 ( .a ({new_AGEMA_signal_987, new_AGEMA_signal_986, n2708}), .b ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, n2493}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2025 ( .a ({new_AGEMA_signal_945, new_AGEMA_signal_944, n2796}), .b ({SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2587}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2028 ( .a ({new_AGEMA_signal_999, new_AGEMA_signal_998, n2719}), .b ({new_AGEMA_signal_1147, new_AGEMA_signal_1146, n2570}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2029 ( .a ({SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({new_AGEMA_signal_989, new_AGEMA_signal_988, n2559}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2035 ( .a ({new_AGEMA_signal_973, new_AGEMA_signal_972, n2765}), .b ({SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_1047, new_AGEMA_signal_1046, n2643}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2036 ( .a ({new_AGEMA_signal_1047, new_AGEMA_signal_1046, n2643}), .b ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, n2442}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2038 ( .a ({new_AGEMA_signal_977, new_AGEMA_signal_976, n2790}), .b ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, n2739}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2044 ( .a ({new_AGEMA_signal_953, new_AGEMA_signal_952, n2462}), .b ({new_AGEMA_signal_945, new_AGEMA_signal_944, n2796}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2437}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2045 ( .a ({SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_991, new_AGEMA_signal_990, n2261}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2046 ( .a ({new_AGEMA_signal_991, new_AGEMA_signal_990, n2261}), .b ({new_AGEMA_signal_1053, new_AGEMA_signal_1052, n2778}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2052 ( .a ({SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({new_AGEMA_signal_961, new_AGEMA_signal_960, n2791}), .clk ( clk ), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({new_AGEMA_signal_1055, new_AGEMA_signal_1054, n2452}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2055 ( .a ({new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2437}), .b ({new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2766}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2068 ( .a ({new_AGEMA_signal_973, new_AGEMA_signal_972, n2765}), .b ({SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_1059, new_AGEMA_signal_1058, n2772}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2070 ( .a ({new_AGEMA_signal_961, new_AGEMA_signal_960, n2791}), .b ({SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, n2824}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2071 ( .a ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, n2824}), .b ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, n2612}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2074 ( .a ({new_AGEMA_signal_1035, new_AGEMA_signal_1034, n2400}), .b ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, n2313}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2089 ( .a ({new_AGEMA_signal_949, new_AGEMA_signal_948, n2810}), .b ({new_AGEMA_signal_957, new_AGEMA_signal_956, n2760}), .clk ( clk ), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2395}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2090 ( .a ({new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2395}), .b ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, n2818}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2094 ( .a ({SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({new_AGEMA_signal_993, new_AGEMA_signal_992, n2779}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2096 ( .a ({new_AGEMA_signal_969, new_AGEMA_signal_968, n2630}), .b ({new_AGEMA_signal_965, new_AGEMA_signal_964, n2813}), .clk ( clk ), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, n2624}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2097 ( .a ({SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({new_AGEMA_signal_995, new_AGEMA_signal_994, n2242}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2100 ( .a ({SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_961, new_AGEMA_signal_960, n2791}), .clk ( clk ), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, n2356}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2119 ( .a ({new_AGEMA_signal_1059, new_AGEMA_signal_1058, n2772}), .b ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, n2823}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2122 ( .a ({new_AGEMA_signal_957, new_AGEMA_signal_956, n2760}), .b ({SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2611}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2131 ( .a ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, n2641}), .b ({new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2828}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2133 ( .a ({new_AGEMA_signal_973, new_AGEMA_signal_972, n2765}), .b ({SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_1071, new_AGEMA_signal_1070, n2616}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2134 ( .a ({new_AGEMA_signal_1071, new_AGEMA_signal_1070, n2616}), .b ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, n2679}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2138 ( .a ({new_AGEMA_signal_973, new_AGEMA_signal_972, n2765}), .b ({new_AGEMA_signal_957, new_AGEMA_signal_956, n2760}), .clk ( clk ), .r ({Fresh[125], Fresh[124], Fresh[123]}), .c ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, n2563}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2139 ( .a ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, n2563}), .b ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, n2809}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2150 ( .a ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2611}), .b ({new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2709}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2163 ( .a ({new_AGEMA_signal_945, new_AGEMA_signal_944, n2796}), .b ({new_AGEMA_signal_949, new_AGEMA_signal_948, n2810}), .clk ( clk ), .r ({Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2401}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2211 ( .a ({new_AGEMA_signal_973, new_AGEMA_signal_972, n2765}), .b ({SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[131], Fresh[130], Fresh[129]}), .c ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, n2061}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2232 ( .a ({new_AGEMA_signal_945, new_AGEMA_signal_944, n2796}), .b ({new_AGEMA_signal_961, new_AGEMA_signal_960, n2791}), .clk ( clk ), .r ({Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2721}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2276 ( .a ({new_AGEMA_signal_961, new_AGEMA_signal_960, n2791}), .b ({new_AGEMA_signal_973, new_AGEMA_signal_972, n2765}), .clk ( clk ), .r ({Fresh[137], Fresh[136], Fresh[135]}), .c ({new_AGEMA_signal_1083, new_AGEMA_signal_1082, n2298}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2278 ( .a ({new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2401}), .b ({new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2118}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2307 ( .a ({SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_969, new_AGEMA_signal_968, n2630}), .clk ( clk ), .r ({Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, n2346}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2341 ( .a ({SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_961, new_AGEMA_signal_960, n2791}), .clk ( clk ), .r ({Fresh[143], Fresh[142], Fresh[141]}), .c ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, n2430}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2383 ( .a ({SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_997, new_AGEMA_signal_996, n2712}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2402 ( .a ({SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_965, new_AGEMA_signal_964, n2813}), .clk ( clk ), .r ({Fresh[149], Fresh[148], Fresh[147]}), .c ({new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2777}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2615 ( .a ({SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_953, new_AGEMA_signal_952, n2462}), .clk ( clk ), .r ({Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, n2463}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2627 ( .a ({new_AGEMA_signal_949, new_AGEMA_signal_948, n2810}), .b ({SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[155], Fresh[154], Fresh[153]}), .c ({new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2474}) ) ;
    buf_clk new_AGEMA_reg_buffer_928 ( .C ( clk ), .D ( new_AGEMA_signal_5416 ), .Q ( new_AGEMA_signal_5417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_930 ( .C ( clk ), .D ( new_AGEMA_signal_5418 ), .Q ( new_AGEMA_signal_5419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_932 ( .C ( clk ), .D ( new_AGEMA_signal_5420 ), .Q ( new_AGEMA_signal_5421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_934 ( .C ( clk ), .D ( new_AGEMA_signal_5422 ), .Q ( new_AGEMA_signal_5423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_936 ( .C ( clk ), .D ( new_AGEMA_signal_5424 ), .Q ( new_AGEMA_signal_5425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_938 ( .C ( clk ), .D ( new_AGEMA_signal_5426 ), .Q ( new_AGEMA_signal_5427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_940 ( .C ( clk ), .D ( new_AGEMA_signal_5428 ), .Q ( new_AGEMA_signal_5429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_942 ( .C ( clk ), .D ( new_AGEMA_signal_5430 ), .Q ( new_AGEMA_signal_5431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_944 ( .C ( clk ), .D ( new_AGEMA_signal_5432 ), .Q ( new_AGEMA_signal_5433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_946 ( .C ( clk ), .D ( new_AGEMA_signal_5434 ), .Q ( new_AGEMA_signal_5435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_948 ( .C ( clk ), .D ( new_AGEMA_signal_5436 ), .Q ( new_AGEMA_signal_5437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_950 ( .C ( clk ), .D ( new_AGEMA_signal_5438 ), .Q ( new_AGEMA_signal_5439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_952 ( .C ( clk ), .D ( new_AGEMA_signal_5440 ), .Q ( new_AGEMA_signal_5441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_954 ( .C ( clk ), .D ( new_AGEMA_signal_5442 ), .Q ( new_AGEMA_signal_5443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_956 ( .C ( clk ), .D ( new_AGEMA_signal_5444 ), .Q ( new_AGEMA_signal_5445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_958 ( .C ( clk ), .D ( new_AGEMA_signal_5446 ), .Q ( new_AGEMA_signal_5447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_960 ( .C ( clk ), .D ( new_AGEMA_signal_5448 ), .Q ( new_AGEMA_signal_5449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_962 ( .C ( clk ), .D ( new_AGEMA_signal_5450 ), .Q ( new_AGEMA_signal_5451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_964 ( .C ( clk ), .D ( new_AGEMA_signal_5452 ), .Q ( new_AGEMA_signal_5453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_966 ( .C ( clk ), .D ( new_AGEMA_signal_5454 ), .Q ( new_AGEMA_signal_5455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_968 ( .C ( clk ), .D ( new_AGEMA_signal_5456 ), .Q ( new_AGEMA_signal_5457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_970 ( .C ( clk ), .D ( new_AGEMA_signal_5458 ), .Q ( new_AGEMA_signal_5459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_972 ( .C ( clk ), .D ( new_AGEMA_signal_5460 ), .Q ( new_AGEMA_signal_5461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_974 ( .C ( clk ), .D ( new_AGEMA_signal_5462 ), .Q ( new_AGEMA_signal_5463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_976 ( .C ( clk ), .D ( new_AGEMA_signal_5464 ), .Q ( new_AGEMA_signal_5465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_978 ( .C ( clk ), .D ( new_AGEMA_signal_5466 ), .Q ( new_AGEMA_signal_5467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_980 ( .C ( clk ), .D ( new_AGEMA_signal_5468 ), .Q ( new_AGEMA_signal_5469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_982 ( .C ( clk ), .D ( new_AGEMA_signal_5470 ), .Q ( new_AGEMA_signal_5471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_984 ( .C ( clk ), .D ( new_AGEMA_signal_5472 ), .Q ( new_AGEMA_signal_5473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_986 ( .C ( clk ), .D ( new_AGEMA_signal_5474 ), .Q ( new_AGEMA_signal_5475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_988 ( .C ( clk ), .D ( new_AGEMA_signal_5476 ), .Q ( new_AGEMA_signal_5477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_990 ( .C ( clk ), .D ( new_AGEMA_signal_5478 ), .Q ( new_AGEMA_signal_5479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_992 ( .C ( clk ), .D ( new_AGEMA_signal_5480 ), .Q ( new_AGEMA_signal_5481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_994 ( .C ( clk ), .D ( new_AGEMA_signal_5482 ), .Q ( new_AGEMA_signal_5483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_996 ( .C ( clk ), .D ( new_AGEMA_signal_5484 ), .Q ( new_AGEMA_signal_5485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_998 ( .C ( clk ), .D ( new_AGEMA_signal_5486 ), .Q ( new_AGEMA_signal_5487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1000 ( .C ( clk ), .D ( new_AGEMA_signal_5488 ), .Q ( new_AGEMA_signal_5489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1002 ( .C ( clk ), .D ( new_AGEMA_signal_5490 ), .Q ( new_AGEMA_signal_5491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1004 ( .C ( clk ), .D ( new_AGEMA_signal_5492 ), .Q ( new_AGEMA_signal_5493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1006 ( .C ( clk ), .D ( new_AGEMA_signal_5494 ), .Q ( new_AGEMA_signal_5495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1008 ( .C ( clk ), .D ( new_AGEMA_signal_5496 ), .Q ( new_AGEMA_signal_5497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1010 ( .C ( clk ), .D ( new_AGEMA_signal_5498 ), .Q ( new_AGEMA_signal_5499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1012 ( .C ( clk ), .D ( new_AGEMA_signal_5500 ), .Q ( new_AGEMA_signal_5501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1014 ( .C ( clk ), .D ( new_AGEMA_signal_5502 ), .Q ( new_AGEMA_signal_5503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1016 ( .C ( clk ), .D ( new_AGEMA_signal_5504 ), .Q ( new_AGEMA_signal_5505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C ( clk ), .D ( new_AGEMA_signal_6274 ), .Q ( new_AGEMA_signal_6275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C ( clk ), .D ( new_AGEMA_signal_6280 ), .Q ( new_AGEMA_signal_6281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C ( clk ), .D ( new_AGEMA_signal_6286 ), .Q ( new_AGEMA_signal_6287 ) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_1017 ( .C ( clk ), .D ( n2769 ), .Q ( new_AGEMA_signal_5506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1019 ( .C ( clk ), .D ( new_AGEMA_signal_1114 ), .Q ( new_AGEMA_signal_5508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1021 ( .C ( clk ), .D ( new_AGEMA_signal_1115 ), .Q ( new_AGEMA_signal_5510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1023 ( .C ( clk ), .D ( new_AGEMA_signal_5489 ), .Q ( new_AGEMA_signal_5512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1025 ( .C ( clk ), .D ( new_AGEMA_signal_5491 ), .Q ( new_AGEMA_signal_5514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1027 ( .C ( clk ), .D ( new_AGEMA_signal_5493 ), .Q ( new_AGEMA_signal_5516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1029 ( .C ( clk ), .D ( new_AGEMA_signal_5423 ), .Q ( new_AGEMA_signal_5518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1031 ( .C ( clk ), .D ( new_AGEMA_signal_5425 ), .Q ( new_AGEMA_signal_5520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1033 ( .C ( clk ), .D ( new_AGEMA_signal_5427 ), .Q ( new_AGEMA_signal_5522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1035 ( .C ( clk ), .D ( n2174 ), .Q ( new_AGEMA_signal_5524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1037 ( .C ( clk ), .D ( new_AGEMA_signal_1140 ), .Q ( new_AGEMA_signal_5526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1039 ( .C ( clk ), .D ( new_AGEMA_signal_1141 ), .Q ( new_AGEMA_signal_5528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1041 ( .C ( clk ), .D ( new_AGEMA_signal_5417 ), .Q ( new_AGEMA_signal_5530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1043 ( .C ( clk ), .D ( new_AGEMA_signal_5419 ), .Q ( new_AGEMA_signal_5532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1045 ( .C ( clk ), .D ( new_AGEMA_signal_5421 ), .Q ( new_AGEMA_signal_5534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1047 ( .C ( clk ), .D ( new_AGEMA_signal_5435 ), .Q ( new_AGEMA_signal_5536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1049 ( .C ( clk ), .D ( new_AGEMA_signal_5437 ), .Q ( new_AGEMA_signal_5538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1051 ( .C ( clk ), .D ( new_AGEMA_signal_5439 ), .Q ( new_AGEMA_signal_5540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1053 ( .C ( clk ), .D ( n2570 ), .Q ( new_AGEMA_signal_5542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1055 ( .C ( clk ), .D ( new_AGEMA_signal_1146 ), .Q ( new_AGEMA_signal_5544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1057 ( .C ( clk ), .D ( new_AGEMA_signal_1147 ), .Q ( new_AGEMA_signal_5546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1059 ( .C ( clk ), .D ( n2792 ), .Q ( new_AGEMA_signal_5548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1061 ( .C ( clk ), .D ( new_AGEMA_signal_1136 ), .Q ( new_AGEMA_signal_5550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1063 ( .C ( clk ), .D ( new_AGEMA_signal_1137 ), .Q ( new_AGEMA_signal_5552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1065 ( .C ( clk ), .D ( n2635 ), .Q ( new_AGEMA_signal_5554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1067 ( .C ( clk ), .D ( new_AGEMA_signal_974 ), .Q ( new_AGEMA_signal_5556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1069 ( .C ( clk ), .D ( new_AGEMA_signal_975 ), .Q ( new_AGEMA_signal_5558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1071 ( .C ( clk ), .D ( n2587 ), .Q ( new_AGEMA_signal_5560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1073 ( .C ( clk ), .D ( new_AGEMA_signal_1044 ), .Q ( new_AGEMA_signal_5562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1075 ( .C ( clk ), .D ( new_AGEMA_signal_1045 ), .Q ( new_AGEMA_signal_5564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1077 ( .C ( clk ), .D ( n2725 ), .Q ( new_AGEMA_signal_5566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1079 ( .C ( clk ), .D ( new_AGEMA_signal_1022 ), .Q ( new_AGEMA_signal_5568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1081 ( .C ( clk ), .D ( new_AGEMA_signal_1023 ), .Q ( new_AGEMA_signal_5570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1083 ( .C ( clk ), .D ( n2708 ), .Q ( new_AGEMA_signal_5572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1085 ( .C ( clk ), .D ( new_AGEMA_signal_986 ), .Q ( new_AGEMA_signal_5574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1087 ( .C ( clk ), .D ( new_AGEMA_signal_987 ), .Q ( new_AGEMA_signal_5576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1089 ( .C ( clk ), .D ( n2818 ), .Q ( new_AGEMA_signal_5578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1091 ( .C ( clk ), .D ( new_AGEMA_signal_1174 ), .Q ( new_AGEMA_signal_5580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1093 ( .C ( clk ), .D ( new_AGEMA_signal_1175 ), .Q ( new_AGEMA_signal_5582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1095 ( .C ( clk ), .D ( n2790 ), .Q ( new_AGEMA_signal_5584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1097 ( .C ( clk ), .D ( new_AGEMA_signal_976 ), .Q ( new_AGEMA_signal_5586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1099 ( .C ( clk ), .D ( new_AGEMA_signal_977 ), .Q ( new_AGEMA_signal_5588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1101 ( .C ( clk ), .D ( n2786 ), .Q ( new_AGEMA_signal_5590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1103 ( .C ( clk ), .D ( new_AGEMA_signal_1128 ), .Q ( new_AGEMA_signal_5592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1105 ( .C ( clk ), .D ( new_AGEMA_signal_1129 ), .Q ( new_AGEMA_signal_5594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1107 ( .C ( clk ), .D ( n2400 ), .Q ( new_AGEMA_signal_5596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1109 ( .C ( clk ), .D ( new_AGEMA_signal_1034 ), .Q ( new_AGEMA_signal_5598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1111 ( .C ( clk ), .D ( new_AGEMA_signal_1035 ), .Q ( new_AGEMA_signal_5600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1113 ( .C ( clk ), .D ( new_AGEMA_signal_5441 ), .Q ( new_AGEMA_signal_5602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1115 ( .C ( clk ), .D ( new_AGEMA_signal_5443 ), .Q ( new_AGEMA_signal_5604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1117 ( .C ( clk ), .D ( new_AGEMA_signal_5445 ), .Q ( new_AGEMA_signal_5606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1119 ( .C ( clk ), .D ( n2815 ), .Q ( new_AGEMA_signal_5608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1121 ( .C ( clk ), .D ( new_AGEMA_signal_1024 ), .Q ( new_AGEMA_signal_5610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1123 ( .C ( clk ), .D ( new_AGEMA_signal_1025 ), .Q ( new_AGEMA_signal_5612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1125 ( .C ( clk ), .D ( n2723 ), .Q ( new_AGEMA_signal_5614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1127 ( .C ( clk ), .D ( new_AGEMA_signal_1020 ), .Q ( new_AGEMA_signal_5616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1129 ( .C ( clk ), .D ( new_AGEMA_signal_1021 ), .Q ( new_AGEMA_signal_5618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1131 ( .C ( clk ), .D ( n2709 ), .Q ( new_AGEMA_signal_5620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1133 ( .C ( clk ), .D ( new_AGEMA_signal_1194 ), .Q ( new_AGEMA_signal_5622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1135 ( .C ( clk ), .D ( new_AGEMA_signal_1195 ), .Q ( new_AGEMA_signal_5624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1137 ( .C ( clk ), .D ( n2753 ), .Q ( new_AGEMA_signal_5626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1139 ( .C ( clk ), .D ( new_AGEMA_signal_1032 ), .Q ( new_AGEMA_signal_5628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1141 ( .C ( clk ), .D ( new_AGEMA_signal_1033 ), .Q ( new_AGEMA_signal_5630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1143 ( .C ( clk ), .D ( n2401 ), .Q ( new_AGEMA_signal_5632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1145 ( .C ( clk ), .D ( new_AGEMA_signal_1074 ), .Q ( new_AGEMA_signal_5634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1147 ( .C ( clk ), .D ( new_AGEMA_signal_1075 ), .Q ( new_AGEMA_signal_5636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1149 ( .C ( clk ), .D ( new_AGEMA_signal_5477 ), .Q ( new_AGEMA_signal_5638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1151 ( .C ( clk ), .D ( new_AGEMA_signal_5479 ), .Q ( new_AGEMA_signal_5640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1153 ( .C ( clk ), .D ( new_AGEMA_signal_5481 ), .Q ( new_AGEMA_signal_5642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1155 ( .C ( clk ), .D ( new_AGEMA_signal_5447 ), .Q ( new_AGEMA_signal_5644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1157 ( .C ( clk ), .D ( new_AGEMA_signal_5449 ), .Q ( new_AGEMA_signal_5646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1159 ( .C ( clk ), .D ( new_AGEMA_signal_5451 ), .Q ( new_AGEMA_signal_5648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1161 ( .C ( clk ), .D ( n2615 ), .Q ( new_AGEMA_signal_5650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1163 ( .C ( clk ), .D ( new_AGEMA_signal_1004 ), .Q ( new_AGEMA_signal_5652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1165 ( .C ( clk ), .D ( new_AGEMA_signal_1005 ), .Q ( new_AGEMA_signal_5654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1167 ( .C ( clk ), .D ( n2643 ), .Q ( new_AGEMA_signal_5656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1169 ( .C ( clk ), .D ( new_AGEMA_signal_1046 ), .Q ( new_AGEMA_signal_5658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1171 ( .C ( clk ), .D ( new_AGEMA_signal_1047 ), .Q ( new_AGEMA_signal_5660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1173 ( .C ( clk ), .D ( n2563 ), .Q ( new_AGEMA_signal_5662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1175 ( .C ( clk ), .D ( new_AGEMA_signal_1072 ), .Q ( new_AGEMA_signal_5664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1177 ( .C ( clk ), .D ( new_AGEMA_signal_1073 ), .Q ( new_AGEMA_signal_5666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1179 ( .C ( clk ), .D ( n2612 ), .Q ( new_AGEMA_signal_5668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1181 ( .C ( clk ), .D ( new_AGEMA_signal_1164 ), .Q ( new_AGEMA_signal_5670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1183 ( .C ( clk ), .D ( new_AGEMA_signal_1165 ), .Q ( new_AGEMA_signal_5672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1185 ( .C ( clk ), .D ( n2824 ), .Q ( new_AGEMA_signal_5674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1187 ( .C ( clk ), .D ( new_AGEMA_signal_1060 ), .Q ( new_AGEMA_signal_5676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1189 ( .C ( clk ), .D ( new_AGEMA_signal_1061 ), .Q ( new_AGEMA_signal_5678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1191 ( .C ( clk ), .D ( n2816 ), .Q ( new_AGEMA_signal_5680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1193 ( .C ( clk ), .D ( new_AGEMA_signal_1008 ), .Q ( new_AGEMA_signal_5682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1195 ( .C ( clk ), .D ( new_AGEMA_signal_1009 ), .Q ( new_AGEMA_signal_5684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1197 ( .C ( clk ), .D ( n2073 ), .Q ( new_AGEMA_signal_5686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1199 ( .C ( clk ), .D ( new_AGEMA_signal_1016 ), .Q ( new_AGEMA_signal_5688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1201 ( .C ( clk ), .D ( new_AGEMA_signal_1017 ), .Q ( new_AGEMA_signal_5690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1203 ( .C ( clk ), .D ( n2519 ), .Q ( new_AGEMA_signal_5692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1205 ( .C ( clk ), .D ( new_AGEMA_signal_978 ), .Q ( new_AGEMA_signal_5694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1207 ( .C ( clk ), .D ( new_AGEMA_signal_979 ), .Q ( new_AGEMA_signal_5696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1209 ( .C ( clk ), .D ( n2616 ), .Q ( new_AGEMA_signal_5698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1211 ( .C ( clk ), .D ( new_AGEMA_signal_1070 ), .Q ( new_AGEMA_signal_5700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1213 ( .C ( clk ), .D ( new_AGEMA_signal_1071 ), .Q ( new_AGEMA_signal_5702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1215 ( .C ( clk ), .D ( new_AGEMA_signal_5483 ), .Q ( new_AGEMA_signal_5704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1217 ( .C ( clk ), .D ( new_AGEMA_signal_5485 ), .Q ( new_AGEMA_signal_5706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1219 ( .C ( clk ), .D ( new_AGEMA_signal_5487 ), .Q ( new_AGEMA_signal_5708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1221 ( .C ( clk ), .D ( n2780 ), .Q ( new_AGEMA_signal_5710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1223 ( .C ( clk ), .D ( new_AGEMA_signal_1010 ), .Q ( new_AGEMA_signal_5712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1225 ( .C ( clk ), .D ( new_AGEMA_signal_1011 ), .Q ( new_AGEMA_signal_5714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1227 ( .C ( clk ), .D ( new_AGEMA_signal_5495 ), .Q ( new_AGEMA_signal_5716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1229 ( .C ( clk ), .D ( new_AGEMA_signal_5497 ), .Q ( new_AGEMA_signal_5718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1231 ( .C ( clk ), .D ( new_AGEMA_signal_5499 ), .Q ( new_AGEMA_signal_5720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1233 ( .C ( clk ), .D ( n2742 ), .Q ( new_AGEMA_signal_5722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1235 ( .C ( clk ), .D ( new_AGEMA_signal_1030 ), .Q ( new_AGEMA_signal_5724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1237 ( .C ( clk ), .D ( new_AGEMA_signal_1031 ), .Q ( new_AGEMA_signal_5726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1239 ( .C ( clk ), .D ( n2724 ), .Q ( new_AGEMA_signal_5728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1241 ( .C ( clk ), .D ( new_AGEMA_signal_1138 ), .Q ( new_AGEMA_signal_5730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1243 ( .C ( clk ), .D ( new_AGEMA_signal_1139 ), .Q ( new_AGEMA_signal_5732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1245 ( .C ( clk ), .D ( n2317 ), .Q ( new_AGEMA_signal_5734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1247 ( .C ( clk ), .D ( new_AGEMA_signal_1012 ), .Q ( new_AGEMA_signal_5736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1249 ( .C ( clk ), .D ( new_AGEMA_signal_1013 ), .Q ( new_AGEMA_signal_5738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1251 ( .C ( clk ), .D ( n2688 ), .Q ( new_AGEMA_signal_5740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1253 ( .C ( clk ), .D ( new_AGEMA_signal_1120 ), .Q ( new_AGEMA_signal_5742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1255 ( .C ( clk ), .D ( new_AGEMA_signal_1121 ), .Q ( new_AGEMA_signal_5744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C ( clk ), .D ( n2609 ), .Q ( new_AGEMA_signal_5746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1259 ( .C ( clk ), .D ( new_AGEMA_signal_1038 ), .Q ( new_AGEMA_signal_5748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C ( clk ), .D ( new_AGEMA_signal_1039 ), .Q ( new_AGEMA_signal_5750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C ( clk ), .D ( n2672 ), .Q ( new_AGEMA_signal_5752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C ( clk ), .D ( new_AGEMA_signal_1104 ), .Q ( new_AGEMA_signal_5754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C ( clk ), .D ( new_AGEMA_signal_1105 ), .Q ( new_AGEMA_signal_5756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C ( clk ), .D ( n2640 ), .Q ( new_AGEMA_signal_5758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C ( clk ), .D ( new_AGEMA_signal_1106 ), .Q ( new_AGEMA_signal_5760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C ( clk ), .D ( new_AGEMA_signal_1107 ), .Q ( new_AGEMA_signal_5762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C ( clk ), .D ( n2713 ), .Q ( new_AGEMA_signal_5764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C ( clk ), .D ( new_AGEMA_signal_1018 ), .Q ( new_AGEMA_signal_5766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C ( clk ), .D ( new_AGEMA_signal_1019 ), .Q ( new_AGEMA_signal_5768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C ( clk ), .D ( n2777 ), .Q ( new_AGEMA_signal_5770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C ( clk ), .D ( new_AGEMA_signal_1092 ), .Q ( new_AGEMA_signal_5772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C ( clk ), .D ( new_AGEMA_signal_1093 ), .Q ( new_AGEMA_signal_5774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C ( clk ), .D ( n2789 ), .Q ( new_AGEMA_signal_5776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C ( clk ), .D ( new_AGEMA_signal_1112 ), .Q ( new_AGEMA_signal_5778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C ( clk ), .D ( new_AGEMA_signal_1113 ), .Q ( new_AGEMA_signal_5780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C ( clk ), .D ( n2661 ), .Q ( new_AGEMA_signal_5782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C ( clk ), .D ( new_AGEMA_signal_1040 ), .Q ( new_AGEMA_signal_5784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C ( clk ), .D ( new_AGEMA_signal_1041 ), .Q ( new_AGEMA_signal_5786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C ( clk ), .D ( new_AGEMA_signal_5459 ), .Q ( new_AGEMA_signal_5788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C ( clk ), .D ( new_AGEMA_signal_5461 ), .Q ( new_AGEMA_signal_5790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C ( clk ), .D ( new_AGEMA_signal_5463 ), .Q ( new_AGEMA_signal_5792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C ( clk ), .D ( n2694 ), .Q ( new_AGEMA_signal_5794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C ( clk ), .D ( new_AGEMA_signal_1014 ), .Q ( new_AGEMA_signal_5796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C ( clk ), .D ( new_AGEMA_signal_1015 ), .Q ( new_AGEMA_signal_5798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C ( clk ), .D ( new_AGEMA_signal_5465 ), .Q ( new_AGEMA_signal_5800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C ( clk ), .D ( new_AGEMA_signal_5467 ), .Q ( new_AGEMA_signal_5802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C ( clk ), .D ( new_AGEMA_signal_5469 ), .Q ( new_AGEMA_signal_5804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C ( clk ), .D ( n2682 ), .Q ( new_AGEMA_signal_5806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1319 ( .C ( clk ), .D ( new_AGEMA_signal_982 ), .Q ( new_AGEMA_signal_5808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1321 ( .C ( clk ), .D ( new_AGEMA_signal_983 ), .Q ( new_AGEMA_signal_5810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1323 ( .C ( clk ), .D ( new_AGEMA_signal_5501 ), .Q ( new_AGEMA_signal_5812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C ( clk ), .D ( new_AGEMA_signal_5503 ), .Q ( new_AGEMA_signal_5814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C ( clk ), .D ( new_AGEMA_signal_5505 ), .Q ( new_AGEMA_signal_5816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C ( clk ), .D ( n2624 ), .Q ( new_AGEMA_signal_5818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C ( clk ), .D ( new_AGEMA_signal_1064 ), .Q ( new_AGEMA_signal_5820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C ( clk ), .D ( new_AGEMA_signal_1065 ), .Q ( new_AGEMA_signal_5822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C ( clk ), .D ( n2356 ), .Q ( new_AGEMA_signal_5824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C ( clk ), .D ( new_AGEMA_signal_1066 ), .Q ( new_AGEMA_signal_5826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C ( clk ), .D ( new_AGEMA_signal_1067 ), .Q ( new_AGEMA_signal_5828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C ( clk ), .D ( n2778 ), .Q ( new_AGEMA_signal_5830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C ( clk ), .D ( new_AGEMA_signal_1052 ), .Q ( new_AGEMA_signal_5832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C ( clk ), .D ( new_AGEMA_signal_1053 ), .Q ( new_AGEMA_signal_5834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C ( clk ), .D ( n2766 ), .Q ( new_AGEMA_signal_5836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C ( clk ), .D ( new_AGEMA_signal_1158 ), .Q ( new_AGEMA_signal_5838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C ( clk ), .D ( new_AGEMA_signal_1159 ), .Q ( new_AGEMA_signal_5840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C ( clk ), .D ( n2767 ), .Q ( new_AGEMA_signal_5842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C ( clk ), .D ( new_AGEMA_signal_1110 ), .Q ( new_AGEMA_signal_5844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C ( clk ), .D ( new_AGEMA_signal_1111 ), .Q ( new_AGEMA_signal_5846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C ( clk ), .D ( n2641 ), .Q ( new_AGEMA_signal_5848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1361 ( .C ( clk ), .D ( new_AGEMA_signal_1000 ), .Q ( new_AGEMA_signal_5850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1363 ( .C ( clk ), .D ( new_AGEMA_signal_1001 ), .Q ( new_AGEMA_signal_5852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1365 ( .C ( clk ), .D ( n2719 ), .Q ( new_AGEMA_signal_5854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1367 ( .C ( clk ), .D ( new_AGEMA_signal_998 ), .Q ( new_AGEMA_signal_5856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1369 ( .C ( clk ), .D ( new_AGEMA_signal_999 ), .Q ( new_AGEMA_signal_5858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1371 ( .C ( clk ), .D ( n2707 ), .Q ( new_AGEMA_signal_5860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1373 ( .C ( clk ), .D ( new_AGEMA_signal_1116 ), .Q ( new_AGEMA_signal_5862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1375 ( .C ( clk ), .D ( new_AGEMA_signal_1117 ), .Q ( new_AGEMA_signal_5864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1377 ( .C ( clk ), .D ( n2493 ), .Q ( new_AGEMA_signal_5866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1379 ( .C ( clk ), .D ( new_AGEMA_signal_1042 ), .Q ( new_AGEMA_signal_5868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1381 ( .C ( clk ), .D ( new_AGEMA_signal_1043 ), .Q ( new_AGEMA_signal_5870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1383 ( .C ( clk ), .D ( n2577 ), .Q ( new_AGEMA_signal_5872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1385 ( .C ( clk ), .D ( new_AGEMA_signal_1132 ), .Q ( new_AGEMA_signal_5874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1387 ( .C ( clk ), .D ( new_AGEMA_signal_1133 ), .Q ( new_AGEMA_signal_5876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1389 ( .C ( clk ), .D ( n2541 ), .Q ( new_AGEMA_signal_5878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1391 ( .C ( clk ), .D ( new_AGEMA_signal_1122 ), .Q ( new_AGEMA_signal_5880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1393 ( .C ( clk ), .D ( new_AGEMA_signal_1123 ), .Q ( new_AGEMA_signal_5882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1395 ( .C ( clk ), .D ( n2679 ), .Q ( new_AGEMA_signal_5884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1397 ( .C ( clk ), .D ( new_AGEMA_signal_1190 ), .Q ( new_AGEMA_signal_5886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1399 ( .C ( clk ), .D ( new_AGEMA_signal_1191 ), .Q ( new_AGEMA_signal_5888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1401 ( .C ( clk ), .D ( n2699 ), .Q ( new_AGEMA_signal_5890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1403 ( .C ( clk ), .D ( new_AGEMA_signal_1006 ), .Q ( new_AGEMA_signal_5892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1405 ( .C ( clk ), .D ( new_AGEMA_signal_1007 ), .Q ( new_AGEMA_signal_5894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1407 ( .C ( clk ), .D ( n2611 ), .Q ( new_AGEMA_signal_5896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1409 ( .C ( clk ), .D ( new_AGEMA_signal_1068 ), .Q ( new_AGEMA_signal_5898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1411 ( .C ( clk ), .D ( new_AGEMA_signal_1069 ), .Q ( new_AGEMA_signal_5900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1413 ( .C ( clk ), .D ( n2739 ), .Q ( new_AGEMA_signal_5902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1415 ( .C ( clk ), .D ( new_AGEMA_signal_1048 ), .Q ( new_AGEMA_signal_5904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1417 ( .C ( clk ), .D ( new_AGEMA_signal_1049 ), .Q ( new_AGEMA_signal_5906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1419 ( .C ( clk ), .D ( n2772 ), .Q ( new_AGEMA_signal_5908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1421 ( .C ( clk ), .D ( new_AGEMA_signal_1058 ), .Q ( new_AGEMA_signal_5910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1423 ( .C ( clk ), .D ( new_AGEMA_signal_1059 ), .Q ( new_AGEMA_signal_5912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1437 ( .C ( clk ), .D ( n2442 ), .Q ( new_AGEMA_signal_5926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1441 ( .C ( clk ), .D ( new_AGEMA_signal_1148 ), .Q ( new_AGEMA_signal_5930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1445 ( .C ( clk ), .D ( new_AGEMA_signal_1149 ), .Q ( new_AGEMA_signal_5934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1515 ( .C ( clk ), .D ( n2779 ), .Q ( new_AGEMA_signal_6004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1519 ( .C ( clk ), .D ( new_AGEMA_signal_992 ), .Q ( new_AGEMA_signal_6008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1523 ( .C ( clk ), .D ( new_AGEMA_signal_993 ), .Q ( new_AGEMA_signal_6012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1569 ( .C ( clk ), .D ( n2721 ), .Q ( new_AGEMA_signal_6058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1573 ( .C ( clk ), .D ( new_AGEMA_signal_1080 ), .Q ( new_AGEMA_signal_6062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1577 ( .C ( clk ), .D ( new_AGEMA_signal_1081 ), .Q ( new_AGEMA_signal_6066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1611 ( .C ( clk ), .D ( n2823 ), .Q ( new_AGEMA_signal_6100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1615 ( .C ( clk ), .D ( new_AGEMA_signal_1184 ), .Q ( new_AGEMA_signal_6104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1619 ( .C ( clk ), .D ( new_AGEMA_signal_1185 ), .Q ( new_AGEMA_signal_6108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1641 ( .C ( clk ), .D ( n2346 ), .Q ( new_AGEMA_signal_6130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1645 ( .C ( clk ), .D ( new_AGEMA_signal_1084 ), .Q ( new_AGEMA_signal_6134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1649 ( .C ( clk ), .D ( new_AGEMA_signal_1085 ), .Q ( new_AGEMA_signal_6138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1671 ( .C ( clk ), .D ( n2315 ), .Q ( new_AGEMA_signal_6160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1675 ( .C ( clk ), .D ( new_AGEMA_signal_980 ), .Q ( new_AGEMA_signal_6164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1679 ( .C ( clk ), .D ( new_AGEMA_signal_981 ), .Q ( new_AGEMA_signal_6168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C ( clk ), .D ( new_AGEMA_signal_6275 ), .Q ( new_AGEMA_signal_6276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C ( clk ), .D ( new_AGEMA_signal_6281 ), .Q ( new_AGEMA_signal_6282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C ( clk ), .D ( new_AGEMA_signal_6287 ), .Q ( new_AGEMA_signal_6288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C ( clk ), .D ( new_AGEMA_signal_5429 ), .Q ( new_AGEMA_signal_6310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C ( clk ), .D ( new_AGEMA_signal_5431 ), .Q ( new_AGEMA_signal_6314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C ( clk ), .D ( new_AGEMA_signal_5433 ), .Q ( new_AGEMA_signal_6318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C ( clk ), .D ( n2600 ), .Q ( new_AGEMA_signal_6340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C ( clk ), .D ( new_AGEMA_signal_1026 ), .Q ( new_AGEMA_signal_6344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C ( clk ), .D ( new_AGEMA_signal_1027 ), .Q ( new_AGEMA_signal_6348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C ( clk ), .D ( n2750 ), .Q ( new_AGEMA_signal_6394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C ( clk ), .D ( new_AGEMA_signal_1002 ), .Q ( new_AGEMA_signal_6398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C ( clk ), .D ( new_AGEMA_signal_1003 ), .Q ( new_AGEMA_signal_6402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C ( clk ), .D ( new_AGEMA_signal_5471 ), .Q ( new_AGEMA_signal_6418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C ( clk ), .D ( new_AGEMA_signal_5473 ), .Q ( new_AGEMA_signal_6422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C ( clk ), .D ( new_AGEMA_signal_5475 ), .Q ( new_AGEMA_signal_6426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2151 ( .C ( clk ), .D ( n2737 ), .Q ( new_AGEMA_signal_6640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C ( clk ), .D ( new_AGEMA_signal_1108 ), .Q ( new_AGEMA_signal_6646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2163 ( .C ( clk ), .D ( new_AGEMA_signal_1109 ), .Q ( new_AGEMA_signal_6652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2229 ( .C ( clk ), .D ( n2785 ), .Q ( new_AGEMA_signal_6718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2235 ( .C ( clk ), .D ( new_AGEMA_signal_1036 ), .Q ( new_AGEMA_signal_6724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2241 ( .C ( clk ), .D ( new_AGEMA_signal_1037 ), .Q ( new_AGEMA_signal_6730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2577 ( .C ( clk ), .D ( n2595 ), .Q ( new_AGEMA_signal_7066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2585 ( .C ( clk ), .D ( new_AGEMA_signal_984 ), .Q ( new_AGEMA_signal_7074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2593 ( .C ( clk ), .D ( new_AGEMA_signal_985 ), .Q ( new_AGEMA_signal_7082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2607 ( .C ( clk ), .D ( n2437 ), .Q ( new_AGEMA_signal_7096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2615 ( .C ( clk ), .D ( new_AGEMA_signal_1050 ), .Q ( new_AGEMA_signal_7104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2623 ( .C ( clk ), .D ( new_AGEMA_signal_1051 ), .Q ( new_AGEMA_signal_7112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2835 ( .C ( clk ), .D ( n2828 ), .Q ( new_AGEMA_signal_7324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2843 ( .C ( clk ), .D ( new_AGEMA_signal_1188 ), .Q ( new_AGEMA_signal_7332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2851 ( .C ( clk ), .D ( new_AGEMA_signal_1189 ), .Q ( new_AGEMA_signal_7340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3093 ( .C ( clk ), .D ( n2538 ), .Q ( new_AGEMA_signal_7582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3101 ( .C ( clk ), .D ( new_AGEMA_signal_1028 ), .Q ( new_AGEMA_signal_7590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3109 ( .C ( clk ), .D ( new_AGEMA_signal_1029 ), .Q ( new_AGEMA_signal_7598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3183 ( .C ( clk ), .D ( n2809 ), .Q ( new_AGEMA_signal_7672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3191 ( .C ( clk ), .D ( new_AGEMA_signal_1192 ), .Q ( new_AGEMA_signal_7680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3199 ( .C ( clk ), .D ( new_AGEMA_signal_1193 ), .Q ( new_AGEMA_signal_7688 ) ) ;

    /* cells in depth 4 */
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1954 ( .a ({new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2750}), .b ({new_AGEMA_signal_1107, new_AGEMA_signal_1106, n2640}), .clk ( clk ), .r ({Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, n2575}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1959 ( .a ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, n2737}), .b ({new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2767}), .clk ( clk ), .r ({Fresh[161], Fresh[160], Fresh[159]}), .c ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, n1962}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1964 ( .a ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, n2789}), .b ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, n2317}), .clk ( clk ), .r ({Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, n1922}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1974 ( .a ({new_AGEMA_signal_981, new_AGEMA_signal_980, n2315}), .b ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2713}), .clk ( clk ), .r ({Fresh[167], Fresh[166], Fresh[165]}), .c ({new_AGEMA_signal_1119, new_AGEMA_signal_1118, n2755}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1977 ( .a ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, n2317}), .b ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, n2688}), .clk ( clk ), .r ({Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, n1926}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1980 ( .a ({new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2767}), .b ({new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2541}), .clk ( clk ), .r ({Fresh[173], Fresh[172], Fresh[171]}), .c ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, n1925}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1986 ( .a ({new_AGEMA_signal_1125, new_AGEMA_signal_1124, n2086}), .b ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, n2317}), .clk ( clk ), .r ({Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, n2151}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1988 ( .a ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, n2641}), .b ({new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2600}), .clk ( clk ), .r ({Fresh[179], Fresh[178], Fresh[177]}), .c ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, n2631}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U1989 ( .a ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, n2631}), .b ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, n2734}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1992 ( .a ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2707}), .b ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2786}), .clk ( clk ), .r ({Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2763}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1997 ( .a ({new_AGEMA_signal_979, new_AGEMA_signal_978, n2519}), .b ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, n2742}), .clk ( clk ), .r ({Fresh[185], Fresh[184], Fresh[183]}), .c ({new_AGEMA_signal_1131, new_AGEMA_signal_1130, n1930}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2005 ( .a ({new_AGEMA_signal_1035, new_AGEMA_signal_1034, n2400}), .b ({new_AGEMA_signal_979, new_AGEMA_signal_978, n2519}), .clk ( clk ), .r ({Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2492}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2006 ( .a ({new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2492}), .b ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, n2732}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2010 ( .a ({new_AGEMA_signal_5421, new_AGEMA_signal_5419, new_AGEMA_signal_5417}), .b ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, n2792}), .clk ( clk ), .r ({Fresh[191], Fresh[190], Fresh[189]}), .c ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, n1937}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2022 ( .a ({new_AGEMA_signal_5427, new_AGEMA_signal_5425, new_AGEMA_signal_5423}), .b ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, n2493}), .clk ( clk ), .r ({Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_1143, new_AGEMA_signal_1142, n1942}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) U2026 ( .a ({new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2587}), .b ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, n2815}), .clk ( clk ), .r ({Fresh[197], Fresh[196], Fresh[195]}), .c ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, n2676}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2030 ( .a ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, n2789}), .b ({new_AGEMA_signal_989, new_AGEMA_signal_988, n2559}), .clk ( clk ), .r ({Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, n1944}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2037 ( .a ({new_AGEMA_signal_1023, new_AGEMA_signal_1022, n2725}), .b ({new_AGEMA_signal_1115, new_AGEMA_signal_1114, n2769}), .clk ( clk ), .r ({Fresh[203], Fresh[202], Fresh[201]}), .c ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, n1950}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2039 ( .a ({new_AGEMA_signal_5433, new_AGEMA_signal_5431, new_AGEMA_signal_5429}), .b ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, n2739}), .clk ( clk ), .r ({Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_1151, new_AGEMA_signal_1150, n1949}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2042 ( .a ({new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2750}), .b ({new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2600}), .clk ( clk ), .r ({Fresh[209], Fresh[208], Fresh[207]}), .c ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, n2677}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2043 ( .a ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, n2677}), .b ({new_AGEMA_signal_1341, new_AGEMA_signal_1340, n2662}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2047 ( .a ({new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2437}), .b ({new_AGEMA_signal_1053, new_AGEMA_signal_1052, n2778}), .clk ( clk ), .r ({Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_1155, new_AGEMA_signal_1154, n2627}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2053 ( .a ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2816}), .b ({new_AGEMA_signal_1055, new_AGEMA_signal_1054, n2452}), .clk ( clk ), .r ({Fresh[215], Fresh[214], Fresh[213]}), .c ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, n1957}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2056 ( .a ({new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2766}), .b ({new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2600}), .clk ( clk ), .r ({Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, n2088}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2062 ( .a ({new_AGEMA_signal_979, new_AGEMA_signal_978, n2519}), .b ({new_AGEMA_signal_987, new_AGEMA_signal_986, n2708}), .clk ( clk ), .r ({Fresh[221], Fresh[220], Fresh[219]}), .c ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, n1964}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2063 ( .a ({new_AGEMA_signal_5439, new_AGEMA_signal_5437, new_AGEMA_signal_5435}), .b ({new_AGEMA_signal_1047, new_AGEMA_signal_1046, n2643}), .clk ( clk ), .r ({Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, n2736}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2069 ( .a ({new_AGEMA_signal_1059, new_AGEMA_signal_1058, n2772}), .b ({new_AGEMA_signal_5445, new_AGEMA_signal_5443, new_AGEMA_signal_5441}), .clk ( clk ), .r ({Fresh[227], Fresh[226], Fresh[225]}), .c ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, n2673}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2072 ( .a ({new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2766}), .b ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, n2612}), .clk ( clk ), .r ({Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, n2761}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2073 ( .a ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, n2761}), .b ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, n2720}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2075 ( .a ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, n2313}), .b ({new_AGEMA_signal_999, new_AGEMA_signal_998, n2719}), .clk ( clk ), .r ({Fresh[233], Fresh[232], Fresh[231]}), .c ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, n2412}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2076 ( .a ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, n2412}), .b ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, n2417}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2079 ( .a ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, n2641}), .b ({new_AGEMA_signal_991, new_AGEMA_signal_990, n2261}), .clk ( clk ), .r ({Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, n2571}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2080 ( .a ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, n2571}), .b ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, n2505}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2081 ( .a ({new_AGEMA_signal_979, new_AGEMA_signal_978, n2519}), .b ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, n2824}), .clk ( clk ), .r ({Fresh[239], Fresh[238], Fresh[237]}), .c ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2651}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2083 ( .a ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, n2792}), .b ({new_AGEMA_signal_5445, new_AGEMA_signal_5443, new_AGEMA_signal_5441}), .clk ( clk ), .r ({Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_1353, new_AGEMA_signal_1352, n2359}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2086 ( .a ({new_AGEMA_signal_979, new_AGEMA_signal_978, n2519}), .b ({new_AGEMA_signal_1053, new_AGEMA_signal_1052, n2778}), .clk ( clk ), .r ({Fresh[245], Fresh[244], Fresh[243]}), .c ({new_AGEMA_signal_1173, new_AGEMA_signal_1172, n2101}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2087 ( .a ({new_AGEMA_signal_1173, new_AGEMA_signal_1172, n2101}), .b ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, n2625}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2091 ( .a ({new_AGEMA_signal_999, new_AGEMA_signal_998, n2719}), .b ({new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2609}), .clk ( clk ), .r ({Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_1177, new_AGEMA_signal_1176, n2190}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2095 ( .a ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, n2739}), .b ({new_AGEMA_signal_993, new_AGEMA_signal_992, n2779}), .clk ( clk ), .r ({Fresh[251], Fresh[250], Fresh[249]}), .c ({new_AGEMA_signal_1179, new_AGEMA_signal_1178, n1976}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2098 ( .a ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2672}), .b ({new_AGEMA_signal_995, new_AGEMA_signal_994, n2242}), .clk ( clk ), .r ({Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_1359, new_AGEMA_signal_1358, n2535}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2101 ( .a ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, n2688}), .b ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, n2356}), .clk ( clk ), .r ({Fresh[257], Fresh[256], Fresh[255]}), .c ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, n1973}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2105 ( .a ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, n2815}), .b ({new_AGEMA_signal_981, new_AGEMA_signal_980, n2315}), .clk ( clk ), .r ({Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, n2690}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2111 ( .a ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, n2493}), .b ({new_AGEMA_signal_5451, new_AGEMA_signal_5449, new_AGEMA_signal_5447}), .clk ( clk ), .r ({Fresh[263], Fresh[262], Fresh[261]}), .c ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2817}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2113 ( .a ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, n2442}), .b ({new_AGEMA_signal_993, new_AGEMA_signal_992, n2779}), .clk ( clk ), .r ({Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_1365, new_AGEMA_signal_1364, n2741}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2118 ( .a ({new_AGEMA_signal_1011, new_AGEMA_signal_1010, n2780}), .b ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, n2818}), .clk ( clk ), .r ({Fresh[269], Fresh[268], Fresh[267]}), .c ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, n1992}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2120 ( .a ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, n2823}), .b ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2672}), .clk ( clk ), .r ({Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, n1991}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2123 ( .a ({new_AGEMA_signal_1047, new_AGEMA_signal_1046, n2643}), .b ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2611}), .clk ( clk ), .r ({Fresh[275], Fresh[274], Fresh[273]}), .c ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, n1993}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2125 ( .a ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, n2737}), .b ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, n2792}), .clk ( clk ), .r ({Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_1371, new_AGEMA_signal_1370, n1995}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2132 ( .a ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, n2818}), .b ({new_AGEMA_signal_987, new_AGEMA_signal_986, n2708}), .clk ( clk ), .r ({Fresh[281], Fresh[280], Fresh[279]}), .c ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, n2241}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2135 ( .a ({new_AGEMA_signal_5457, new_AGEMA_signal_5455, new_AGEMA_signal_5453}), .b ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, n2679}), .clk ( clk ), .r ({Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, n2003}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2140 ( .a ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, n2612}), .b ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, n2809}), .clk ( clk ), .r ({Fresh[287], Fresh[286], Fresh[285]}), .c ({new_AGEMA_signal_1377, new_AGEMA_signal_1376, n2008}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2141 ( .a ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, n2679}), .b ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, n2688}), .clk ( clk ), .r ({Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, n2572}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2143 ( .a ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, n2809}), .b ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, n2356}), .clk ( clk ), .r ({Fresh[293], Fresh[292], Fresh[291]}), .c ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, n2004}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2147 ( .a ({new_AGEMA_signal_975, new_AGEMA_signal_974, n2635}), .b ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2672}), .clk ( clk ), .r ({Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_1383, new_AGEMA_signal_1382, n2009}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2151 ( .a ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, n2789}), .b ({new_AGEMA_signal_5451, new_AGEMA_signal_5449, new_AGEMA_signal_5447}), .clk ( clk ), .r ({Fresh[299], Fresh[298], Fresh[297]}), .c ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, n2533}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2157 ( .a ({new_AGEMA_signal_999, new_AGEMA_signal_998, n2719}), .b ({new_AGEMA_signal_983, new_AGEMA_signal_982, n2682}), .clk ( clk ), .r ({Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_1197, new_AGEMA_signal_1196, n2026}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2158 ( .a ({new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2766}), .b ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, n2493}), .clk ( clk ), .r ({Fresh[305], Fresh[304], Fresh[303]}), .c ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, n2022}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2159 ( .a ({new_AGEMA_signal_5463, new_AGEMA_signal_5461, new_AGEMA_signal_5459}), .b ({new_AGEMA_signal_1023, new_AGEMA_signal_1022, n2725}), .clk ( clk ), .r ({Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, n2227}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2167 ( .a ({new_AGEMA_signal_977, new_AGEMA_signal_976, n2790}), .b ({new_AGEMA_signal_5451, new_AGEMA_signal_5449, new_AGEMA_signal_5447}), .clk ( clk ), .r ({Fresh[311], Fresh[310], Fresh[309]}), .c ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, n2027}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2171 ( .a ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, n2818}), .b ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, n2442}), .clk ( clk ), .r ({Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, n2214}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2173 ( .a ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, n2442}), .b ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2707}), .clk ( clk ), .r ({Fresh[317], Fresh[316], Fresh[315]}), .c ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, n2290}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2174 ( .a ({new_AGEMA_signal_5439, new_AGEMA_signal_5437, new_AGEMA_signal_5435}), .b ({new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2767}), .clk ( clk ), .r ({Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, n2376}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2178 ( .a ({new_AGEMA_signal_987, new_AGEMA_signal_986, n2708}), .b ({new_AGEMA_signal_1035, new_AGEMA_signal_1034, n2400}), .clk ( clk ), .r ({Fresh[323], Fresh[322], Fresh[321]}), .c ({new_AGEMA_signal_1203, new_AGEMA_signal_1202, n2034}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2182 ( .a ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2611}), .b ({new_AGEMA_signal_999, new_AGEMA_signal_998, n2719}), .clk ( clk ), .r ({Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, n2171}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2183 ( .a ({new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2828}), .b ({new_AGEMA_signal_1115, new_AGEMA_signal_1114, n2769}), .clk ( clk ), .r ({Fresh[329], Fresh[328], Fresh[327]}), .c ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2039}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2188 ( .a ({new_AGEMA_signal_1023, new_AGEMA_signal_1022, n2725}), .b ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2707}), .clk ( clk ), .r ({Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, n2042}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2191 ( .a ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2707}), .b ({new_AGEMA_signal_981, new_AGEMA_signal_980, n2315}), .clk ( clk ), .r ({Fresh[335], Fresh[334], Fresh[333]}), .c ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, n2754}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2192 ( .a ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, n2313}), .b ({new_AGEMA_signal_977, new_AGEMA_signal_976, n2790}), .clk ( clk ), .r ({Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_1407, new_AGEMA_signal_1406, n2044}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2198 ( .a ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, n2313}), .b ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, n2641}), .clk ( clk ), .r ({Fresh[341], Fresh[340], Fresh[339]}), .c ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, n2654}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2202 ( .a ({new_AGEMA_signal_975, new_AGEMA_signal_974, n2635}), .b ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, n2577}), .clk ( clk ), .r ({Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, n2055}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2205 ( .a ({new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2395}), .b ({new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2767}), .clk ( clk ), .r ({Fresh[347], Fresh[346], Fresh[345]}), .c ({new_AGEMA_signal_1413, new_AGEMA_signal_1412, n2057}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2208 ( .a ({new_AGEMA_signal_1191, new_AGEMA_signal_1190, n2679}), .b ({new_AGEMA_signal_983, new_AGEMA_signal_982, n2682}), .clk ( clk ), .r ({Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, n2407}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2212 ( .a ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, n2688}), .b ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, n2061}), .clk ( clk ), .r ({Fresh[353], Fresh[352], Fresh[351]}), .c ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, n2062}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2216 ( .a ({new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2766}), .b ({new_AGEMA_signal_989, new_AGEMA_signal_988, n2559}), .clk ( clk ), .r ({Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_1419, new_AGEMA_signal_1418, n2731}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2220 ( .a ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, n2690}), .b ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, n2068}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2224 ( .a ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2611}), .b ({new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2750}), .clk ( clk ), .r ({Fresh[359], Fresh[358], Fresh[357]}), .c ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, n2642}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2225 ( .a ({new_AGEMA_signal_1023, new_AGEMA_signal_1022, n2725}), .b ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2786}), .clk ( clk ), .r ({Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, n2252}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2228 ( .a ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, n2739}), .b ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, n2815}), .clk ( clk ), .r ({Fresh[365], Fresh[364], Fresh[363]}), .c ({new_AGEMA_signal_1209, new_AGEMA_signal_1208, n2075}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) U2233 ( .a ({new_AGEMA_signal_975, new_AGEMA_signal_974, n2635}), .b ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2723}), .clk ( clk ), .r ({Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, n2081}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2234 ( .a ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, n2792}), .b ({new_AGEMA_signal_983, new_AGEMA_signal_982, n2682}), .clk ( clk ), .r ({Fresh[371], Fresh[370], Fresh[369]}), .c ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, n2080}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2237 ( .a ({new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2600}), .b ({new_AGEMA_signal_999, new_AGEMA_signal_998, n2719}), .clk ( clk ), .r ({Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, n2498}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2238 ( .a ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, n2498}), .b ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, n2773}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2239 ( .a ({new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2767}), .b ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, n2792}), .clk ( clk ), .r ({Fresh[377], Fresh[376], Fresh[375]}), .c ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, n2083}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2244 ( .a ({new_AGEMA_signal_5457, new_AGEMA_signal_5455, new_AGEMA_signal_5453}), .b ({new_AGEMA_signal_1125, new_AGEMA_signal_1124, n2086}), .clk ( clk ), .r ({Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_1431, new_AGEMA_signal_1430, n2562}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2247 ( .a ({new_AGEMA_signal_5439, new_AGEMA_signal_5437, new_AGEMA_signal_5435}), .b ({new_AGEMA_signal_1041, new_AGEMA_signal_1040, n2661}), .clk ( clk ), .r ({Fresh[383], Fresh[382], Fresh[381]}), .c ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, n2087}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2251 ( .a ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, n2563}), .b ({new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2174}), .clk ( clk ), .r ({Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, n2156}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2260 ( .a ({new_AGEMA_signal_1115, new_AGEMA_signal_1114, n2769}), .b ({new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2401}), .clk ( clk ), .r ({Fresh[389], Fresh[388], Fresh[387]}), .c ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, n2100}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2277 ( .a ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, n2739}), .b ({new_AGEMA_signal_1083, new_AGEMA_signal_1082, n2298}), .clk ( clk ), .r ({Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, n2544}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2279 ( .a ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, n2356}), .b ({new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2118}), .clk ( clk ), .r ({Fresh[395], Fresh[394], Fresh[393]}), .c ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, n2121}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2284 ( .a ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2707}), .b ({new_AGEMA_signal_1147, new_AGEMA_signal_1146, n2570}), .clk ( clk ), .r ({Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, n2122}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2286 ( .a ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, n2792}), .b ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, n2612}), .clk ( clk ), .r ({Fresh[401], Fresh[400], Fresh[399]}), .c ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, n2811}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2294 ( .a ({new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2437}), .b ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, n2742}), .clk ( clk ), .r ({Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_1221, new_AGEMA_signal_1220, n2647}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2297 ( .a ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, n2742}), .b ({new_AGEMA_signal_981, new_AGEMA_signal_980, n2315}), .clk ( clk ), .r ({Fresh[407], Fresh[406], Fresh[405]}), .c ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, n2132}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2304 ( .a ({new_AGEMA_signal_1071, new_AGEMA_signal_1070, n2616}), .b ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2707}), .clk ( clk ), .r ({Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, n2220}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2305 ( .a ({new_AGEMA_signal_5421, new_AGEMA_signal_5419, new_AGEMA_signal_5417}), .b ({new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2767}), .clk ( clk ), .r ({Fresh[413], Fresh[412], Fresh[411]}), .c ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, n2138}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2312 ( .a ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, n2612}), .b ({new_AGEMA_signal_5469, new_AGEMA_signal_5467, new_AGEMA_signal_5465}), .clk ( clk ), .r ({Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, n2555}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2322 ( .a ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, n2612}), .b ({new_AGEMA_signal_5475, new_AGEMA_signal_5473, new_AGEMA_signal_5471}), .clk ( clk ), .r ({Fresh[419], Fresh[418], Fresh[417]}), .c ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, n2429}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2328 ( .a ({new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2437}), .b ({new_AGEMA_signal_5451, new_AGEMA_signal_5449, new_AGEMA_signal_5447}), .clk ( clk ), .r ({Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_1225, new_AGEMA_signal_1224, n2162}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2337 ( .a ({new_AGEMA_signal_981, new_AGEMA_signal_980, n2315}), .b ({new_AGEMA_signal_995, new_AGEMA_signal_994, n2242}), .clk ( clk ), .r ({Fresh[425], Fresh[424], Fresh[423]}), .c ({new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2545}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2340 ( .a ({new_AGEMA_signal_989, new_AGEMA_signal_988, n2559}), .b ({new_AGEMA_signal_1047, new_AGEMA_signal_1046, n2643}), .clk ( clk ), .r ({Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, n2178}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2342 ( .a ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, n2430}), .b ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2707}), .clk ( clk ), .r ({Fresh[431], Fresh[430], Fresh[429]}), .c ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, n2176}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2343 ( .a ({new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2174}), .b ({new_AGEMA_signal_5457, new_AGEMA_signal_5455, new_AGEMA_signal_5453}), .clk ( clk ), .r ({Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, n2175}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2348 ( .a ({new_AGEMA_signal_991, new_AGEMA_signal_990, n2261}), .b ({new_AGEMA_signal_5475, new_AGEMA_signal_5473, new_AGEMA_signal_5471}), .clk ( clk ), .r ({Fresh[437], Fresh[436], Fresh[435]}), .c ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, n2182}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2353 ( .a ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2786}), .b ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, n2430}), .clk ( clk ), .r ({Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, n2188}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2355 ( .a ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, n2792}), .b ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, n2612}), .clk ( clk ), .r ({Fresh[443], Fresh[442], Fresh[441]}), .c ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, n2189}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2357 ( .a ({new_AGEMA_signal_975, new_AGEMA_signal_974, n2635}), .b ({new_AGEMA_signal_1115, new_AGEMA_signal_1114, n2769}), .clk ( clk ), .r ({Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, n2446}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2362 ( .a ({new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2750}), .b ({new_AGEMA_signal_989, new_AGEMA_signal_988, n2559}), .clk ( clk ), .r ({Fresh[449], Fresh[448], Fresh[447]}), .c ({new_AGEMA_signal_1233, new_AGEMA_signal_1232, n2576}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2363 ( .a ({new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2609}), .b ({new_AGEMA_signal_5481, new_AGEMA_signal_5479, new_AGEMA_signal_5477}), .clk ( clk ), .r ({Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, n2748}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) U2368 ( .a ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, n2654}), .b ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, n2674}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2378 ( .a ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, n2815}), .b ({new_AGEMA_signal_987, new_AGEMA_signal_986, n2708}), .clk ( clk ), .r ({Fresh[455], Fresh[454], Fresh[453]}), .c ({new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2213}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2380 ( .a ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2816}), .b ({new_AGEMA_signal_5439, new_AGEMA_signal_5437, new_AGEMA_signal_5435}), .clk ( clk ), .r ({Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, n2215}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2384 ( .a ({new_AGEMA_signal_997, new_AGEMA_signal_996, n2712}), .b ({new_AGEMA_signal_1115, new_AGEMA_signal_1114, n2769}), .clk ( clk ), .r ({Fresh[461], Fresh[460], Fresh[459]}), .c ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, n2218}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2386 ( .a ({new_AGEMA_signal_1083, new_AGEMA_signal_1082, n2298}), .b ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2672}), .clk ( clk ), .r ({Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, n2219}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2405 ( .a ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2707}), .b ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2713}), .clk ( clk ), .r ({Fresh[467], Fresh[466], Fresh[465]}), .c ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, n2240}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2407 ( .a ({new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2709}), .b ({new_AGEMA_signal_995, new_AGEMA_signal_994, n2242}), .clk ( clk ), .r ({Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, n2561}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2408 ( .a ({new_AGEMA_signal_5457, new_AGEMA_signal_5455, new_AGEMA_signal_5453}), .b ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, n2442}), .clk ( clk ), .r ({Fresh[473], Fresh[472], Fresh[471]}), .c ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, n2243}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2411 ( .a ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, n2615}), .b ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, n2442}), .clk ( clk ), .r ({Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, n2245}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2422 ( .a ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2672}), .b ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, n2430}), .clk ( clk ), .r ({Fresh[479], Fresh[478], Fresh[477]}), .c ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, n2540}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2423 ( .a ({new_AGEMA_signal_991, new_AGEMA_signal_990, n2261}), .b ({new_AGEMA_signal_1107, new_AGEMA_signal_1106, n2640}), .clk ( clk ), .r ({Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_1503, new_AGEMA_signal_1502, n2259}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2426 ( .a ({new_AGEMA_signal_991, new_AGEMA_signal_990, n2261}), .b ({new_AGEMA_signal_1041, new_AGEMA_signal_1040, n2661}), .clk ( clk ), .r ({Fresh[485], Fresh[484], Fresh[483]}), .c ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, n2262}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2431 ( .a ({new_AGEMA_signal_981, new_AGEMA_signal_980, n2315}), .b ({new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2777}), .clk ( clk ), .r ({Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_1243, new_AGEMA_signal_1242, n2266}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2432 ( .a ({new_AGEMA_signal_1059, new_AGEMA_signal_1058, n2772}), .b ({new_AGEMA_signal_5475, new_AGEMA_signal_5473, new_AGEMA_signal_5471}), .clk ( clk ), .r ({Fresh[491], Fresh[490], Fresh[489]}), .c ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, n2645}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2436 ( .a ({new_AGEMA_signal_5421, new_AGEMA_signal_5419, new_AGEMA_signal_5417}), .b ({new_AGEMA_signal_1023, new_AGEMA_signal_1022, n2725}), .clk ( clk ), .r ({Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, n2268}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2443 ( .a ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2816}), .b ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2786}), .clk ( clk ), .r ({Fresh[497], Fresh[496], Fresh[495]}), .c ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, n2278}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2448 ( .a ({new_AGEMA_signal_5487, new_AGEMA_signal_5485, new_AGEMA_signal_5483}), .b ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2713}), .clk ( clk ), .r ({Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2383}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2455 ( .a ({new_AGEMA_signal_1053, new_AGEMA_signal_1052, n2778}), .b ({new_AGEMA_signal_1147, new_AGEMA_signal_1146, n2570}), .clk ( clk ), .r ({Fresh[503], Fresh[502], Fresh[501]}), .c ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, n2774}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2458 ( .a ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, n2823}), .b ({new_AGEMA_signal_1053, new_AGEMA_signal_1052, n2778}), .clk ( clk ), .r ({Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, n2287}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2470 ( .a ({new_AGEMA_signal_979, new_AGEMA_signal_978, n2519}), .b ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2707}), .clk ( clk ), .r ({Fresh[509], Fresh[508], Fresh[507]}), .c ({new_AGEMA_signal_1521, new_AGEMA_signal_1520, n2438}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2471 ( .a ({new_AGEMA_signal_1083, new_AGEMA_signal_1082, n2298}), .b ({new_AGEMA_signal_981, new_AGEMA_signal_980, n2315}), .clk ( clk ), .r ({Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, n2299}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2481 ( .a ({new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2766}), .b ({new_AGEMA_signal_1167, new_AGEMA_signal_1166, n2313}), .clk ( clk ), .r ({Fresh[515], Fresh[514], Fresh[513]}), .c ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, n2371}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2484 ( .a ({new_AGEMA_signal_981, new_AGEMA_signal_980, n2315}), .b ({new_AGEMA_signal_979, new_AGEMA_signal_978, n2519}), .clk ( clk ), .r ({Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_1095, new_AGEMA_signal_1094, n2316}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2486 ( .a ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, n2624}), .b ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, n2317}), .clk ( clk ), .r ({Fresh[521], Fresh[520], Fresh[519]}), .c ({new_AGEMA_signal_1255, new_AGEMA_signal_1254, n2318}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2492 ( .a ({new_AGEMA_signal_987, new_AGEMA_signal_986, n2708}), .b ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2672}), .clk ( clk ), .r ({Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, n2325}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2494 ( .a ({new_AGEMA_signal_987, new_AGEMA_signal_986, n2708}), .b ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2707}), .clk ( clk ), .r ({Fresh[527], Fresh[526], Fresh[525]}), .c ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, n2328}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2495 ( .a ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, n2742}), .b ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2723}), .clk ( clk ), .r ({Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_1257, new_AGEMA_signal_1256, n2327}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2505 ( .a ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, n2737}), .b ({new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2694}), .clk ( clk ), .r ({Fresh[533], Fresh[532], Fresh[531]}), .c ({new_AGEMA_signal_1533, new_AGEMA_signal_1532, n2343}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2510 ( .a ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, n2563}), .b ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2672}), .clk ( clk ), .r ({Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, n2344}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) U2512 ( .a ({new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2395}), .b ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, n2346}), .clk ( clk ), .r ({Fresh[539], Fresh[538], Fresh[537]}), .c ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, n2348}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2513 ( .a ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, n2742}), .b ({new_AGEMA_signal_1011, new_AGEMA_signal_1010, n2780}), .clk ( clk ), .r ({Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2347}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2520 ( .a ({new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2694}), .b ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2753}), .clk ( clk ), .r ({Fresh[545], Fresh[544], Fresh[543]}), .c ({new_AGEMA_signal_1263, new_AGEMA_signal_1262, n2363}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2521 ( .a ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, n2809}), .b ({new_AGEMA_signal_5445, new_AGEMA_signal_5443, new_AGEMA_signal_5441}), .clk ( clk ), .r ({Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, n2353}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2524 ( .a ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, n2818}), .b ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2713}), .clk ( clk ), .r ({Fresh[551], Fresh[550], Fresh[549]}), .c ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, n2355}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2530 ( .a ({new_AGEMA_signal_997, new_AGEMA_signal_996, n2712}), .b ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2672}), .clk ( clk ), .r ({Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2364}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2543 ( .a ({new_AGEMA_signal_5421, new_AGEMA_signal_5419, new_AGEMA_signal_5417}), .b ({new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2401}), .clk ( clk ), .r ({Fresh[557], Fresh[556], Fresh[555]}), .c ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, n2415}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2558 ( .a ({new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2395}), .b ({new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2750}), .clk ( clk ), .r ({Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2700}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2563 ( .a ({new_AGEMA_signal_5493, new_AGEMA_signal_5491, new_AGEMA_signal_5489}), .b ({new_AGEMA_signal_1035, new_AGEMA_signal_1034, n2400}), .clk ( clk ), .r ({Fresh[563], Fresh[562], Fresh[561]}), .c ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, n2594}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2564 ( .a ({new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2401}), .b ({new_AGEMA_signal_5451, new_AGEMA_signal_5449, new_AGEMA_signal_5447}), .clk ( clk ), .r ({Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, n2402}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2585 ( .a ({new_AGEMA_signal_997, new_AGEMA_signal_996, n2712}), .b ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, n2823}), .clk ( clk ), .r ({Fresh[569], Fresh[568], Fresh[567]}), .c ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, n2428}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2588 ( .a ({new_AGEMA_signal_1089, new_AGEMA_signal_1088, n2430}), .b ({new_AGEMA_signal_1147, new_AGEMA_signal_1146, n2570}), .clk ( clk ), .r ({Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, n2431}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2594 ( .a ({new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2437}), .b ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, n2615}), .clk ( clk ), .r ({Fresh[575], Fresh[574], Fresh[573]}), .c ({new_AGEMA_signal_1273, new_AGEMA_signal_1272, n2483}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2599 ( .a ({new_AGEMA_signal_1149, new_AGEMA_signal_1148, n2442}), .b ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2713}), .clk ( clk ), .r ({Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, n2443}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2606 ( .a ({new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2766}), .b ({new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2609}), .clk ( clk ), .r ({Fresh[581], Fresh[580], Fresh[579]}), .c ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, n2693}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2608 ( .a ({new_AGEMA_signal_1055, new_AGEMA_signal_1054, n2452}), .b ({new_AGEMA_signal_5499, new_AGEMA_signal_5497, new_AGEMA_signal_5495}), .clk ( clk ), .r ({Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_1275, new_AGEMA_signal_1274, n2453}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2616 ( .a ({new_AGEMA_signal_977, new_AGEMA_signal_976, n2790}), .b ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, n2463}), .clk ( clk ), .r ({Fresh[587], Fresh[586], Fresh[585]}), .c ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, n2464}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2620 ( .a ({new_AGEMA_signal_1023, new_AGEMA_signal_1022, n2725}), .b ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, n2742}), .clk ( clk ), .r ({Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2468}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2624 ( .a ({new_AGEMA_signal_1053, new_AGEMA_signal_1052, n2778}), .b ({new_AGEMA_signal_5445, new_AGEMA_signal_5443, new_AGEMA_signal_5441}), .clk ( clk ), .r ({Fresh[593], Fresh[592], Fresh[591]}), .c ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, n2473}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2625 ( .a ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, n2815}), .b ({new_AGEMA_signal_1011, new_AGEMA_signal_1010, n2780}), .clk ( clk ), .r ({Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, n2472}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2628 ( .a ({new_AGEMA_signal_1041, new_AGEMA_signal_1040, n2661}), .b ({new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2474}), .clk ( clk ), .r ({Fresh[599], Fresh[598], Fresh[597]}), .c ({new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2475}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2632 ( .a ({new_AGEMA_signal_5505, new_AGEMA_signal_5503, new_AGEMA_signal_5501}), .b ({new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2828}), .clk ( clk ), .r ({Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, n2480}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2638 ( .a ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, n2577}), .b ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, n2615}), .clk ( clk ), .r ({Fresh[605], Fresh[604], Fresh[603]}), .c ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, n2487}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2641 ( .a ({new_AGEMA_signal_1071, new_AGEMA_signal_1070, n2616}), .b ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, n2824}), .clk ( clk ), .r ({Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, n2488}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2665 ( .a ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2786}), .b ({new_AGEMA_signal_979, new_AGEMA_signal_978, n2519}), .clk ( clk ), .r ({Fresh[611], Fresh[610], Fresh[609]}), .c ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, n2520}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2667 ( .a ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2713}), .b ({new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2587}), .clk ( clk ), .r ({Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, n2521}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2674 ( .a ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, n2737}), .b ({new_AGEMA_signal_985, new_AGEMA_signal_984, n2595}), .clk ( clk ), .r ({Fresh[617], Fresh[616], Fresh[615]}), .c ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, n2531}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2689 ( .a ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, n2824}), .b ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, n2818}), .clk ( clk ), .r ({Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, n2553}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2691 ( .a ({new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2694}), .b ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, n2792}), .clk ( clk ), .r ({Fresh[623], Fresh[622], Fresh[621]}), .c ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, n2554}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) U2695 ( .a ({new_AGEMA_signal_989, new_AGEMA_signal_988, n2559}), .b ({new_AGEMA_signal_1047, new_AGEMA_signal_1046, n2643}), .clk ( clk ), .r ({Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2560}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2698 ( .a ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, n2724}), .b ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, n2563}), .clk ( clk ), .r ({Fresh[629], Fresh[628], Fresh[627]}), .c ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, n2564}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2714 ( .a ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, n2688}), .b ({new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2694}), .clk ( clk ), .r ({Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, n2586}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2720 ( .a ({new_AGEMA_signal_985, new_AGEMA_signal_984, n2595}), .b ({new_AGEMA_signal_1047, new_AGEMA_signal_1046, n2643}), .clk ( clk ), .r ({Fresh[635], Fresh[634], Fresh[633]}), .c ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, n2597}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2721 ( .a ({new_AGEMA_signal_1107, new_AGEMA_signal_1106, n2640}), .b ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, n2789}), .clk ( clk ), .r ({Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, n2596}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2723 ( .a ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, n2724}), .b ({new_AGEMA_signal_1011, new_AGEMA_signal_1010, n2780}), .clk ( clk ), .r ({Fresh[641], Fresh[640], Fresh[639]}), .c ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, n2598}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2725 ( .a ({new_AGEMA_signal_975, new_AGEMA_signal_974, n2635}), .b ({new_AGEMA_signal_5439, new_AGEMA_signal_5437, new_AGEMA_signal_5435}), .clk ( clk ), .r ({Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_1101, new_AGEMA_signal_1100, n2599}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2732 ( .a ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2707}), .b ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, n2818}), .clk ( clk ), .r ({Fresh[647], Fresh[646], Fresh[645]}), .c ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, n2610}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2734 ( .a ({new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2767}), .b ({new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2611}), .clk ( clk ), .r ({Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, n2614}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2735 ( .a ({new_AGEMA_signal_1165, new_AGEMA_signal_1164, n2612}), .b ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, n2789}), .clk ( clk ), .r ({Fresh[653], Fresh[652], Fresh[651]}), .c ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, n2613}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2737 ( .a ({new_AGEMA_signal_1071, new_AGEMA_signal_1070, n2616}), .b ({new_AGEMA_signal_1005, new_AGEMA_signal_1004, n2615}), .clk ( clk ), .r ({Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, n2617}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2742 ( .a ({new_AGEMA_signal_1065, new_AGEMA_signal_1064, n2624}), .b ({new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2750}), .clk ( clk ), .r ({Fresh[659], Fresh[658], Fresh[657]}), .c ({new_AGEMA_signal_1299, new_AGEMA_signal_1298, n2629}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2751 ( .a ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, n2641}), .b ({new_AGEMA_signal_1107, new_AGEMA_signal_1106, n2640}), .clk ( clk ), .r ({Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, n2784}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2757 ( .a ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, n2785}), .b ({new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2777}), .clk ( clk ), .r ({Fresh[665], Fresh[664], Fresh[663]}), .c ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, n2650}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2775 ( .a ({new_AGEMA_signal_5469, new_AGEMA_signal_5467, new_AGEMA_signal_5465}), .b ({new_AGEMA_signal_983, new_AGEMA_signal_982, n2682}), .clk ( clk ), .r ({Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, n2683}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2789 ( .a ({new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2723}), .b ({new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2707}), .clk ( clk ), .r ({Fresh[671], Fresh[670], Fresh[669]}), .c ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, n2711}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2790 ( .a ({new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2709}), .b ({new_AGEMA_signal_987, new_AGEMA_signal_986, n2708}), .clk ( clk ), .r ({Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, n2710}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2792 ( .a ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, n2713}), .b ({new_AGEMA_signal_997, new_AGEMA_signal_996, n2712}), .clk ( clk ), .r ({Fresh[677], Fresh[676], Fresh[675]}), .c ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2714}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2797 ( .a ({new_AGEMA_signal_977, new_AGEMA_signal_976, n2790}), .b ({new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2721}), .clk ( clk ), .r ({Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_1305, new_AGEMA_signal_1304, n2722}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2799 ( .a ({new_AGEMA_signal_1023, new_AGEMA_signal_1022, n2725}), .b ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, n2724}), .clk ( clk ), .r ({Fresh[683], Fresh[682], Fresh[681]}), .c ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, n2726}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2806 ( .a ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, n2737}), .b ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2753}), .clk ( clk ), .r ({Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, n2738}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2822 ( .a ({new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2767}), .b ({new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2766}), .clk ( clk ), .r ({Fresh[689], Fresh[688], Fresh[687]}), .c ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, n2768}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2828 ( .a ({new_AGEMA_signal_1053, new_AGEMA_signal_1052, n2778}), .b ({new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2777}), .clk ( clk ), .r ({Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, n2782}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2829 ( .a ({new_AGEMA_signal_1011, new_AGEMA_signal_1010, n2780}), .b ({new_AGEMA_signal_993, new_AGEMA_signal_992, n2779}), .clk ( clk ), .r ({Fresh[695], Fresh[694], Fresh[693]}), .c ({new_AGEMA_signal_1309, new_AGEMA_signal_1308, n2781}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2832 ( .a ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2786}), .b ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, n2785}), .clk ( clk ), .r ({Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, n2787}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2834 ( .a ({new_AGEMA_signal_977, new_AGEMA_signal_976, n2790}), .b ({new_AGEMA_signal_1113, new_AGEMA_signal_1112, n2789}), .clk ( clk ), .r ({Fresh[701], Fresh[700], Fresh[699]}), .c ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, n2794}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2835 ( .a ({new_AGEMA_signal_1137, new_AGEMA_signal_1136, n2792}), .b ({new_AGEMA_signal_5487, new_AGEMA_signal_5485, new_AGEMA_signal_5483}), .clk ( clk ), .r ({Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, n2793}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2844 ( .a ({new_AGEMA_signal_5505, new_AGEMA_signal_5503, new_AGEMA_signal_5501}), .b ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, n2809}), .clk ( clk ), .r ({Fresh[707], Fresh[706], Fresh[705]}), .c ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, n2812}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2847 ( .a ({new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2816}), .b ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, n2815}), .clk ( clk ), .r ({Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_1311, new_AGEMA_signal_1310, n2820}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2851 ( .a ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, n2824}), .b ({new_AGEMA_signal_1185, new_AGEMA_signal_1184, n2823}), .clk ( clk ), .r ({Fresh[713], Fresh[712], Fresh[711]}), .c ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, n2825}) ) ;
    buf_clk new_AGEMA_reg_buffer_1018 ( .C ( clk ), .D ( new_AGEMA_signal_5506 ), .Q ( new_AGEMA_signal_5507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1020 ( .C ( clk ), .D ( new_AGEMA_signal_5508 ), .Q ( new_AGEMA_signal_5509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1022 ( .C ( clk ), .D ( new_AGEMA_signal_5510 ), .Q ( new_AGEMA_signal_5511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1024 ( .C ( clk ), .D ( new_AGEMA_signal_5512 ), .Q ( new_AGEMA_signal_5513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1026 ( .C ( clk ), .D ( new_AGEMA_signal_5514 ), .Q ( new_AGEMA_signal_5515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1028 ( .C ( clk ), .D ( new_AGEMA_signal_5516 ), .Q ( new_AGEMA_signal_5517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1030 ( .C ( clk ), .D ( new_AGEMA_signal_5518 ), .Q ( new_AGEMA_signal_5519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1032 ( .C ( clk ), .D ( new_AGEMA_signal_5520 ), .Q ( new_AGEMA_signal_5521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1034 ( .C ( clk ), .D ( new_AGEMA_signal_5522 ), .Q ( new_AGEMA_signal_5523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1036 ( .C ( clk ), .D ( new_AGEMA_signal_5524 ), .Q ( new_AGEMA_signal_5525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1038 ( .C ( clk ), .D ( new_AGEMA_signal_5526 ), .Q ( new_AGEMA_signal_5527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1040 ( .C ( clk ), .D ( new_AGEMA_signal_5528 ), .Q ( new_AGEMA_signal_5529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1042 ( .C ( clk ), .D ( new_AGEMA_signal_5530 ), .Q ( new_AGEMA_signal_5531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1044 ( .C ( clk ), .D ( new_AGEMA_signal_5532 ), .Q ( new_AGEMA_signal_5533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1046 ( .C ( clk ), .D ( new_AGEMA_signal_5534 ), .Q ( new_AGEMA_signal_5535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1048 ( .C ( clk ), .D ( new_AGEMA_signal_5536 ), .Q ( new_AGEMA_signal_5537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1050 ( .C ( clk ), .D ( new_AGEMA_signal_5538 ), .Q ( new_AGEMA_signal_5539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1052 ( .C ( clk ), .D ( new_AGEMA_signal_5540 ), .Q ( new_AGEMA_signal_5541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1054 ( .C ( clk ), .D ( new_AGEMA_signal_5542 ), .Q ( new_AGEMA_signal_5543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1056 ( .C ( clk ), .D ( new_AGEMA_signal_5544 ), .Q ( new_AGEMA_signal_5545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1058 ( .C ( clk ), .D ( new_AGEMA_signal_5546 ), .Q ( new_AGEMA_signal_5547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1060 ( .C ( clk ), .D ( new_AGEMA_signal_5548 ), .Q ( new_AGEMA_signal_5549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1062 ( .C ( clk ), .D ( new_AGEMA_signal_5550 ), .Q ( new_AGEMA_signal_5551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1064 ( .C ( clk ), .D ( new_AGEMA_signal_5552 ), .Q ( new_AGEMA_signal_5553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1066 ( .C ( clk ), .D ( new_AGEMA_signal_5554 ), .Q ( new_AGEMA_signal_5555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1068 ( .C ( clk ), .D ( new_AGEMA_signal_5556 ), .Q ( new_AGEMA_signal_5557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1070 ( .C ( clk ), .D ( new_AGEMA_signal_5558 ), .Q ( new_AGEMA_signal_5559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1072 ( .C ( clk ), .D ( new_AGEMA_signal_5560 ), .Q ( new_AGEMA_signal_5561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1074 ( .C ( clk ), .D ( new_AGEMA_signal_5562 ), .Q ( new_AGEMA_signal_5563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1076 ( .C ( clk ), .D ( new_AGEMA_signal_5564 ), .Q ( new_AGEMA_signal_5565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1078 ( .C ( clk ), .D ( new_AGEMA_signal_5566 ), .Q ( new_AGEMA_signal_5567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1080 ( .C ( clk ), .D ( new_AGEMA_signal_5568 ), .Q ( new_AGEMA_signal_5569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1082 ( .C ( clk ), .D ( new_AGEMA_signal_5570 ), .Q ( new_AGEMA_signal_5571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1084 ( .C ( clk ), .D ( new_AGEMA_signal_5572 ), .Q ( new_AGEMA_signal_5573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1086 ( .C ( clk ), .D ( new_AGEMA_signal_5574 ), .Q ( new_AGEMA_signal_5575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1088 ( .C ( clk ), .D ( new_AGEMA_signal_5576 ), .Q ( new_AGEMA_signal_5577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1090 ( .C ( clk ), .D ( new_AGEMA_signal_5578 ), .Q ( new_AGEMA_signal_5579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1092 ( .C ( clk ), .D ( new_AGEMA_signal_5580 ), .Q ( new_AGEMA_signal_5581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1094 ( .C ( clk ), .D ( new_AGEMA_signal_5582 ), .Q ( new_AGEMA_signal_5583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1096 ( .C ( clk ), .D ( new_AGEMA_signal_5584 ), .Q ( new_AGEMA_signal_5585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1098 ( .C ( clk ), .D ( new_AGEMA_signal_5586 ), .Q ( new_AGEMA_signal_5587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1100 ( .C ( clk ), .D ( new_AGEMA_signal_5588 ), .Q ( new_AGEMA_signal_5589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1102 ( .C ( clk ), .D ( new_AGEMA_signal_5590 ), .Q ( new_AGEMA_signal_5591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1104 ( .C ( clk ), .D ( new_AGEMA_signal_5592 ), .Q ( new_AGEMA_signal_5593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1106 ( .C ( clk ), .D ( new_AGEMA_signal_5594 ), .Q ( new_AGEMA_signal_5595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1108 ( .C ( clk ), .D ( new_AGEMA_signal_5596 ), .Q ( new_AGEMA_signal_5597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1110 ( .C ( clk ), .D ( new_AGEMA_signal_5598 ), .Q ( new_AGEMA_signal_5599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1112 ( .C ( clk ), .D ( new_AGEMA_signal_5600 ), .Q ( new_AGEMA_signal_5601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1114 ( .C ( clk ), .D ( new_AGEMA_signal_5602 ), .Q ( new_AGEMA_signal_5603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1116 ( .C ( clk ), .D ( new_AGEMA_signal_5604 ), .Q ( new_AGEMA_signal_5605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1118 ( .C ( clk ), .D ( new_AGEMA_signal_5606 ), .Q ( new_AGEMA_signal_5607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1120 ( .C ( clk ), .D ( new_AGEMA_signal_5608 ), .Q ( new_AGEMA_signal_5609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1122 ( .C ( clk ), .D ( new_AGEMA_signal_5610 ), .Q ( new_AGEMA_signal_5611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1124 ( .C ( clk ), .D ( new_AGEMA_signal_5612 ), .Q ( new_AGEMA_signal_5613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1126 ( .C ( clk ), .D ( new_AGEMA_signal_5614 ), .Q ( new_AGEMA_signal_5615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1128 ( .C ( clk ), .D ( new_AGEMA_signal_5616 ), .Q ( new_AGEMA_signal_5617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1130 ( .C ( clk ), .D ( new_AGEMA_signal_5618 ), .Q ( new_AGEMA_signal_5619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1132 ( .C ( clk ), .D ( new_AGEMA_signal_5620 ), .Q ( new_AGEMA_signal_5621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1134 ( .C ( clk ), .D ( new_AGEMA_signal_5622 ), .Q ( new_AGEMA_signal_5623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1136 ( .C ( clk ), .D ( new_AGEMA_signal_5624 ), .Q ( new_AGEMA_signal_5625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1138 ( .C ( clk ), .D ( new_AGEMA_signal_5626 ), .Q ( new_AGEMA_signal_5627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1140 ( .C ( clk ), .D ( new_AGEMA_signal_5628 ), .Q ( new_AGEMA_signal_5629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1142 ( .C ( clk ), .D ( new_AGEMA_signal_5630 ), .Q ( new_AGEMA_signal_5631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1144 ( .C ( clk ), .D ( new_AGEMA_signal_5632 ), .Q ( new_AGEMA_signal_5633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1146 ( .C ( clk ), .D ( new_AGEMA_signal_5634 ), .Q ( new_AGEMA_signal_5635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1148 ( .C ( clk ), .D ( new_AGEMA_signal_5636 ), .Q ( new_AGEMA_signal_5637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1150 ( .C ( clk ), .D ( new_AGEMA_signal_5638 ), .Q ( new_AGEMA_signal_5639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1152 ( .C ( clk ), .D ( new_AGEMA_signal_5640 ), .Q ( new_AGEMA_signal_5641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1154 ( .C ( clk ), .D ( new_AGEMA_signal_5642 ), .Q ( new_AGEMA_signal_5643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1156 ( .C ( clk ), .D ( new_AGEMA_signal_5644 ), .Q ( new_AGEMA_signal_5645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1158 ( .C ( clk ), .D ( new_AGEMA_signal_5646 ), .Q ( new_AGEMA_signal_5647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1160 ( .C ( clk ), .D ( new_AGEMA_signal_5648 ), .Q ( new_AGEMA_signal_5649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1162 ( .C ( clk ), .D ( new_AGEMA_signal_5650 ), .Q ( new_AGEMA_signal_5651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1164 ( .C ( clk ), .D ( new_AGEMA_signal_5652 ), .Q ( new_AGEMA_signal_5653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1166 ( .C ( clk ), .D ( new_AGEMA_signal_5654 ), .Q ( new_AGEMA_signal_5655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1168 ( .C ( clk ), .D ( new_AGEMA_signal_5656 ), .Q ( new_AGEMA_signal_5657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1170 ( .C ( clk ), .D ( new_AGEMA_signal_5658 ), .Q ( new_AGEMA_signal_5659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1172 ( .C ( clk ), .D ( new_AGEMA_signal_5660 ), .Q ( new_AGEMA_signal_5661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1174 ( .C ( clk ), .D ( new_AGEMA_signal_5662 ), .Q ( new_AGEMA_signal_5663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1176 ( .C ( clk ), .D ( new_AGEMA_signal_5664 ), .Q ( new_AGEMA_signal_5665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1178 ( .C ( clk ), .D ( new_AGEMA_signal_5666 ), .Q ( new_AGEMA_signal_5667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1180 ( .C ( clk ), .D ( new_AGEMA_signal_5668 ), .Q ( new_AGEMA_signal_5669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1182 ( .C ( clk ), .D ( new_AGEMA_signal_5670 ), .Q ( new_AGEMA_signal_5671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1184 ( .C ( clk ), .D ( new_AGEMA_signal_5672 ), .Q ( new_AGEMA_signal_5673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1186 ( .C ( clk ), .D ( new_AGEMA_signal_5674 ), .Q ( new_AGEMA_signal_5675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1188 ( .C ( clk ), .D ( new_AGEMA_signal_5676 ), .Q ( new_AGEMA_signal_5677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1190 ( .C ( clk ), .D ( new_AGEMA_signal_5678 ), .Q ( new_AGEMA_signal_5679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1192 ( .C ( clk ), .D ( new_AGEMA_signal_5680 ), .Q ( new_AGEMA_signal_5681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1194 ( .C ( clk ), .D ( new_AGEMA_signal_5682 ), .Q ( new_AGEMA_signal_5683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1196 ( .C ( clk ), .D ( new_AGEMA_signal_5684 ), .Q ( new_AGEMA_signal_5685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1198 ( .C ( clk ), .D ( new_AGEMA_signal_5686 ), .Q ( new_AGEMA_signal_5687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1200 ( .C ( clk ), .D ( new_AGEMA_signal_5688 ), .Q ( new_AGEMA_signal_5689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1202 ( .C ( clk ), .D ( new_AGEMA_signal_5690 ), .Q ( new_AGEMA_signal_5691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1204 ( .C ( clk ), .D ( new_AGEMA_signal_5692 ), .Q ( new_AGEMA_signal_5693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1206 ( .C ( clk ), .D ( new_AGEMA_signal_5694 ), .Q ( new_AGEMA_signal_5695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1208 ( .C ( clk ), .D ( new_AGEMA_signal_5696 ), .Q ( new_AGEMA_signal_5697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1210 ( .C ( clk ), .D ( new_AGEMA_signal_5698 ), .Q ( new_AGEMA_signal_5699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1212 ( .C ( clk ), .D ( new_AGEMA_signal_5700 ), .Q ( new_AGEMA_signal_5701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1214 ( .C ( clk ), .D ( new_AGEMA_signal_5702 ), .Q ( new_AGEMA_signal_5703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1216 ( .C ( clk ), .D ( new_AGEMA_signal_5704 ), .Q ( new_AGEMA_signal_5705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1218 ( .C ( clk ), .D ( new_AGEMA_signal_5706 ), .Q ( new_AGEMA_signal_5707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1220 ( .C ( clk ), .D ( new_AGEMA_signal_5708 ), .Q ( new_AGEMA_signal_5709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1222 ( .C ( clk ), .D ( new_AGEMA_signal_5710 ), .Q ( new_AGEMA_signal_5711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1224 ( .C ( clk ), .D ( new_AGEMA_signal_5712 ), .Q ( new_AGEMA_signal_5713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1226 ( .C ( clk ), .D ( new_AGEMA_signal_5714 ), .Q ( new_AGEMA_signal_5715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1228 ( .C ( clk ), .D ( new_AGEMA_signal_5716 ), .Q ( new_AGEMA_signal_5717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1230 ( .C ( clk ), .D ( new_AGEMA_signal_5718 ), .Q ( new_AGEMA_signal_5719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1232 ( .C ( clk ), .D ( new_AGEMA_signal_5720 ), .Q ( new_AGEMA_signal_5721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1234 ( .C ( clk ), .D ( new_AGEMA_signal_5722 ), .Q ( new_AGEMA_signal_5723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1236 ( .C ( clk ), .D ( new_AGEMA_signal_5724 ), .Q ( new_AGEMA_signal_5725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1238 ( .C ( clk ), .D ( new_AGEMA_signal_5726 ), .Q ( new_AGEMA_signal_5727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1240 ( .C ( clk ), .D ( new_AGEMA_signal_5728 ), .Q ( new_AGEMA_signal_5729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1242 ( .C ( clk ), .D ( new_AGEMA_signal_5730 ), .Q ( new_AGEMA_signal_5731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1244 ( .C ( clk ), .D ( new_AGEMA_signal_5732 ), .Q ( new_AGEMA_signal_5733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1246 ( .C ( clk ), .D ( new_AGEMA_signal_5734 ), .Q ( new_AGEMA_signal_5735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1248 ( .C ( clk ), .D ( new_AGEMA_signal_5736 ), .Q ( new_AGEMA_signal_5737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1250 ( .C ( clk ), .D ( new_AGEMA_signal_5738 ), .Q ( new_AGEMA_signal_5739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1252 ( .C ( clk ), .D ( new_AGEMA_signal_5740 ), .Q ( new_AGEMA_signal_5741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1254 ( .C ( clk ), .D ( new_AGEMA_signal_5742 ), .Q ( new_AGEMA_signal_5743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C ( clk ), .D ( new_AGEMA_signal_5744 ), .Q ( new_AGEMA_signal_5745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C ( clk ), .D ( new_AGEMA_signal_5746 ), .Q ( new_AGEMA_signal_5747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C ( clk ), .D ( new_AGEMA_signal_5748 ), .Q ( new_AGEMA_signal_5749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C ( clk ), .D ( new_AGEMA_signal_5750 ), .Q ( new_AGEMA_signal_5751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C ( clk ), .D ( new_AGEMA_signal_5752 ), .Q ( new_AGEMA_signal_5753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C ( clk ), .D ( new_AGEMA_signal_5754 ), .Q ( new_AGEMA_signal_5755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C ( clk ), .D ( new_AGEMA_signal_5756 ), .Q ( new_AGEMA_signal_5757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C ( clk ), .D ( new_AGEMA_signal_5758 ), .Q ( new_AGEMA_signal_5759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C ( clk ), .D ( new_AGEMA_signal_5760 ), .Q ( new_AGEMA_signal_5761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C ( clk ), .D ( new_AGEMA_signal_5762 ), .Q ( new_AGEMA_signal_5763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C ( clk ), .D ( new_AGEMA_signal_5764 ), .Q ( new_AGEMA_signal_5765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C ( clk ), .D ( new_AGEMA_signal_5766 ), .Q ( new_AGEMA_signal_5767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C ( clk ), .D ( new_AGEMA_signal_5768 ), .Q ( new_AGEMA_signal_5769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C ( clk ), .D ( new_AGEMA_signal_5770 ), .Q ( new_AGEMA_signal_5771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C ( clk ), .D ( new_AGEMA_signal_5772 ), .Q ( new_AGEMA_signal_5773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C ( clk ), .D ( new_AGEMA_signal_5774 ), .Q ( new_AGEMA_signal_5775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C ( clk ), .D ( new_AGEMA_signal_5776 ), .Q ( new_AGEMA_signal_5777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C ( clk ), .D ( new_AGEMA_signal_5778 ), .Q ( new_AGEMA_signal_5779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C ( clk ), .D ( new_AGEMA_signal_5780 ), .Q ( new_AGEMA_signal_5781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C ( clk ), .D ( new_AGEMA_signal_5782 ), .Q ( new_AGEMA_signal_5783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C ( clk ), .D ( new_AGEMA_signal_5784 ), .Q ( new_AGEMA_signal_5785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C ( clk ), .D ( new_AGEMA_signal_5786 ), .Q ( new_AGEMA_signal_5787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C ( clk ), .D ( new_AGEMA_signal_5788 ), .Q ( new_AGEMA_signal_5789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C ( clk ), .D ( new_AGEMA_signal_5790 ), .Q ( new_AGEMA_signal_5791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C ( clk ), .D ( new_AGEMA_signal_5792 ), .Q ( new_AGEMA_signal_5793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C ( clk ), .D ( new_AGEMA_signal_5794 ), .Q ( new_AGEMA_signal_5795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C ( clk ), .D ( new_AGEMA_signal_5796 ), .Q ( new_AGEMA_signal_5797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C ( clk ), .D ( new_AGEMA_signal_5798 ), .Q ( new_AGEMA_signal_5799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C ( clk ), .D ( new_AGEMA_signal_5800 ), .Q ( new_AGEMA_signal_5801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C ( clk ), .D ( new_AGEMA_signal_5802 ), .Q ( new_AGEMA_signal_5803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C ( clk ), .D ( new_AGEMA_signal_5804 ), .Q ( new_AGEMA_signal_5805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C ( clk ), .D ( new_AGEMA_signal_5806 ), .Q ( new_AGEMA_signal_5807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C ( clk ), .D ( new_AGEMA_signal_5808 ), .Q ( new_AGEMA_signal_5809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1322 ( .C ( clk ), .D ( new_AGEMA_signal_5810 ), .Q ( new_AGEMA_signal_5811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C ( clk ), .D ( new_AGEMA_signal_5812 ), .Q ( new_AGEMA_signal_5813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C ( clk ), .D ( new_AGEMA_signal_5814 ), .Q ( new_AGEMA_signal_5815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C ( clk ), .D ( new_AGEMA_signal_5816 ), .Q ( new_AGEMA_signal_5817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C ( clk ), .D ( new_AGEMA_signal_5818 ), .Q ( new_AGEMA_signal_5819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C ( clk ), .D ( new_AGEMA_signal_5820 ), .Q ( new_AGEMA_signal_5821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C ( clk ), .D ( new_AGEMA_signal_5822 ), .Q ( new_AGEMA_signal_5823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C ( clk ), .D ( new_AGEMA_signal_5824 ), .Q ( new_AGEMA_signal_5825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C ( clk ), .D ( new_AGEMA_signal_5826 ), .Q ( new_AGEMA_signal_5827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C ( clk ), .D ( new_AGEMA_signal_5828 ), .Q ( new_AGEMA_signal_5829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C ( clk ), .D ( new_AGEMA_signal_5830 ), .Q ( new_AGEMA_signal_5831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C ( clk ), .D ( new_AGEMA_signal_5832 ), .Q ( new_AGEMA_signal_5833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C ( clk ), .D ( new_AGEMA_signal_5834 ), .Q ( new_AGEMA_signal_5835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C ( clk ), .D ( new_AGEMA_signal_5836 ), .Q ( new_AGEMA_signal_5837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C ( clk ), .D ( new_AGEMA_signal_5838 ), .Q ( new_AGEMA_signal_5839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C ( clk ), .D ( new_AGEMA_signal_5840 ), .Q ( new_AGEMA_signal_5841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C ( clk ), .D ( new_AGEMA_signal_5842 ), .Q ( new_AGEMA_signal_5843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C ( clk ), .D ( new_AGEMA_signal_5844 ), .Q ( new_AGEMA_signal_5845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C ( clk ), .D ( new_AGEMA_signal_5846 ), .Q ( new_AGEMA_signal_5847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1360 ( .C ( clk ), .D ( new_AGEMA_signal_5848 ), .Q ( new_AGEMA_signal_5849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1362 ( .C ( clk ), .D ( new_AGEMA_signal_5850 ), .Q ( new_AGEMA_signal_5851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1364 ( .C ( clk ), .D ( new_AGEMA_signal_5852 ), .Q ( new_AGEMA_signal_5853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1366 ( .C ( clk ), .D ( new_AGEMA_signal_5854 ), .Q ( new_AGEMA_signal_5855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1368 ( .C ( clk ), .D ( new_AGEMA_signal_5856 ), .Q ( new_AGEMA_signal_5857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1370 ( .C ( clk ), .D ( new_AGEMA_signal_5858 ), .Q ( new_AGEMA_signal_5859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1372 ( .C ( clk ), .D ( new_AGEMA_signal_5860 ), .Q ( new_AGEMA_signal_5861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1374 ( .C ( clk ), .D ( new_AGEMA_signal_5862 ), .Q ( new_AGEMA_signal_5863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1376 ( .C ( clk ), .D ( new_AGEMA_signal_5864 ), .Q ( new_AGEMA_signal_5865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1378 ( .C ( clk ), .D ( new_AGEMA_signal_5866 ), .Q ( new_AGEMA_signal_5867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1380 ( .C ( clk ), .D ( new_AGEMA_signal_5868 ), .Q ( new_AGEMA_signal_5869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1382 ( .C ( clk ), .D ( new_AGEMA_signal_5870 ), .Q ( new_AGEMA_signal_5871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1384 ( .C ( clk ), .D ( new_AGEMA_signal_5872 ), .Q ( new_AGEMA_signal_5873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1386 ( .C ( clk ), .D ( new_AGEMA_signal_5874 ), .Q ( new_AGEMA_signal_5875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1388 ( .C ( clk ), .D ( new_AGEMA_signal_5876 ), .Q ( new_AGEMA_signal_5877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1390 ( .C ( clk ), .D ( new_AGEMA_signal_5878 ), .Q ( new_AGEMA_signal_5879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1392 ( .C ( clk ), .D ( new_AGEMA_signal_5880 ), .Q ( new_AGEMA_signal_5881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1394 ( .C ( clk ), .D ( new_AGEMA_signal_5882 ), .Q ( new_AGEMA_signal_5883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1396 ( .C ( clk ), .D ( new_AGEMA_signal_5884 ), .Q ( new_AGEMA_signal_5885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1398 ( .C ( clk ), .D ( new_AGEMA_signal_5886 ), .Q ( new_AGEMA_signal_5887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1400 ( .C ( clk ), .D ( new_AGEMA_signal_5888 ), .Q ( new_AGEMA_signal_5889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1402 ( .C ( clk ), .D ( new_AGEMA_signal_5890 ), .Q ( new_AGEMA_signal_5891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1404 ( .C ( clk ), .D ( new_AGEMA_signal_5892 ), .Q ( new_AGEMA_signal_5893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1406 ( .C ( clk ), .D ( new_AGEMA_signal_5894 ), .Q ( new_AGEMA_signal_5895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1408 ( .C ( clk ), .D ( new_AGEMA_signal_5896 ), .Q ( new_AGEMA_signal_5897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1410 ( .C ( clk ), .D ( new_AGEMA_signal_5898 ), .Q ( new_AGEMA_signal_5899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1412 ( .C ( clk ), .D ( new_AGEMA_signal_5900 ), .Q ( new_AGEMA_signal_5901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1414 ( .C ( clk ), .D ( new_AGEMA_signal_5902 ), .Q ( new_AGEMA_signal_5903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1416 ( .C ( clk ), .D ( new_AGEMA_signal_5904 ), .Q ( new_AGEMA_signal_5905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1418 ( .C ( clk ), .D ( new_AGEMA_signal_5906 ), .Q ( new_AGEMA_signal_5907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1420 ( .C ( clk ), .D ( new_AGEMA_signal_5908 ), .Q ( new_AGEMA_signal_5909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1422 ( .C ( clk ), .D ( new_AGEMA_signal_5910 ), .Q ( new_AGEMA_signal_5911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1424 ( .C ( clk ), .D ( new_AGEMA_signal_5912 ), .Q ( new_AGEMA_signal_5913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1438 ( .C ( clk ), .D ( new_AGEMA_signal_5926 ), .Q ( new_AGEMA_signal_5927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1442 ( .C ( clk ), .D ( new_AGEMA_signal_5930 ), .Q ( new_AGEMA_signal_5931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1446 ( .C ( clk ), .D ( new_AGEMA_signal_5934 ), .Q ( new_AGEMA_signal_5935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1516 ( .C ( clk ), .D ( new_AGEMA_signal_6004 ), .Q ( new_AGEMA_signal_6005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1520 ( .C ( clk ), .D ( new_AGEMA_signal_6008 ), .Q ( new_AGEMA_signal_6009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1524 ( .C ( clk ), .D ( new_AGEMA_signal_6012 ), .Q ( new_AGEMA_signal_6013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1570 ( .C ( clk ), .D ( new_AGEMA_signal_6058 ), .Q ( new_AGEMA_signal_6059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1574 ( .C ( clk ), .D ( new_AGEMA_signal_6062 ), .Q ( new_AGEMA_signal_6063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1578 ( .C ( clk ), .D ( new_AGEMA_signal_6066 ), .Q ( new_AGEMA_signal_6067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1612 ( .C ( clk ), .D ( new_AGEMA_signal_6100 ), .Q ( new_AGEMA_signal_6101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1616 ( .C ( clk ), .D ( new_AGEMA_signal_6104 ), .Q ( new_AGEMA_signal_6105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1620 ( .C ( clk ), .D ( new_AGEMA_signal_6108 ), .Q ( new_AGEMA_signal_6109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1642 ( .C ( clk ), .D ( new_AGEMA_signal_6130 ), .Q ( new_AGEMA_signal_6131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1646 ( .C ( clk ), .D ( new_AGEMA_signal_6134 ), .Q ( new_AGEMA_signal_6135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1650 ( .C ( clk ), .D ( new_AGEMA_signal_6138 ), .Q ( new_AGEMA_signal_6139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1672 ( .C ( clk ), .D ( new_AGEMA_signal_6160 ), .Q ( new_AGEMA_signal_6161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1676 ( .C ( clk ), .D ( new_AGEMA_signal_6164 ), .Q ( new_AGEMA_signal_6165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1680 ( .C ( clk ), .D ( new_AGEMA_signal_6168 ), .Q ( new_AGEMA_signal_6169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C ( clk ), .D ( new_AGEMA_signal_6276 ), .Q ( new_AGEMA_signal_6277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C ( clk ), .D ( new_AGEMA_signal_6282 ), .Q ( new_AGEMA_signal_6283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C ( clk ), .D ( new_AGEMA_signal_6288 ), .Q ( new_AGEMA_signal_6289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C ( clk ), .D ( new_AGEMA_signal_6310 ), .Q ( new_AGEMA_signal_6311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C ( clk ), .D ( new_AGEMA_signal_6314 ), .Q ( new_AGEMA_signal_6315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C ( clk ), .D ( new_AGEMA_signal_6318 ), .Q ( new_AGEMA_signal_6319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C ( clk ), .D ( new_AGEMA_signal_6340 ), .Q ( new_AGEMA_signal_6341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C ( clk ), .D ( new_AGEMA_signal_6344 ), .Q ( new_AGEMA_signal_6345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C ( clk ), .D ( new_AGEMA_signal_6348 ), .Q ( new_AGEMA_signal_6349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C ( clk ), .D ( new_AGEMA_signal_6394 ), .Q ( new_AGEMA_signal_6395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C ( clk ), .D ( new_AGEMA_signal_6398 ), .Q ( new_AGEMA_signal_6399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C ( clk ), .D ( new_AGEMA_signal_6402 ), .Q ( new_AGEMA_signal_6403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C ( clk ), .D ( new_AGEMA_signal_6418 ), .Q ( new_AGEMA_signal_6419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C ( clk ), .D ( new_AGEMA_signal_6422 ), .Q ( new_AGEMA_signal_6423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C ( clk ), .D ( new_AGEMA_signal_6426 ), .Q ( new_AGEMA_signal_6427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2152 ( .C ( clk ), .D ( new_AGEMA_signal_6640 ), .Q ( new_AGEMA_signal_6641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C ( clk ), .D ( new_AGEMA_signal_6646 ), .Q ( new_AGEMA_signal_6647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2164 ( .C ( clk ), .D ( new_AGEMA_signal_6652 ), .Q ( new_AGEMA_signal_6653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2230 ( .C ( clk ), .D ( new_AGEMA_signal_6718 ), .Q ( new_AGEMA_signal_6719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2236 ( .C ( clk ), .D ( new_AGEMA_signal_6724 ), .Q ( new_AGEMA_signal_6725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2242 ( .C ( clk ), .D ( new_AGEMA_signal_6730 ), .Q ( new_AGEMA_signal_6731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2578 ( .C ( clk ), .D ( new_AGEMA_signal_7066 ), .Q ( new_AGEMA_signal_7067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2586 ( .C ( clk ), .D ( new_AGEMA_signal_7074 ), .Q ( new_AGEMA_signal_7075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2594 ( .C ( clk ), .D ( new_AGEMA_signal_7082 ), .Q ( new_AGEMA_signal_7083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2608 ( .C ( clk ), .D ( new_AGEMA_signal_7096 ), .Q ( new_AGEMA_signal_7097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2616 ( .C ( clk ), .D ( new_AGEMA_signal_7104 ), .Q ( new_AGEMA_signal_7105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2624 ( .C ( clk ), .D ( new_AGEMA_signal_7112 ), .Q ( new_AGEMA_signal_7113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2836 ( .C ( clk ), .D ( new_AGEMA_signal_7324 ), .Q ( new_AGEMA_signal_7325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2844 ( .C ( clk ), .D ( new_AGEMA_signal_7332 ), .Q ( new_AGEMA_signal_7333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2852 ( .C ( clk ), .D ( new_AGEMA_signal_7340 ), .Q ( new_AGEMA_signal_7341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3094 ( .C ( clk ), .D ( new_AGEMA_signal_7582 ), .Q ( new_AGEMA_signal_7583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3102 ( .C ( clk ), .D ( new_AGEMA_signal_7590 ), .Q ( new_AGEMA_signal_7591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3110 ( .C ( clk ), .D ( new_AGEMA_signal_7598 ), .Q ( new_AGEMA_signal_7599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3184 ( .C ( clk ), .D ( new_AGEMA_signal_7672 ), .Q ( new_AGEMA_signal_7673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3192 ( .C ( clk ), .D ( new_AGEMA_signal_7680 ), .Q ( new_AGEMA_signal_7681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3200 ( .C ( clk ), .D ( new_AGEMA_signal_7688 ), .Q ( new_AGEMA_signal_7689 ) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_1425 ( .C ( clk ), .D ( n2755 ), .Q ( new_AGEMA_signal_5914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1427 ( .C ( clk ), .D ( new_AGEMA_signal_1118 ), .Q ( new_AGEMA_signal_5916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1429 ( .C ( clk ), .D ( new_AGEMA_signal_1119 ), .Q ( new_AGEMA_signal_5918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1431 ( .C ( clk ), .D ( n2151 ), .Q ( new_AGEMA_signal_5920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1433 ( .C ( clk ), .D ( new_AGEMA_signal_1322 ), .Q ( new_AGEMA_signal_5922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1435 ( .C ( clk ), .D ( new_AGEMA_signal_1323 ), .Q ( new_AGEMA_signal_5924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1439 ( .C ( clk ), .D ( new_AGEMA_signal_5927 ), .Q ( new_AGEMA_signal_5928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1443 ( .C ( clk ), .D ( new_AGEMA_signal_5931 ), .Q ( new_AGEMA_signal_5932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1447 ( .C ( clk ), .D ( new_AGEMA_signal_5935 ), .Q ( new_AGEMA_signal_5936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1449 ( .C ( clk ), .D ( new_AGEMA_signal_5555 ), .Q ( new_AGEMA_signal_5938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1451 ( .C ( clk ), .D ( new_AGEMA_signal_5557 ), .Q ( new_AGEMA_signal_5940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1453 ( .C ( clk ), .D ( new_AGEMA_signal_5559 ), .Q ( new_AGEMA_signal_5942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1455 ( .C ( clk ), .D ( new_AGEMA_signal_5537 ), .Q ( new_AGEMA_signal_5944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1457 ( .C ( clk ), .D ( new_AGEMA_signal_5539 ), .Q ( new_AGEMA_signal_5946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1459 ( .C ( clk ), .D ( new_AGEMA_signal_5541 ), .Q ( new_AGEMA_signal_5948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1461 ( .C ( clk ), .D ( n1964 ), .Q ( new_AGEMA_signal_5950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1463 ( .C ( clk ), .D ( new_AGEMA_signal_1056 ), .Q ( new_AGEMA_signal_5952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1465 ( .C ( clk ), .D ( new_AGEMA_signal_1057 ), .Q ( new_AGEMA_signal_5954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1467 ( .C ( clk ), .D ( n2673 ), .Q ( new_AGEMA_signal_5956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1469 ( .C ( clk ), .D ( new_AGEMA_signal_1162 ), .Q ( new_AGEMA_signal_5958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1471 ( .C ( clk ), .D ( new_AGEMA_signal_1163 ), .Q ( new_AGEMA_signal_5960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1473 ( .C ( clk ), .D ( n2359 ), .Q ( new_AGEMA_signal_5962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1475 ( .C ( clk ), .D ( new_AGEMA_signal_1352 ), .Q ( new_AGEMA_signal_5964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1477 ( .C ( clk ), .D ( new_AGEMA_signal_1353 ), .Q ( new_AGEMA_signal_5966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1479 ( .C ( clk ), .D ( n1973 ), .Q ( new_AGEMA_signal_5968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1481 ( .C ( clk ), .D ( new_AGEMA_signal_1360 ), .Q ( new_AGEMA_signal_5970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1483 ( .C ( clk ), .D ( new_AGEMA_signal_1361 ), .Q ( new_AGEMA_signal_5972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1485 ( .C ( clk ), .D ( n2690 ), .Q ( new_AGEMA_signal_5974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1487 ( .C ( clk ), .D ( new_AGEMA_signal_1180 ), .Q ( new_AGEMA_signal_5976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1489 ( .C ( clk ), .D ( new_AGEMA_signal_1181 ), .Q ( new_AGEMA_signal_5978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1491 ( .C ( clk ), .D ( n2741 ), .Q ( new_AGEMA_signal_5980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1493 ( .C ( clk ), .D ( new_AGEMA_signal_1364 ), .Q ( new_AGEMA_signal_5982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1495 ( .C ( clk ), .D ( new_AGEMA_signal_1365 ), .Q ( new_AGEMA_signal_5984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1497 ( .C ( clk ), .D ( n1993 ), .Q ( new_AGEMA_signal_5986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1499 ( .C ( clk ), .D ( new_AGEMA_signal_1186 ), .Q ( new_AGEMA_signal_5988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1501 ( .C ( clk ), .D ( new_AGEMA_signal_1187 ), .Q ( new_AGEMA_signal_5990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1503 ( .C ( clk ), .D ( n2241 ), .Q ( new_AGEMA_signal_5992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1505 ( .C ( clk ), .D ( new_AGEMA_signal_1372 ), .Q ( new_AGEMA_signal_5994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1507 ( .C ( clk ), .D ( new_AGEMA_signal_1373 ), .Q ( new_AGEMA_signal_5996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1509 ( .C ( clk ), .D ( new_AGEMA_signal_5717 ), .Q ( new_AGEMA_signal_5998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1511 ( .C ( clk ), .D ( new_AGEMA_signal_5719 ), .Q ( new_AGEMA_signal_6000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1513 ( .C ( clk ), .D ( new_AGEMA_signal_5721 ), .Q ( new_AGEMA_signal_6002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1517 ( .C ( clk ), .D ( new_AGEMA_signal_6005 ), .Q ( new_AGEMA_signal_6006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1521 ( .C ( clk ), .D ( new_AGEMA_signal_6009 ), .Q ( new_AGEMA_signal_6010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1525 ( .C ( clk ), .D ( new_AGEMA_signal_6013 ), .Q ( new_AGEMA_signal_6014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1527 ( .C ( clk ), .D ( n2290 ), .Q ( new_AGEMA_signal_6016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1529 ( .C ( clk ), .D ( new_AGEMA_signal_1394 ), .Q ( new_AGEMA_signal_6018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1531 ( .C ( clk ), .D ( new_AGEMA_signal_1395 ), .Q ( new_AGEMA_signal_6020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1533 ( .C ( clk ), .D ( n2171 ), .Q ( new_AGEMA_signal_6022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1535 ( .C ( clk ), .D ( new_AGEMA_signal_1204 ), .Q ( new_AGEMA_signal_6024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1537 ( .C ( clk ), .D ( new_AGEMA_signal_1205 ), .Q ( new_AGEMA_signal_6026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1539 ( .C ( clk ), .D ( n2042 ), .Q ( new_AGEMA_signal_6028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1541 ( .C ( clk ), .D ( new_AGEMA_signal_1402 ), .Q ( new_AGEMA_signal_6030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1543 ( .C ( clk ), .D ( new_AGEMA_signal_1403 ), .Q ( new_AGEMA_signal_6032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1545 ( .C ( clk ), .D ( n2754 ), .Q ( new_AGEMA_signal_6034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1547 ( .C ( clk ), .D ( new_AGEMA_signal_1404 ), .Q ( new_AGEMA_signal_6036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1549 ( .C ( clk ), .D ( new_AGEMA_signal_1405 ), .Q ( new_AGEMA_signal_6038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1551 ( .C ( clk ), .D ( new_AGEMA_signal_5507 ), .Q ( new_AGEMA_signal_6040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1553 ( .C ( clk ), .D ( new_AGEMA_signal_5509 ), .Q ( new_AGEMA_signal_6042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1555 ( .C ( clk ), .D ( new_AGEMA_signal_5511 ), .Q ( new_AGEMA_signal_6044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1557 ( .C ( clk ), .D ( n2535 ), .Q ( new_AGEMA_signal_6046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1559 ( .C ( clk ), .D ( new_AGEMA_signal_1358 ), .Q ( new_AGEMA_signal_6048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1561 ( .C ( clk ), .D ( new_AGEMA_signal_1359 ), .Q ( new_AGEMA_signal_6050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1563 ( .C ( clk ), .D ( n2642 ), .Q ( new_AGEMA_signal_6052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1565 ( .C ( clk ), .D ( new_AGEMA_signal_1206 ), .Q ( new_AGEMA_signal_6054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1567 ( .C ( clk ), .D ( new_AGEMA_signal_1207 ), .Q ( new_AGEMA_signal_6056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1571 ( .C ( clk ), .D ( new_AGEMA_signal_6059 ), .Q ( new_AGEMA_signal_6060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1575 ( .C ( clk ), .D ( new_AGEMA_signal_6063 ), .Q ( new_AGEMA_signal_6064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1579 ( .C ( clk ), .D ( new_AGEMA_signal_6067 ), .Q ( new_AGEMA_signal_6068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1581 ( .C ( clk ), .D ( n2773 ), .Q ( new_AGEMA_signal_6070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1583 ( .C ( clk ), .D ( new_AGEMA_signal_1426 ), .Q ( new_AGEMA_signal_6072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1585 ( .C ( clk ), .D ( new_AGEMA_signal_1427 ), .Q ( new_AGEMA_signal_6074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1587 ( .C ( clk ), .D ( n2627 ), .Q ( new_AGEMA_signal_6076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1589 ( .C ( clk ), .D ( new_AGEMA_signal_1154 ), .Q ( new_AGEMA_signal_6078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1591 ( .C ( clk ), .D ( new_AGEMA_signal_1155 ), .Q ( new_AGEMA_signal_6080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1593 ( .C ( clk ), .D ( new_AGEMA_signal_5627 ), .Q ( new_AGEMA_signal_6082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1595 ( .C ( clk ), .D ( new_AGEMA_signal_5629 ), .Q ( new_AGEMA_signal_6084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1597 ( .C ( clk ), .D ( new_AGEMA_signal_5631 ), .Q ( new_AGEMA_signal_6086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1599 ( .C ( clk ), .D ( n2631 ), .Q ( new_AGEMA_signal_6088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1601 ( .C ( clk ), .D ( new_AGEMA_signal_1126 ), .Q ( new_AGEMA_signal_6090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1603 ( .C ( clk ), .D ( new_AGEMA_signal_1127 ), .Q ( new_AGEMA_signal_6092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1605 ( .C ( clk ), .D ( n2376 ), .Q ( new_AGEMA_signal_6094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1607 ( .C ( clk ), .D ( new_AGEMA_signal_1396 ), .Q ( new_AGEMA_signal_6096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1609 ( .C ( clk ), .D ( new_AGEMA_signal_1397 ), .Q ( new_AGEMA_signal_6098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1613 ( .C ( clk ), .D ( new_AGEMA_signal_6101 ), .Q ( new_AGEMA_signal_6102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1617 ( .C ( clk ), .D ( new_AGEMA_signal_6105 ), .Q ( new_AGEMA_signal_6106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1621 ( .C ( clk ), .D ( new_AGEMA_signal_6109 ), .Q ( new_AGEMA_signal_6110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1623 ( .C ( clk ), .D ( new_AGEMA_signal_5765 ), .Q ( new_AGEMA_signal_6112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1625 ( .C ( clk ), .D ( new_AGEMA_signal_5767 ), .Q ( new_AGEMA_signal_6114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1627 ( .C ( clk ), .D ( new_AGEMA_signal_5769 ), .Q ( new_AGEMA_signal_6116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1629 ( .C ( clk ), .D ( new_AGEMA_signal_5657 ), .Q ( new_AGEMA_signal_6118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1631 ( .C ( clk ), .D ( new_AGEMA_signal_5659 ), .Q ( new_AGEMA_signal_6120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1633 ( .C ( clk ), .D ( new_AGEMA_signal_5661 ), .Q ( new_AGEMA_signal_6122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1635 ( .C ( clk ), .D ( new_AGEMA_signal_5681 ), .Q ( new_AGEMA_signal_6124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1637 ( .C ( clk ), .D ( new_AGEMA_signal_5683 ), .Q ( new_AGEMA_signal_6126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1639 ( .C ( clk ), .D ( new_AGEMA_signal_5685 ), .Q ( new_AGEMA_signal_6128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1643 ( .C ( clk ), .D ( new_AGEMA_signal_6131 ), .Q ( new_AGEMA_signal_6132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1647 ( .C ( clk ), .D ( new_AGEMA_signal_6135 ), .Q ( new_AGEMA_signal_6136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1651 ( .C ( clk ), .D ( new_AGEMA_signal_6139 ), .Q ( new_AGEMA_signal_6140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1653 ( .C ( clk ), .D ( new_AGEMA_signal_5885 ), .Q ( new_AGEMA_signal_6142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1655 ( .C ( clk ), .D ( new_AGEMA_signal_5887 ), .Q ( new_AGEMA_signal_6144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1657 ( .C ( clk ), .D ( new_AGEMA_signal_5889 ), .Q ( new_AGEMA_signal_6146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1659 ( .C ( clk ), .D ( n2498 ), .Q ( new_AGEMA_signal_6148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1661 ( .C ( clk ), .D ( new_AGEMA_signal_1212 ), .Q ( new_AGEMA_signal_6150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1663 ( .C ( clk ), .D ( new_AGEMA_signal_1213 ), .Q ( new_AGEMA_signal_6152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1665 ( .C ( clk ), .D ( n2178 ), .Q ( new_AGEMA_signal_6154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1667 ( .C ( clk ), .D ( new_AGEMA_signal_1228 ), .Q ( new_AGEMA_signal_6156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1669 ( .C ( clk ), .D ( new_AGEMA_signal_1229 ), .Q ( new_AGEMA_signal_6158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1673 ( .C ( clk ), .D ( new_AGEMA_signal_6161 ), .Q ( new_AGEMA_signal_6162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1677 ( .C ( clk ), .D ( new_AGEMA_signal_6165 ), .Q ( new_AGEMA_signal_6166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1681 ( .C ( clk ), .D ( new_AGEMA_signal_6169 ), .Q ( new_AGEMA_signal_6170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1683 ( .C ( clk ), .D ( n2505 ), .Q ( new_AGEMA_signal_6172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1685 ( .C ( clk ), .D ( new_AGEMA_signal_1350 ), .Q ( new_AGEMA_signal_6174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1687 ( .C ( clk ), .D ( new_AGEMA_signal_1351 ), .Q ( new_AGEMA_signal_6176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1689 ( .C ( clk ), .D ( n2540 ), .Q ( new_AGEMA_signal_6178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1691 ( .C ( clk ), .D ( new_AGEMA_signal_1500 ), .Q ( new_AGEMA_signal_6180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1693 ( .C ( clk ), .D ( new_AGEMA_signal_1501 ), .Q ( new_AGEMA_signal_6182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1695 ( .C ( clk ), .D ( n2266 ), .Q ( new_AGEMA_signal_6184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1697 ( .C ( clk ), .D ( new_AGEMA_signal_1242 ), .Q ( new_AGEMA_signal_6186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1699 ( .C ( clk ), .D ( new_AGEMA_signal_1243 ), .Q ( new_AGEMA_signal_6188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1701 ( .C ( clk ), .D ( n2278 ), .Q ( new_AGEMA_signal_6190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1703 ( .C ( clk ), .D ( new_AGEMA_signal_1508 ), .Q ( new_AGEMA_signal_6192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1705 ( .C ( clk ), .D ( new_AGEMA_signal_1509 ), .Q ( new_AGEMA_signal_6194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1707 ( .C ( clk ), .D ( new_AGEMA_signal_5753 ), .Q ( new_AGEMA_signal_6196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1709 ( .C ( clk ), .D ( new_AGEMA_signal_5755 ), .Q ( new_AGEMA_signal_6198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1711 ( .C ( clk ), .D ( new_AGEMA_signal_5757 ), .Q ( new_AGEMA_signal_6200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1713 ( .C ( clk ), .D ( new_AGEMA_signal_5819 ), .Q ( new_AGEMA_signal_6202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C ( clk ), .D ( new_AGEMA_signal_5821 ), .Q ( new_AGEMA_signal_6204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C ( clk ), .D ( new_AGEMA_signal_5823 ), .Q ( new_AGEMA_signal_6206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C ( clk ), .D ( new_AGEMA_signal_5615 ), .Q ( new_AGEMA_signal_6208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C ( clk ), .D ( new_AGEMA_signal_5617 ), .Q ( new_AGEMA_signal_6210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C ( clk ), .D ( new_AGEMA_signal_5619 ), .Q ( new_AGEMA_signal_6212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C ( clk ), .D ( new_AGEMA_signal_5603 ), .Q ( new_AGEMA_signal_6214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C ( clk ), .D ( new_AGEMA_signal_5605 ), .Q ( new_AGEMA_signal_6216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C ( clk ), .D ( new_AGEMA_signal_5607 ), .Q ( new_AGEMA_signal_6218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C ( clk ), .D ( n2318 ), .Q ( new_AGEMA_signal_6220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C ( clk ), .D ( new_AGEMA_signal_1254 ), .Q ( new_AGEMA_signal_6222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C ( clk ), .D ( new_AGEMA_signal_1255 ), .Q ( new_AGEMA_signal_6224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C ( clk ), .D ( n2325 ), .Q ( new_AGEMA_signal_6226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C ( clk ), .D ( new_AGEMA_signal_1528 ), .Q ( new_AGEMA_signal_6228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C ( clk ), .D ( new_AGEMA_signal_1529 ), .Q ( new_AGEMA_signal_6230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C ( clk ), .D ( n2677 ), .Q ( new_AGEMA_signal_6232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C ( clk ), .D ( new_AGEMA_signal_1152 ), .Q ( new_AGEMA_signal_6234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C ( clk ), .D ( new_AGEMA_signal_1153 ), .Q ( new_AGEMA_signal_6236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C ( clk ), .D ( new_AGEMA_signal_5873 ), .Q ( new_AGEMA_signal_6238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C ( clk ), .D ( new_AGEMA_signal_5875 ), .Q ( new_AGEMA_signal_6240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C ( clk ), .D ( new_AGEMA_signal_5877 ), .Q ( new_AGEMA_signal_6242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C ( clk ), .D ( new_AGEMA_signal_5897 ), .Q ( new_AGEMA_signal_6244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1757 ( .C ( clk ), .D ( new_AGEMA_signal_5899 ), .Q ( new_AGEMA_signal_6246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C ( clk ), .D ( new_AGEMA_signal_5901 ), .Q ( new_AGEMA_signal_6248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C ( clk ), .D ( new_AGEMA_signal_5669 ), .Q ( new_AGEMA_signal_6250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C ( clk ), .D ( new_AGEMA_signal_5671 ), .Q ( new_AGEMA_signal_6252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C ( clk ), .D ( new_AGEMA_signal_5673 ), .Q ( new_AGEMA_signal_6254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C ( clk ), .D ( new_AGEMA_signal_5519 ), .Q ( new_AGEMA_signal_6256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C ( clk ), .D ( new_AGEMA_signal_5521 ), .Q ( new_AGEMA_signal_6258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C ( clk ), .D ( new_AGEMA_signal_5523 ), .Q ( new_AGEMA_signal_6260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C ( clk ), .D ( n2625 ), .Q ( new_AGEMA_signal_6262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C ( clk ), .D ( new_AGEMA_signal_1354 ), .Q ( new_AGEMA_signal_6264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C ( clk ), .D ( new_AGEMA_signal_1355 ), .Q ( new_AGEMA_signal_6266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C ( clk ), .D ( n2431 ), .Q ( new_AGEMA_signal_6268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C ( clk ), .D ( new_AGEMA_signal_1570 ), .Q ( new_AGEMA_signal_6270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C ( clk ), .D ( new_AGEMA_signal_1571 ), .Q ( new_AGEMA_signal_6272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C ( clk ), .D ( new_AGEMA_signal_6277 ), .Q ( new_AGEMA_signal_6278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C ( clk ), .D ( new_AGEMA_signal_6283 ), .Q ( new_AGEMA_signal_6284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C ( clk ), .D ( new_AGEMA_signal_6289 ), .Q ( new_AGEMA_signal_6290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C ( clk ), .D ( n2453 ), .Q ( new_AGEMA_signal_6292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C ( clk ), .D ( new_AGEMA_signal_1274 ), .Q ( new_AGEMA_signal_6294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C ( clk ), .D ( new_AGEMA_signal_1275 ), .Q ( new_AGEMA_signal_6296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C ( clk ), .D ( n2475 ), .Q ( new_AGEMA_signal_6298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C ( clk ), .D ( new_AGEMA_signal_1284 ), .Q ( new_AGEMA_signal_6300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C ( clk ), .D ( new_AGEMA_signal_1285 ), .Q ( new_AGEMA_signal_6302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C ( clk ), .D ( n2487 ), .Q ( new_AGEMA_signal_6304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C ( clk ), .D ( new_AGEMA_signal_1586 ), .Q ( new_AGEMA_signal_6306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C ( clk ), .D ( new_AGEMA_signal_1587 ), .Q ( new_AGEMA_signal_6308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C ( clk ), .D ( new_AGEMA_signal_6311 ), .Q ( new_AGEMA_signal_6312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C ( clk ), .D ( new_AGEMA_signal_6315 ), .Q ( new_AGEMA_signal_6316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C ( clk ), .D ( new_AGEMA_signal_6319 ), .Q ( new_AGEMA_signal_6320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C ( clk ), .D ( new_AGEMA_signal_5729 ), .Q ( new_AGEMA_signal_6322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C ( clk ), .D ( new_AGEMA_signal_5731 ), .Q ( new_AGEMA_signal_6324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C ( clk ), .D ( new_AGEMA_signal_5733 ), .Q ( new_AGEMA_signal_6326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C ( clk ), .D ( new_AGEMA_signal_5741 ), .Q ( new_AGEMA_signal_6328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C ( clk ), .D ( new_AGEMA_signal_5743 ), .Q ( new_AGEMA_signal_6330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C ( clk ), .D ( new_AGEMA_signal_5745 ), .Q ( new_AGEMA_signal_6332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C ( clk ), .D ( n2564 ), .Q ( new_AGEMA_signal_6334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C ( clk ), .D ( new_AGEMA_signal_1608 ), .Q ( new_AGEMA_signal_6336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C ( clk ), .D ( new_AGEMA_signal_1609 ), .Q ( new_AGEMA_signal_6338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C ( clk ), .D ( new_AGEMA_signal_6341 ), .Q ( new_AGEMA_signal_6342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C ( clk ), .D ( new_AGEMA_signal_6345 ), .Q ( new_AGEMA_signal_6346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C ( clk ), .D ( new_AGEMA_signal_6349 ), .Q ( new_AGEMA_signal_6350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C ( clk ), .D ( n2617 ), .Q ( new_AGEMA_signal_6352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C ( clk ), .D ( new_AGEMA_signal_1296 ), .Q ( new_AGEMA_signal_6354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C ( clk ), .D ( new_AGEMA_signal_1297 ), .Q ( new_AGEMA_signal_6356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C ( clk ), .D ( n2647 ), .Q ( new_AGEMA_signal_6358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C ( clk ), .D ( new_AGEMA_signal_1220 ), .Q ( new_AGEMA_signal_6360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C ( clk ), .D ( new_AGEMA_signal_1221 ), .Q ( new_AGEMA_signal_6362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C ( clk ), .D ( n2674 ), .Q ( new_AGEMA_signal_6364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C ( clk ), .D ( new_AGEMA_signal_1808 ), .Q ( new_AGEMA_signal_6366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C ( clk ), .D ( new_AGEMA_signal_1809 ), .Q ( new_AGEMA_signal_6368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C ( clk ), .D ( n2683 ), .Q ( new_AGEMA_signal_6370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C ( clk ), .D ( new_AGEMA_signal_1102 ), .Q ( new_AGEMA_signal_6372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C ( clk ), .D ( new_AGEMA_signal_1103 ), .Q ( new_AGEMA_signal_6374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C ( clk ), .D ( n2714 ), .Q ( new_AGEMA_signal_6376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C ( clk ), .D ( new_AGEMA_signal_1302 ), .Q ( new_AGEMA_signal_6378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C ( clk ), .D ( new_AGEMA_signal_1303 ), .Q ( new_AGEMA_signal_6380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C ( clk ), .D ( n2726 ), .Q ( new_AGEMA_signal_6382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C ( clk ), .D ( new_AGEMA_signal_1652 ), .Q ( new_AGEMA_signal_6384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C ( clk ), .D ( new_AGEMA_signal_1653 ), .Q ( new_AGEMA_signal_6386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C ( clk ), .D ( n2734 ), .Q ( new_AGEMA_signal_6388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C ( clk ), .D ( new_AGEMA_signal_1324 ), .Q ( new_AGEMA_signal_6390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C ( clk ), .D ( new_AGEMA_signal_1325 ), .Q ( new_AGEMA_signal_6392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C ( clk ), .D ( new_AGEMA_signal_6395 ), .Q ( new_AGEMA_signal_6396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C ( clk ), .D ( new_AGEMA_signal_6399 ), .Q ( new_AGEMA_signal_6400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C ( clk ), .D ( new_AGEMA_signal_6403 ), .Q ( new_AGEMA_signal_6404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C ( clk ), .D ( n2763 ), .Q ( new_AGEMA_signal_6406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C ( clk ), .D ( new_AGEMA_signal_1326 ), .Q ( new_AGEMA_signal_6408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C ( clk ), .D ( new_AGEMA_signal_1327 ), .Q ( new_AGEMA_signal_6410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C ( clk ), .D ( n2784 ), .Q ( new_AGEMA_signal_6412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C ( clk ), .D ( new_AGEMA_signal_1632 ), .Q ( new_AGEMA_signal_6414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C ( clk ), .D ( new_AGEMA_signal_1633 ), .Q ( new_AGEMA_signal_6416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C ( clk ), .D ( new_AGEMA_signal_6419 ), .Q ( new_AGEMA_signal_6420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C ( clk ), .D ( new_AGEMA_signal_6423 ), .Q ( new_AGEMA_signal_6424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C ( clk ), .D ( new_AGEMA_signal_6427 ), .Q ( new_AGEMA_signal_6428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C ( clk ), .D ( n2820 ), .Q ( new_AGEMA_signal_6430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C ( clk ), .D ( new_AGEMA_signal_1310 ), .Q ( new_AGEMA_signal_6432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C ( clk ), .D ( new_AGEMA_signal_1311 ), .Q ( new_AGEMA_signal_6434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C ( clk ), .D ( new_AGEMA_signal_5861 ), .Q ( new_AGEMA_signal_6436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C ( clk ), .D ( new_AGEMA_signal_5863 ), .Q ( new_AGEMA_signal_6440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C ( clk ), .D ( new_AGEMA_signal_5865 ), .Q ( new_AGEMA_signal_6444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C ( clk ), .D ( n1930 ), .Q ( new_AGEMA_signal_6448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C ( clk ), .D ( new_AGEMA_signal_1130 ), .Q ( new_AGEMA_signal_6452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C ( clk ), .D ( new_AGEMA_signal_1131 ), .Q ( new_AGEMA_signal_6456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C ( clk ), .D ( n1976 ), .Q ( new_AGEMA_signal_6472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C ( clk ), .D ( new_AGEMA_signal_1178 ), .Q ( new_AGEMA_signal_6476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C ( clk ), .D ( new_AGEMA_signal_1179 ), .Q ( new_AGEMA_signal_6480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C ( clk ), .D ( new_AGEMA_signal_5609 ), .Q ( new_AGEMA_signal_6490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C ( clk ), .D ( new_AGEMA_signal_5611 ), .Q ( new_AGEMA_signal_6494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C ( clk ), .D ( new_AGEMA_signal_5613 ), .Q ( new_AGEMA_signal_6498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C ( clk ), .D ( n2008 ), .Q ( new_AGEMA_signal_6508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C ( clk ), .D ( new_AGEMA_signal_1376 ), .Q ( new_AGEMA_signal_6512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C ( clk ), .D ( new_AGEMA_signal_1377 ), .Q ( new_AGEMA_signal_6516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C ( clk ), .D ( n2022 ), .Q ( new_AGEMA_signal_6520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C ( clk ), .D ( new_AGEMA_signal_1386 ), .Q ( new_AGEMA_signal_6524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C ( clk ), .D ( new_AGEMA_signal_1387 ), .Q ( new_AGEMA_signal_6528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C ( clk ), .D ( n2057 ), .Q ( new_AGEMA_signal_6556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C ( clk ), .D ( new_AGEMA_signal_1412 ), .Q ( new_AGEMA_signal_6560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C ( clk ), .D ( new_AGEMA_signal_1413 ), .Q ( new_AGEMA_signal_6564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C ( clk ), .D ( n2062 ), .Q ( new_AGEMA_signal_6568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C ( clk ), .D ( new_AGEMA_signal_1416 ), .Q ( new_AGEMA_signal_6572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C ( clk ), .D ( new_AGEMA_signal_1417 ), .Q ( new_AGEMA_signal_6576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C ( clk ), .D ( n2075 ), .Q ( new_AGEMA_signal_6580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C ( clk ), .D ( new_AGEMA_signal_1208 ), .Q ( new_AGEMA_signal_6584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C ( clk ), .D ( new_AGEMA_signal_1209 ), .Q ( new_AGEMA_signal_6588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C ( clk ), .D ( n2121 ), .Q ( new_AGEMA_signal_6610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C ( clk ), .D ( new_AGEMA_signal_1440 ), .Q ( new_AGEMA_signal_6614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C ( clk ), .D ( new_AGEMA_signal_1441 ), .Q ( new_AGEMA_signal_6618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C ( clk ), .D ( new_AGEMA_signal_5579 ), .Q ( new_AGEMA_signal_6628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2143 ( .C ( clk ), .D ( new_AGEMA_signal_5581 ), .Q ( new_AGEMA_signal_6632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2147 ( .C ( clk ), .D ( new_AGEMA_signal_5583 ), .Q ( new_AGEMA_signal_6636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2153 ( .C ( clk ), .D ( new_AGEMA_signal_6641 ), .Q ( new_AGEMA_signal_6642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C ( clk ), .D ( new_AGEMA_signal_6647 ), .Q ( new_AGEMA_signal_6648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2165 ( .C ( clk ), .D ( new_AGEMA_signal_6653 ), .Q ( new_AGEMA_signal_6654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2169 ( .C ( clk ), .D ( new_AGEMA_signal_5795 ), .Q ( new_AGEMA_signal_6658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2173 ( .C ( clk ), .D ( new_AGEMA_signal_5797 ), .Q ( new_AGEMA_signal_6662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2177 ( .C ( clk ), .D ( new_AGEMA_signal_5799 ), .Q ( new_AGEMA_signal_6666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2181 ( .C ( clk ), .D ( new_AGEMA_signal_5837 ), .Q ( new_AGEMA_signal_6670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2185 ( .C ( clk ), .D ( new_AGEMA_signal_5839 ), .Q ( new_AGEMA_signal_6674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2189 ( .C ( clk ), .D ( new_AGEMA_signal_5841 ), .Q ( new_AGEMA_signal_6678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2217 ( .C ( clk ), .D ( n2245 ), .Q ( new_AGEMA_signal_6706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2221 ( .C ( clk ), .D ( new_AGEMA_signal_1498 ), .Q ( new_AGEMA_signal_6710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2225 ( .C ( clk ), .D ( new_AGEMA_signal_1499 ), .Q ( new_AGEMA_signal_6714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2231 ( .C ( clk ), .D ( new_AGEMA_signal_6719 ), .Q ( new_AGEMA_signal_6720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2237 ( .C ( clk ), .D ( new_AGEMA_signal_6725 ), .Q ( new_AGEMA_signal_6726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2243 ( .C ( clk ), .D ( new_AGEMA_signal_6731 ), .Q ( new_AGEMA_signal_6732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2247 ( .C ( clk ), .D ( n2262 ), .Q ( new_AGEMA_signal_6736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2251 ( .C ( clk ), .D ( new_AGEMA_signal_1240 ), .Q ( new_AGEMA_signal_6740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C ( clk ), .D ( new_AGEMA_signal_1241 ), .Q ( new_AGEMA_signal_6744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2277 ( .C ( clk ), .D ( n2343 ), .Q ( new_AGEMA_signal_6766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2281 ( .C ( clk ), .D ( new_AGEMA_signal_1532 ), .Q ( new_AGEMA_signal_6770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2285 ( .C ( clk ), .D ( new_AGEMA_signal_1533 ), .Q ( new_AGEMA_signal_6774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2301 ( .C ( clk ), .D ( new_AGEMA_signal_5801 ), .Q ( new_AGEMA_signal_6790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2305 ( .C ( clk ), .D ( new_AGEMA_signal_5803 ), .Q ( new_AGEMA_signal_6794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2309 ( .C ( clk ), .D ( new_AGEMA_signal_5805 ), .Q ( new_AGEMA_signal_6798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2313 ( .C ( clk ), .D ( new_AGEMA_signal_5777 ), .Q ( new_AGEMA_signal_6802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2317 ( .C ( clk ), .D ( new_AGEMA_signal_5779 ), .Q ( new_AGEMA_signal_6806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2321 ( .C ( clk ), .D ( new_AGEMA_signal_5781 ), .Q ( new_AGEMA_signal_6810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2325 ( .C ( clk ), .D ( new_AGEMA_signal_5567 ), .Q ( new_AGEMA_signal_6814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2329 ( .C ( clk ), .D ( new_AGEMA_signal_5569 ), .Q ( new_AGEMA_signal_6818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2333 ( .C ( clk ), .D ( new_AGEMA_signal_5571 ), .Q ( new_AGEMA_signal_6822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2337 ( .C ( clk ), .D ( new_AGEMA_signal_5645 ), .Q ( new_AGEMA_signal_6826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2341 ( .C ( clk ), .D ( new_AGEMA_signal_5647 ), .Q ( new_AGEMA_signal_6830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2345 ( .C ( clk ), .D ( new_AGEMA_signal_5649 ), .Q ( new_AGEMA_signal_6834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2349 ( .C ( clk ), .D ( n2417 ), .Q ( new_AGEMA_signal_6838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2353 ( .C ( clk ), .D ( new_AGEMA_signal_1706 ), .Q ( new_AGEMA_signal_6842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2357 ( .C ( clk ), .D ( new_AGEMA_signal_1707 ), .Q ( new_AGEMA_signal_6846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2385 ( .C ( clk ), .D ( new_AGEMA_signal_5855 ), .Q ( new_AGEMA_signal_6874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2389 ( .C ( clk ), .D ( new_AGEMA_signal_5857 ), .Q ( new_AGEMA_signal_6878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2393 ( .C ( clk ), .D ( new_AGEMA_signal_5859 ), .Q ( new_AGEMA_signal_6882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2397 ( .C ( clk ), .D ( n2483 ), .Q ( new_AGEMA_signal_6886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2401 ( .C ( clk ), .D ( new_AGEMA_signal_1272 ), .Q ( new_AGEMA_signal_6890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2405 ( .C ( clk ), .D ( new_AGEMA_signal_1273 ), .Q ( new_AGEMA_signal_6894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2463 ( .C ( clk ), .D ( n2629 ), .Q ( new_AGEMA_signal_6952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2467 ( .C ( clk ), .D ( new_AGEMA_signal_1298 ), .Q ( new_AGEMA_signal_6956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2471 ( .C ( clk ), .D ( new_AGEMA_signal_1299 ), .Q ( new_AGEMA_signal_6960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2505 ( .C ( clk ), .D ( n2736 ), .Q ( new_AGEMA_signal_6994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2509 ( .C ( clk ), .D ( new_AGEMA_signal_1160 ), .Q ( new_AGEMA_signal_6998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2513 ( .C ( clk ), .D ( new_AGEMA_signal_1161 ), .Q ( new_AGEMA_signal_7002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2517 ( .C ( clk ), .D ( new_AGEMA_signal_5723 ), .Q ( new_AGEMA_signal_7006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2521 ( .C ( clk ), .D ( new_AGEMA_signal_5725 ), .Q ( new_AGEMA_signal_7010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2525 ( .C ( clk ), .D ( new_AGEMA_signal_5727 ), .Q ( new_AGEMA_signal_7014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2529 ( .C ( clk ), .D ( new_AGEMA_signal_5639 ), .Q ( new_AGEMA_signal_7018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2533 ( .C ( clk ), .D ( new_AGEMA_signal_5641 ), .Q ( new_AGEMA_signal_7022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2537 ( .C ( clk ), .D ( new_AGEMA_signal_5643 ), .Q ( new_AGEMA_signal_7026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2541 ( .C ( clk ), .D ( n2787 ), .Q ( new_AGEMA_signal_7030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2545 ( .C ( clk ), .D ( new_AGEMA_signal_1664 ), .Q ( new_AGEMA_signal_7034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2549 ( .C ( clk ), .D ( new_AGEMA_signal_1665 ), .Q ( new_AGEMA_signal_7038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2579 ( .C ( clk ), .D ( new_AGEMA_signal_7067 ), .Q ( new_AGEMA_signal_7068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2587 ( .C ( clk ), .D ( new_AGEMA_signal_7075 ), .Q ( new_AGEMA_signal_7076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2595 ( .C ( clk ), .D ( new_AGEMA_signal_7083 ), .Q ( new_AGEMA_signal_7084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2609 ( .C ( clk ), .D ( new_AGEMA_signal_7097 ), .Q ( new_AGEMA_signal_7098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2617 ( .C ( clk ), .D ( new_AGEMA_signal_7105 ), .Q ( new_AGEMA_signal_7106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2625 ( .C ( clk ), .D ( new_AGEMA_signal_7113 ), .Q ( new_AGEMA_signal_7114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2631 ( .C ( clk ), .D ( n2009 ), .Q ( new_AGEMA_signal_7120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2637 ( .C ( clk ), .D ( new_AGEMA_signal_1382 ), .Q ( new_AGEMA_signal_7126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2643 ( .C ( clk ), .D ( new_AGEMA_signal_1383 ), .Q ( new_AGEMA_signal_7132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2661 ( .C ( clk ), .D ( n2034 ), .Q ( new_AGEMA_signal_7150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2667 ( .C ( clk ), .D ( new_AGEMA_signal_1202 ), .Q ( new_AGEMA_signal_7156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2673 ( .C ( clk ), .D ( new_AGEMA_signal_1203 ), .Q ( new_AGEMA_signal_7162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2685 ( .C ( clk ), .D ( new_AGEMA_signal_5849 ), .Q ( new_AGEMA_signal_7174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2691 ( .C ( clk ), .D ( new_AGEMA_signal_5851 ), .Q ( new_AGEMA_signal_7180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2697 ( .C ( clk ), .D ( new_AGEMA_signal_5853 ), .Q ( new_AGEMA_signal_7186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2703 ( .C ( clk ), .D ( new_AGEMA_signal_5891 ), .Q ( new_AGEMA_signal_7192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2709 ( .C ( clk ), .D ( new_AGEMA_signal_5893 ), .Q ( new_AGEMA_signal_7198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2715 ( .C ( clk ), .D ( new_AGEMA_signal_5895 ), .Q ( new_AGEMA_signal_7204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2739 ( .C ( clk ), .D ( new_AGEMA_signal_5513 ), .Q ( new_AGEMA_signal_7228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2745 ( .C ( clk ), .D ( new_AGEMA_signal_5515 ), .Q ( new_AGEMA_signal_7234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2751 ( .C ( clk ), .D ( new_AGEMA_signal_5517 ), .Q ( new_AGEMA_signal_7240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2757 ( .C ( clk ), .D ( n2122 ), .Q ( new_AGEMA_signal_7246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2763 ( .C ( clk ), .D ( new_AGEMA_signal_1444 ), .Q ( new_AGEMA_signal_7252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2769 ( .C ( clk ), .D ( new_AGEMA_signal_1445 ), .Q ( new_AGEMA_signal_7258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2781 ( .C ( clk ), .D ( n2220 ), .Q ( new_AGEMA_signal_7270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2787 ( .C ( clk ), .D ( new_AGEMA_signal_1456 ), .Q ( new_AGEMA_signal_7276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2793 ( .C ( clk ), .D ( new_AGEMA_signal_1457 ), .Q ( new_AGEMA_signal_7282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2837 ( .C ( clk ), .D ( new_AGEMA_signal_7325 ), .Q ( new_AGEMA_signal_7326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2845 ( .C ( clk ), .D ( new_AGEMA_signal_7333 ), .Q ( new_AGEMA_signal_7334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2853 ( .C ( clk ), .D ( new_AGEMA_signal_7341 ), .Q ( new_AGEMA_signal_7342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2859 ( .C ( clk ), .D ( new_AGEMA_signal_5663 ), .Q ( new_AGEMA_signal_7348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2865 ( .C ( clk ), .D ( new_AGEMA_signal_5665 ), .Q ( new_AGEMA_signal_7354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2871 ( .C ( clk ), .D ( new_AGEMA_signal_5667 ), .Q ( new_AGEMA_signal_7360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2943 ( .C ( clk ), .D ( n2344 ), .Q ( new_AGEMA_signal_7432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2949 ( .C ( clk ), .D ( new_AGEMA_signal_1536 ), .Q ( new_AGEMA_signal_7438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2955 ( .C ( clk ), .D ( new_AGEMA_signal_1537 ), .Q ( new_AGEMA_signal_7444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3039 ( .C ( clk ), .D ( n2468 ), .Q ( new_AGEMA_signal_7528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3045 ( .C ( clk ), .D ( new_AGEMA_signal_1278 ), .Q ( new_AGEMA_signal_7534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3051 ( .C ( clk ), .D ( new_AGEMA_signal_1279 ), .Q ( new_AGEMA_signal_7540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3057 ( .C ( clk ), .D ( n2761 ), .Q ( new_AGEMA_signal_7546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3063 ( .C ( clk ), .D ( new_AGEMA_signal_1346 ), .Q ( new_AGEMA_signal_7552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3069 ( .C ( clk ), .D ( new_AGEMA_signal_1347 ), .Q ( new_AGEMA_signal_7558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3095 ( .C ( clk ), .D ( new_AGEMA_signal_7583 ), .Q ( new_AGEMA_signal_7584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3103 ( .C ( clk ), .D ( new_AGEMA_signal_7591 ), .Q ( new_AGEMA_signal_7592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3111 ( .C ( clk ), .D ( new_AGEMA_signal_7599 ), .Q ( new_AGEMA_signal_7600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3185 ( .C ( clk ), .D ( new_AGEMA_signal_7673 ), .Q ( new_AGEMA_signal_7674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3193 ( .C ( clk ), .D ( new_AGEMA_signal_7681 ), .Q ( new_AGEMA_signal_7682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3201 ( .C ( clk ), .D ( new_AGEMA_signal_7689 ), .Q ( new_AGEMA_signal_7690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3231 ( .C ( clk ), .D ( n2825 ), .Q ( new_AGEMA_signal_7720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3237 ( .C ( clk ), .D ( new_AGEMA_signal_1674 ), .Q ( new_AGEMA_signal_7726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3243 ( .C ( clk ), .D ( new_AGEMA_signal_1675 ), .Q ( new_AGEMA_signal_7732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3255 ( .C ( clk ), .D ( n1957 ), .Q ( new_AGEMA_signal_7744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3263 ( .C ( clk ), .D ( new_AGEMA_signal_1156 ), .Q ( new_AGEMA_signal_7752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3271 ( .C ( clk ), .D ( new_AGEMA_signal_1157 ), .Q ( new_AGEMA_signal_7760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3297 ( .C ( clk ), .D ( n2026 ), .Q ( new_AGEMA_signal_7786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3305 ( .C ( clk ), .D ( new_AGEMA_signal_1196 ), .Q ( new_AGEMA_signal_7794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3313 ( .C ( clk ), .D ( new_AGEMA_signal_1197 ), .Q ( new_AGEMA_signal_7802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3357 ( .C ( clk ), .D ( n2811 ), .Q ( new_AGEMA_signal_7846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3365 ( .C ( clk ), .D ( new_AGEMA_signal_1446 ), .Q ( new_AGEMA_signal_7854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3373 ( .C ( clk ), .D ( new_AGEMA_signal_1447 ), .Q ( new_AGEMA_signal_7862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3495 ( .C ( clk ), .D ( new_AGEMA_signal_5909 ), .Q ( new_AGEMA_signal_7984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3503 ( .C ( clk ), .D ( new_AGEMA_signal_5911 ), .Q ( new_AGEMA_signal_7992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3511 ( .C ( clk ), .D ( new_AGEMA_signal_5913 ), .Q ( new_AGEMA_signal_8000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3549 ( .C ( clk ), .D ( n2363 ), .Q ( new_AGEMA_signal_8038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3557 ( .C ( clk ), .D ( new_AGEMA_signal_1262 ), .Q ( new_AGEMA_signal_8046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3565 ( .C ( clk ), .D ( new_AGEMA_signal_1263 ), .Q ( new_AGEMA_signal_8054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3645 ( .C ( clk ), .D ( new_AGEMA_signal_5843 ), .Q ( new_AGEMA_signal_8134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3653 ( .C ( clk ), .D ( new_AGEMA_signal_5845 ), .Q ( new_AGEMA_signal_8142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3661 ( .C ( clk ), .D ( new_AGEMA_signal_5847 ), .Q ( new_AGEMA_signal_8150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3669 ( .C ( clk ), .D ( new_AGEMA_signal_5543 ), .Q ( new_AGEMA_signal_8158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3677 ( .C ( clk ), .D ( new_AGEMA_signal_5545 ), .Q ( new_AGEMA_signal_8166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3685 ( .C ( clk ), .D ( new_AGEMA_signal_5547 ), .Q ( new_AGEMA_signal_8174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3927 ( .C ( clk ), .D ( n2544 ), .Q ( new_AGEMA_signal_8416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3937 ( .C ( clk ), .D ( new_AGEMA_signal_1216 ), .Q ( new_AGEMA_signal_8426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3947 ( .C ( clk ), .D ( new_AGEMA_signal_1217 ), .Q ( new_AGEMA_signal_8436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4077 ( .C ( clk ), .D ( n2364 ), .Q ( new_AGEMA_signal_8566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4087 ( .C ( clk ), .D ( new_AGEMA_signal_1548 ), .Q ( new_AGEMA_signal_8576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4097 ( .C ( clk ), .D ( new_AGEMA_signal_1549 ), .Q ( new_AGEMA_signal_8586 ) ) ;

    /* cells in depth 6 */
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1960 ( .a ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, n2575}), .b ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, n1962}), .clk ( clk ), .r ({Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, n1924}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1967 ( .a ({new_AGEMA_signal_1317, new_AGEMA_signal_1316, n1922}), .b ({new_AGEMA_signal_5511, new_AGEMA_signal_5509, new_AGEMA_signal_5507}), .clk ( clk ), .r ({Fresh[719], Fresh[718], Fresh[717]}), .c ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, n1923}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1981 ( .a ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, n1926}), .b ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, n1925}), .clk ( clk ), .r ({Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, n1927}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1993 ( .a ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, n2734}), .b ({new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2763}), .clk ( clk ), .r ({Fresh[725], Fresh[724], Fresh[723]}), .c ({new_AGEMA_signal_1683, new_AGEMA_signal_1682, n1929}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2007 ( .a ({new_AGEMA_signal_5517, new_AGEMA_signal_5515, new_AGEMA_signal_5513}), .b ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, n2732}), .clk ( clk ), .r ({Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, n2665}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2011 ( .a ({new_AGEMA_signal_5523, new_AGEMA_signal_5521, new_AGEMA_signal_5519}), .b ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, n1937}), .clk ( clk ), .r ({Fresh[731], Fresh[730], Fresh[729]}), .c ({new_AGEMA_signal_1687, new_AGEMA_signal_1686, n1938}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2019 ( .a ({new_AGEMA_signal_5529, new_AGEMA_signal_5527, new_AGEMA_signal_5525}), .b ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, n2732}), .clk ( clk ), .r ({Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, n2235}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2023 ( .a ({new_AGEMA_signal_5535, new_AGEMA_signal_5533, new_AGEMA_signal_5531}), .b ({new_AGEMA_signal_1143, new_AGEMA_signal_1142, n1942}), .clk ( clk ), .r ({Fresh[737], Fresh[736], Fresh[735]}), .c ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, n1943}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2027 ( .a ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, n2676}), .b ({new_AGEMA_signal_5541, new_AGEMA_signal_5539, new_AGEMA_signal_5537}), .clk ( clk ), .r ({Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, n1946}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2031 ( .a ({new_AGEMA_signal_5547, new_AGEMA_signal_5545, new_AGEMA_signal_5543}), .b ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, n1944}), .clk ( clk ), .r ({Fresh[743], Fresh[742], Fresh[741]}), .c ({new_AGEMA_signal_1691, new_AGEMA_signal_1690, n1945}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2034 ( .a ({new_AGEMA_signal_5553, new_AGEMA_signal_5551, new_AGEMA_signal_5549}), .b ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, n2734}), .clk ( clk ), .r ({Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_1693, new_AGEMA_signal_1692, n1956}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2040 ( .a ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, n1950}), .b ({new_AGEMA_signal_1151, new_AGEMA_signal_1150, n1949}), .clk ( clk ), .r ({Fresh[749], Fresh[748], Fresh[747]}), .c ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, n1951}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2048 ( .a ({new_AGEMA_signal_1341, new_AGEMA_signal_1340, n2662}), .b ({new_AGEMA_signal_1155, new_AGEMA_signal_1154, n2627}), .clk ( clk ), .r ({Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, n1952}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2057 ( .a ({new_AGEMA_signal_5559, new_AGEMA_signal_5557, new_AGEMA_signal_5555}), .b ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, n2088}), .clk ( clk ), .r ({Fresh[755], Fresh[754], Fresh[753]}), .c ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, n2687}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) U2061 ( .a ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, n1962}), .b ({new_AGEMA_signal_5565, new_AGEMA_signal_5563, new_AGEMA_signal_5561}), .clk ( clk ), .r ({Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, n1966}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2064 ( .a ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, n2736}), .b ({new_AGEMA_signal_5571, new_AGEMA_signal_5569, new_AGEMA_signal_5567}), .clk ( clk ), .r ({Fresh[761], Fresh[760], Fresh[759]}), .c ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, n1963}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2077 ( .a ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, n2720}), .b ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, n2417}), .clk ( clk ), .r ({Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, n1968}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2082 ( .a ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, n2505}), .b ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2651}), .clk ( clk ), .r ({Fresh[767], Fresh[766], Fresh[765]}), .c ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, n2684}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2088 ( .a ({new_AGEMA_signal_5577, new_AGEMA_signal_5575, new_AGEMA_signal_5573}), .b ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, n2625}), .clk ( clk ), .r ({Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_1711, new_AGEMA_signal_1710, n1972}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2092 ( .a ({new_AGEMA_signal_5583, new_AGEMA_signal_5581, new_AGEMA_signal_5579}), .b ({new_AGEMA_signal_1177, new_AGEMA_signal_1176, n2190}), .clk ( clk ), .r ({Fresh[773], Fresh[772], Fresh[771]}), .c ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, n1971}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2099 ( .a ({new_AGEMA_signal_5589, new_AGEMA_signal_5587, new_AGEMA_signal_5585}), .b ({new_AGEMA_signal_1359, new_AGEMA_signal_1358, n2535}), .clk ( clk ), .r ({Fresh[776], Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, n1974}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2106 ( .a ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, n2732}), .b ({new_AGEMA_signal_5559, new_AGEMA_signal_5557, new_AGEMA_signal_5555}), .clk ( clk ), .r ({Fresh[779], Fresh[778], Fresh[777]}), .c ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, n1979}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2112 ( .a ({new_AGEMA_signal_5595, new_AGEMA_signal_5593, new_AGEMA_signal_5591}), .b ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2817}), .clk ( clk ), .r ({Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, n1985}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2121 ( .a ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, n1992}), .b ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, n1991}), .clk ( clk ), .r ({Fresh[785], Fresh[784], Fresh[783]}), .c ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, n1994}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2126 ( .a ({new_AGEMA_signal_5601, new_AGEMA_signal_5599, new_AGEMA_signal_5597}), .b ({new_AGEMA_signal_1371, new_AGEMA_signal_1370, n1995}), .clk ( clk ), .r ({Fresh[788], Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, n1996}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2136 ( .a ({new_AGEMA_signal_5607, new_AGEMA_signal_5605, new_AGEMA_signal_5603}), .b ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, n2003}), .clk ( clk ), .r ({Fresh[791], Fresh[790], Fresh[789]}), .c ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, n2137}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2142 ( .a ({new_AGEMA_signal_5613, new_AGEMA_signal_5611, new_AGEMA_signal_5609}), .b ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, n2572}), .clk ( clk ), .r ({Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, n2006}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2144 ( .a ({new_AGEMA_signal_5619, new_AGEMA_signal_5617, new_AGEMA_signal_5615}), .b ({new_AGEMA_signal_1381, new_AGEMA_signal_1380, n2004}), .clk ( clk ), .r ({Fresh[797], Fresh[796], Fresh[795]}), .c ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, n2005}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2152 ( .a ({new_AGEMA_signal_5625, new_AGEMA_signal_5623, new_AGEMA_signal_5621}), .b ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, n2533}), .clk ( clk ), .r ({Fresh[800], Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_1729, new_AGEMA_signal_1728, n2013}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2160 ( .a ({new_AGEMA_signal_5631, new_AGEMA_signal_5629, new_AGEMA_signal_5627}), .b ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, n2227}), .clk ( clk ), .r ({Fresh[803], Fresh[802], Fresh[801]}), .c ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, n2020}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2164 ( .a ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2817}), .b ({new_AGEMA_signal_5637, new_AGEMA_signal_5635, new_AGEMA_signal_5633}), .clk ( clk ), .r ({Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, n2023}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2168 ( .a ({new_AGEMA_signal_1077, new_AGEMA_signal_1076, n2027}), .b ({new_AGEMA_signal_5643, new_AGEMA_signal_5641, new_AGEMA_signal_5639}), .clk ( clk ), .r ({Fresh[809], Fresh[808], Fresh[807]}), .c ({new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2028}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2172 ( .a ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, n2214}), .b ({new_AGEMA_signal_5649, new_AGEMA_signal_5647, new_AGEMA_signal_5645}), .clk ( clk ), .r ({Fresh[812], Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, n2033}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2175 ( .a ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, n2376}), .b ({new_AGEMA_signal_5655, new_AGEMA_signal_5653, new_AGEMA_signal_5651}), .clk ( clk ), .r ({Fresh[815], Fresh[814], Fresh[813]}), .c ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, n2031}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2184 ( .a ({new_AGEMA_signal_1155, new_AGEMA_signal_1154, n2627}), .b ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2039}), .clk ( clk ), .r ({Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, n2040}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2187 ( .a ({new_AGEMA_signal_5661, new_AGEMA_signal_5659, new_AGEMA_signal_5657}), .b ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2651}), .clk ( clk ), .r ({Fresh[821], Fresh[820], Fresh[819]}), .c ({new_AGEMA_signal_1401, new_AGEMA_signal_1400, n2050}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2193 ( .a ({new_AGEMA_signal_5667, new_AGEMA_signal_5665, new_AGEMA_signal_5663}), .b ({new_AGEMA_signal_1407, new_AGEMA_signal_1406, n2044}), .clk ( clk ), .r ({Fresh[824], Fresh[823], Fresh[822]}), .c ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, n2045}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2199 ( .a ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, n2654}), .b ({new_AGEMA_signal_5559, new_AGEMA_signal_5557, new_AGEMA_signal_5555}), .clk ( clk ), .r ({Fresh[827], Fresh[826], Fresh[825]}), .c ({new_AGEMA_signal_1741, new_AGEMA_signal_1740, n2051}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2203 ( .a ({new_AGEMA_signal_5673, new_AGEMA_signal_5671, new_AGEMA_signal_5669}), .b ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, n2055}), .clk ( clk ), .r ({Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, n2056}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2209 ( .a ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, n2407}), .b ({new_AGEMA_signal_5679, new_AGEMA_signal_5677, new_AGEMA_signal_5675}), .clk ( clk ), .r ({Fresh[833], Fresh[832], Fresh[831]}), .c ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, n2060}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2215 ( .a ({new_AGEMA_signal_5685, new_AGEMA_signal_5683, new_AGEMA_signal_5681}), .b ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, n2654}), .clk ( clk ), .r ({Fresh[836], Fresh[835], Fresh[834]}), .c ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, n2066}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2217 ( .a ({new_AGEMA_signal_5643, new_AGEMA_signal_5641, new_AGEMA_signal_5639}), .b ({new_AGEMA_signal_1419, new_AGEMA_signal_1418, n2731}), .clk ( clk ), .r ({Fresh[839], Fresh[838], Fresh[837]}), .c ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, n2065}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2221 ( .a ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, n2068}), .b ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2817}), .clk ( clk ), .r ({Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, n2069}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2226 ( .a ({new_AGEMA_signal_5691, new_AGEMA_signal_5689, new_AGEMA_signal_5687}), .b ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, n2252}), .clk ( clk ), .r ({Fresh[845], Fresh[844], Fresh[843]}), .c ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, n2074}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2235 ( .a ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, n2081}), .b ({new_AGEMA_signal_1425, new_AGEMA_signal_1424, n2080}), .clk ( clk ), .r ({Fresh[848], Fresh[847], Fresh[846]}), .c ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, n2082}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2240 ( .a ({new_AGEMA_signal_5619, new_AGEMA_signal_5617, new_AGEMA_signal_5615}), .b ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, n2083}), .clk ( clk ), .r ({Fresh[851], Fresh[850], Fresh[849]}), .c ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, n2084}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2242 ( .a ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, n2533}), .b ({new_AGEMA_signal_5517, new_AGEMA_signal_5515, new_AGEMA_signal_5513}), .clk ( clk ), .r ({Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_1759, new_AGEMA_signal_1758, n2085}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2245 ( .a ({new_AGEMA_signal_5697, new_AGEMA_signal_5695, new_AGEMA_signal_5693}), .b ({new_AGEMA_signal_1431, new_AGEMA_signal_1430, n2562}), .clk ( clk ), .r ({Fresh[857], Fresh[856], Fresh[855]}), .c ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, n2131}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2248 ( .a ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, n2088}), .b ({new_AGEMA_signal_1215, new_AGEMA_signal_1214, n2087}), .clk ( clk ), .r ({Fresh[860], Fresh[859], Fresh[858]}), .c ({new_AGEMA_signal_1763, new_AGEMA_signal_1762, n2089}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2252 ( .a ({new_AGEMA_signal_5649, new_AGEMA_signal_5647, new_AGEMA_signal_5645}), .b ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, n2156}), .clk ( clk ), .r ({Fresh[863], Fresh[862], Fresh[861]}), .c ({new_AGEMA_signal_1765, new_AGEMA_signal_1764, n2330}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2254 ( .a ({new_AGEMA_signal_5703, new_AGEMA_signal_5701, new_AGEMA_signal_5699}), .b ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, n2151}), .clk ( clk ), .r ({Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, n2092}) ) ;
    or_HPC2 #(.security_order(2), .pipeline(1)) U2256 ( .a ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, n2761}), .b ({new_AGEMA_signal_1353, new_AGEMA_signal_1352, n2359}), .clk ( clk ), .r ({Fresh[869], Fresh[868], Fresh[867]}), .c ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, n2094}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2261 ( .a ({new_AGEMA_signal_1173, new_AGEMA_signal_1172, n2101}), .b ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, n2100}), .clk ( clk ), .r ({Fresh[872], Fresh[871], Fresh[870]}), .c ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, n2160}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2265 ( .a ({new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2492}), .b ({new_AGEMA_signal_5649, new_AGEMA_signal_5647, new_AGEMA_signal_5645}), .clk ( clk ), .r ({Fresh[875], Fresh[874], Fresh[873]}), .c ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, n2504}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2271 ( .a ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, n2417}), .b ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2651}), .clk ( clk ), .r ({Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, n2114}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2273 ( .a ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, n2677}), .b ({new_AGEMA_signal_5619, new_AGEMA_signal_5617, new_AGEMA_signal_5615}), .clk ( clk ), .r ({Fresh[881], Fresh[880], Fresh[879]}), .c ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, n2115}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2280 ( .a ({new_AGEMA_signal_5709, new_AGEMA_signal_5707, new_AGEMA_signal_5705}), .b ({new_AGEMA_signal_1419, new_AGEMA_signal_1418, n2731}), .clk ( clk ), .r ({Fresh[884], Fresh[883], Fresh[882]}), .c ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, n2291}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2281 ( .a ({new_AGEMA_signal_5517, new_AGEMA_signal_5515, new_AGEMA_signal_5513}), .b ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, n2498}), .clk ( clk ), .r ({Fresh[887], Fresh[886], Fresh[885]}), .c ({new_AGEMA_signal_1443, new_AGEMA_signal_1442, n2119}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2291 ( .a ({new_AGEMA_signal_5715, new_AGEMA_signal_5713, new_AGEMA_signal_5711}), .b ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, n2498}), .clk ( clk ), .r ({Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, n2130}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2292 ( .a ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2817}), .b ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, n2631}), .clk ( clk ), .r ({Fresh[893], Fresh[892], Fresh[891]}), .c ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, n2129}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2295 ( .a ({new_AGEMA_signal_1221, new_AGEMA_signal_1220, n2647}), .b ({new_AGEMA_signal_5721, new_AGEMA_signal_5719, new_AGEMA_signal_5717}), .clk ( clk ), .r ({Fresh[896], Fresh[895], Fresh[894]}), .c ({new_AGEMA_signal_1453, new_AGEMA_signal_1452, n2150}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2298 ( .a ({new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2492}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, n2132}), .clk ( clk ), .r ({Fresh[899], Fresh[898], Fresh[897]}), .c ({new_AGEMA_signal_1455, new_AGEMA_signal_1454, n2133}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2302 ( .a ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, n2533}), .b ({new_AGEMA_signal_5727, new_AGEMA_signal_5725, new_AGEMA_signal_5723}), .clk ( clk ), .r ({Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, n2136}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2306 ( .a ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, n2572}), .b ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, n2138}), .clk ( clk ), .r ({Fresh[905], Fresh[904], Fresh[903]}), .c ({new_AGEMA_signal_1783, new_AGEMA_signal_1782, n2139}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2313 ( .a ({new_AGEMA_signal_5733, new_AGEMA_signal_5731, new_AGEMA_signal_5729}), .b ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, n2555}), .clk ( clk ), .r ({Fresh[908], Fresh[907], Fresh[906]}), .c ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, n2144}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2318 ( .a ({new_AGEMA_signal_1323, new_AGEMA_signal_1322, n2151}), .b ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, n2533}), .clk ( clk ), .r ({Fresh[911], Fresh[910], Fresh[909]}), .c ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, n2152}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2321 ( .a ({new_AGEMA_signal_1155, new_AGEMA_signal_1154, n2627}), .b ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, n2156}), .clk ( clk ), .r ({Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, n2170}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2323 ( .a ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, n2429}), .b ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, n2732}), .clk ( clk ), .r ({Fresh[917], Fresh[916], Fresh[915]}), .c ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, n2157}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2329 ( .a ({new_AGEMA_signal_5739, new_AGEMA_signal_5737, new_AGEMA_signal_5735}), .b ({new_AGEMA_signal_1225, new_AGEMA_signal_1224, n2162}), .clk ( clk ), .r ({Fresh[920], Fresh[919], Fresh[918]}), .c ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, n2163}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2335 ( .a ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, n2171}), .b ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, n2376}), .clk ( clk ), .r ({Fresh[923], Fresh[922], Fresh[921]}), .c ({new_AGEMA_signal_1795, new_AGEMA_signal_1794, n2172}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2338 ( .a ({new_AGEMA_signal_5517, new_AGEMA_signal_5515, new_AGEMA_signal_5513}), .b ({new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2545}), .clk ( clk ), .r ({Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_1227, new_AGEMA_signal_1226, n2186}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2339 ( .a ({new_AGEMA_signal_5589, new_AGEMA_signal_5587, new_AGEMA_signal_5585}), .b ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, n2290}), .clk ( clk ), .r ({Fresh[929], Fresh[928], Fresh[927]}), .c ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, n2181}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2344 ( .a ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, n2176}), .b ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, n2175}), .clk ( clk ), .r ({Fresh[932], Fresh[931], Fresh[930]}), .c ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, n2177}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2349 ( .a ({new_AGEMA_signal_5559, new_AGEMA_signal_5557, new_AGEMA_signal_5555}), .b ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, n2182}), .clk ( clk ), .r ({Fresh[935], Fresh[934], Fresh[933]}), .c ({new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2183}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2354 ( .a ({new_AGEMA_signal_5745, new_AGEMA_signal_5743, new_AGEMA_signal_5741}), .b ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, n2188}), .clk ( clk ), .r ({Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_1801, new_AGEMA_signal_1800, n2195}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2356 ( .a ({new_AGEMA_signal_1177, new_AGEMA_signal_1176, n2190}), .b ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, n2189}), .clk ( clk ), .r ({Fresh[941], Fresh[940], Fresh[939]}), .c ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, n2193}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2358 ( .a ({new_AGEMA_signal_5751, new_AGEMA_signal_5749, new_AGEMA_signal_5747}), .b ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, n2446}), .clk ( clk ), .r ({Fresh[944], Fresh[943], Fresh[942]}), .c ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, n2191}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2364 ( .a ({new_AGEMA_signal_1233, new_AGEMA_signal_1232, n2576}), .b ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, n2748}), .clk ( clk ), .r ({Fresh[947], Fresh[946], Fresh[945]}), .c ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, n2196}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2367 ( .a ({new_AGEMA_signal_5541, new_AGEMA_signal_5539, new_AGEMA_signal_5537}), .b ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, n2505}), .clk ( clk ), .r ({Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, n2201}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2369 ( .a ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, n2674}), .b ({new_AGEMA_signal_5757, new_AGEMA_signal_5755, new_AGEMA_signal_5753}), .clk ( clk ), .r ({Fresh[953], Fresh[952], Fresh[951]}), .c ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2200}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) U2371 ( .s ({new_AGEMA_signal_5721, new_AGEMA_signal_5719, new_AGEMA_signal_5717}), .b ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, n2734}), .a ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, n2417}), .clk ( clk ), .r ({Fresh[956], Fresh[955], Fresh[954]}), .c ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, n2202}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2379 ( .a ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, n2214}), .b ({new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2213}), .clk ( clk ), .r ({Fresh[959], Fresh[958], Fresh[957]}), .c ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, n2217}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2381 ( .a ({new_AGEMA_signal_5763, new_AGEMA_signal_5761, new_AGEMA_signal_5759}), .b ({new_AGEMA_signal_1239, new_AGEMA_signal_1238, n2215}), .clk ( clk ), .r ({Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, n2216}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2385 ( .a ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, n2218}), .b ({new_AGEMA_signal_5751, new_AGEMA_signal_5749, new_AGEMA_signal_5747}), .clk ( clk ), .r ({Fresh[965], Fresh[964], Fresh[963]}), .c ({new_AGEMA_signal_1813, new_AGEMA_signal_1812, n2222}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2387 ( .a ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, n2220}), .b ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, n2219}), .clk ( clk ), .r ({Fresh[968], Fresh[967], Fresh[966]}), .c ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, n2221}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2391 ( .a ({new_AGEMA_signal_1155, new_AGEMA_signal_1154, n2627}), .b ({new_AGEMA_signal_5769, new_AGEMA_signal_5767, new_AGEMA_signal_5765}), .clk ( clk ), .r ({Fresh[971], Fresh[970], Fresh[969]}), .c ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, n2226}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) U2393 ( .s ({new_AGEMA_signal_5721, new_AGEMA_signal_5719, new_AGEMA_signal_5717}), .b ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2651}), .a ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, n2227}), .clk ( clk ), .r ({Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, n2228}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2397 ( .a ({new_AGEMA_signal_5631, new_AGEMA_signal_5629, new_AGEMA_signal_5627}), .b ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2651}), .clk ( clk ), .r ({Fresh[977], Fresh[976], Fresh[975]}), .c ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, n2237}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2398 ( .a ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, n2417}), .b ({new_AGEMA_signal_5721, new_AGEMA_signal_5719, new_AGEMA_signal_5717}), .clk ( clk ), .r ({Fresh[980], Fresh[979], Fresh[978]}), .c ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, n2233}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2403 ( .a ({new_AGEMA_signal_5775, new_AGEMA_signal_5773, new_AGEMA_signal_5771}), .b ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, n2631}), .clk ( clk ), .r ({Fresh[983], Fresh[982], Fresh[981]}), .c ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, n2238}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2406 ( .a ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, n2241}), .b ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, n2240}), .clk ( clk ), .r ({Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_1819, new_AGEMA_signal_1818, n2248}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2409 ( .a ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, n2561}), .b ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, n2243}), .clk ( clk ), .r ({Fresh[989], Fresh[988], Fresh[987]}), .c ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, n2244}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2414 ( .a ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, n2376}), .b ({new_AGEMA_signal_5511, new_AGEMA_signal_5509, new_AGEMA_signal_5507}), .clk ( clk ), .r ({Fresh[992], Fresh[991], Fresh[990]}), .c ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, n2249}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) U2417 ( .s ({new_AGEMA_signal_5721, new_AGEMA_signal_5719, new_AGEMA_signal_5717}), .b ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, n2252}), .a ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2651}), .clk ( clk ), .r ({Fresh[995], Fresh[994], Fresh[993]}), .c ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, n2253}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2424 ( .a ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, n2533}), .b ({new_AGEMA_signal_1503, new_AGEMA_signal_1502, n2259}), .clk ( clk ), .r ({Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, n2260}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2429 ( .a ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, n2417}), .b ({new_AGEMA_signal_5781, new_AGEMA_signal_5779, new_AGEMA_signal_5777}), .clk ( clk ), .r ({Fresh[1001], Fresh[1000], Fresh[999]}), .c ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, n2273}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2430 ( .a ({new_AGEMA_signal_5787, new_AGEMA_signal_5785, new_AGEMA_signal_5783}), .b ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, n2720}), .clk ( clk ), .r ({Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, n2752}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2433 ( .a ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, n2645}), .b ({new_AGEMA_signal_5709, new_AGEMA_signal_5707, new_AGEMA_signal_5705}), .clk ( clk ), .r ({Fresh[1007], Fresh[1006], Fresh[1005]}), .c ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, n2265}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2437 ( .a ({new_AGEMA_signal_5793, new_AGEMA_signal_5791, new_AGEMA_signal_5789}), .b ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, n2268}), .clk ( clk ), .r ({Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, n2269}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2444 ( .a ({new_AGEMA_signal_5571, new_AGEMA_signal_5569, new_AGEMA_signal_5567}), .b ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2817}), .clk ( clk ), .r ({Fresh[1013], Fresh[1012], Fresh[1011]}), .c ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, n2277}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2449 ( .a ({new_AGEMA_signal_5799, new_AGEMA_signal_5797, new_AGEMA_signal_5795}), .b ({new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2383}), .clk ( clk ), .r ({Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, n2282}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2452 ( .a ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, n2736}), .b ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, n2533}), .clk ( clk ), .r ({Fresh[1019], Fresh[1018], Fresh[1017]}), .c ({new_AGEMA_signal_1837, new_AGEMA_signal_1836, n2284}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2456 ( .a ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, n2774}), .b ({new_AGEMA_signal_5805, new_AGEMA_signal_5803, new_AGEMA_signal_5801}), .clk ( clk ), .r ({Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, n2459}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2459 ( .a ({new_AGEMA_signal_5523, new_AGEMA_signal_5521, new_AGEMA_signal_5519}), .b ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, n2287}), .clk ( clk ), .r ({Fresh[1025], Fresh[1024], Fresh[1023]}), .c ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, n2288}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2462 ( .a ({new_AGEMA_signal_5517, new_AGEMA_signal_5515, new_AGEMA_signal_5513}), .b ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, n2761}), .clk ( clk ), .r ({Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, n2458}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2464 ( .a ({new_AGEMA_signal_5739, new_AGEMA_signal_5737, new_AGEMA_signal_5735}), .b ({new_AGEMA_signal_1395, new_AGEMA_signal_1394, n2290}), .clk ( clk ), .r ({Fresh[1031], Fresh[1030], Fresh[1029]}), .c ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, n2293}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2467 ( .a ({new_AGEMA_signal_5703, new_AGEMA_signal_5701, new_AGEMA_signal_5699}), .b ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, n2642}), .clk ( clk ), .r ({Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, n2294}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2472 ( .a ({new_AGEMA_signal_1521, new_AGEMA_signal_1520, n2438}), .b ({new_AGEMA_signal_1251, new_AGEMA_signal_1250, n2299}), .clk ( clk ), .r ({Fresh[1037], Fresh[1036], Fresh[1035]}), .c ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, n2300}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2480 ( .a ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, n2734}), .b ({new_AGEMA_signal_5751, new_AGEMA_signal_5749, new_AGEMA_signal_5747}), .clk ( clk ), .r ({Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, n2323}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) U2482 ( .a ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, n2571}), .b ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, n2371}), .clk ( clk ), .r ({Fresh[1043], Fresh[1042], Fresh[1041]}), .c ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, n2314}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2485 ( .a ({new_AGEMA_signal_1095, new_AGEMA_signal_1094, n2316}), .b ({new_AGEMA_signal_5811, new_AGEMA_signal_5809, new_AGEMA_signal_5807}), .clk ( clk ), .r ({Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, n2319}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2491 ( .a ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, n2642}), .b ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, n2498}), .clk ( clk ), .r ({Fresh[1049], Fresh[1048], Fresh[1047]}), .c ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, n2326}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2496 ( .a ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, n2328}), .b ({new_AGEMA_signal_1257, new_AGEMA_signal_1256, n2327}), .clk ( clk ), .r ({Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, n2329}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2501 ( .a ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, n2417}), .b ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, n2674}), .clk ( clk ), .r ({Fresh[1055], Fresh[1054], Fresh[1053]}), .c ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, n2335}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2506 ( .a ({new_AGEMA_signal_5625, new_AGEMA_signal_5623, new_AGEMA_signal_5621}), .b ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, n2376}), .clk ( clk ), .r ({Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, n2341}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2507 ( .a ({new_AGEMA_signal_5817, new_AGEMA_signal_5815, new_AGEMA_signal_5813}), .b ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, n2736}), .clk ( clk ), .r ({Fresh[1061], Fresh[1060], Fresh[1059]}), .c ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, n2340}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2514 ( .a ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, n2348}), .b ({new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2347}), .clk ( clk ), .r ({Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, n2349}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2517 ( .a ({new_AGEMA_signal_5823, new_AGEMA_signal_5821, new_AGEMA_signal_5819}), .b ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, n2690}), .clk ( clk ), .r ({Fresh[1067], Fresh[1066], Fresh[1065]}), .c ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, n2375}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2518 ( .a ({new_AGEMA_signal_5733, new_AGEMA_signal_5731, new_AGEMA_signal_5729}), .b ({new_AGEMA_signal_1161, new_AGEMA_signal_1160, n2736}), .clk ( clk ), .r ({Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, n2352}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2522 ( .a ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, n2353}), .b ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, n2533}), .clk ( clk ), .r ({Fresh[1073], Fresh[1072], Fresh[1071]}), .c ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, n2354}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2525 ( .a ({new_AGEMA_signal_5829, new_AGEMA_signal_5827, new_AGEMA_signal_5825}), .b ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, n2355}), .clk ( clk ), .r ({Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, n2357}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2527 ( .a ({new_AGEMA_signal_1353, new_AGEMA_signal_1352, n2359}), .b ({new_AGEMA_signal_5835, new_AGEMA_signal_5833, new_AGEMA_signal_5831}), .clk ( clk ), .r ({Fresh[1079], Fresh[1078], Fresh[1077]}), .c ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, n2360}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2534 ( .a ({new_AGEMA_signal_5517, new_AGEMA_signal_5515, new_AGEMA_signal_5513}), .b ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, n2674}), .clk ( clk ), .r ({Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, n2369}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2536 ( .a ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, n2371}), .b ({new_AGEMA_signal_5769, new_AGEMA_signal_5767, new_AGEMA_signal_5765}), .clk ( clk ), .r ({Fresh[1085], Fresh[1084], Fresh[1083]}), .c ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, n2372}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2539 ( .a ({new_AGEMA_signal_1233, new_AGEMA_signal_1232, n2576}), .b ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, n2376}), .clk ( clk ), .r ({Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, n2377}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2544 ( .a ({new_AGEMA_signal_5751, new_AGEMA_signal_5749, new_AGEMA_signal_5747}), .b ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, n2415}), .clk ( clk ), .r ({Fresh[1091], Fresh[1090], Fresh[1089]}), .c ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, n2467}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2545 ( .a ({new_AGEMA_signal_5841, new_AGEMA_signal_5839, new_AGEMA_signal_5837}), .b ({new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2383}), .clk ( clk ), .r ({Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, n2385}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2546 ( .a ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2651}), .b ({new_AGEMA_signal_5649, new_AGEMA_signal_5647, new_AGEMA_signal_5645}), .clk ( clk ), .r ({Fresh[1097], Fresh[1096], Fresh[1095]}), .c ({new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2384}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2548 ( .a ({new_AGEMA_signal_5619, new_AGEMA_signal_5617, new_AGEMA_signal_5615}), .b ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, n2429}), .clk ( clk ), .r ({Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, n2386}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2552 ( .a ({new_AGEMA_signal_5745, new_AGEMA_signal_5743, new_AGEMA_signal_5741}), .b ({new_AGEMA_signal_1221, new_AGEMA_signal_1220, n2647}), .clk ( clk ), .r ({Fresh[1103], Fresh[1102], Fresh[1101]}), .c ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, n2394}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2553 ( .a ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2651}), .b ({new_AGEMA_signal_5751, new_AGEMA_signal_5749, new_AGEMA_signal_5747}), .clk ( clk ), .r ({Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, n2391}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2554 ( .a ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, n2505}), .b ({new_AGEMA_signal_5649, new_AGEMA_signal_5647, new_AGEMA_signal_5645}), .clk ( clk ), .r ({Fresh[1109], Fresh[1108], Fresh[1107]}), .c ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, n2390}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2559 ( .a ({new_AGEMA_signal_5703, new_AGEMA_signal_5701, new_AGEMA_signal_5699}), .b ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2700}), .clk ( clk ), .r ({Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2396}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2562 ( .a ({new_AGEMA_signal_5847, new_AGEMA_signal_5845, new_AGEMA_signal_5843}), .b ({new_AGEMA_signal_1521, new_AGEMA_signal_1520, n2438}), .clk ( clk ), .r ({Fresh[1115], Fresh[1114], Fresh[1113]}), .c ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, n2406}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2565 ( .a ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, n2594}), .b ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, n2402}), .clk ( clk ), .r ({Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, n2403}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2569 ( .a ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, n2407}), .b ({new_AGEMA_signal_5727, new_AGEMA_signal_5725, new_AGEMA_signal_5723}), .clk ( clk ), .r ({Fresh[1121], Fresh[1120], Fresh[1119]}), .c ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, n2408}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2573 ( .a ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, n2412}), .b ({new_AGEMA_signal_5775, new_AGEMA_signal_5773, new_AGEMA_signal_5771}), .clk ( clk ), .r ({Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, n2574}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2574 ( .a ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, n2498}), .b ({new_AGEMA_signal_5667, new_AGEMA_signal_5665, new_AGEMA_signal_5663}), .clk ( clk ), .r ({Fresh[1127], Fresh[1126], Fresh[1125]}), .c ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, n2413}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2577 ( .a ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, n2415}), .b ({new_AGEMA_signal_5649, new_AGEMA_signal_5647, new_AGEMA_signal_5645}), .clk ( clk ), .r ({Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, n2416}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2586 ( .a ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, n2428}), .b ({new_AGEMA_signal_5853, new_AGEMA_signal_5851, new_AGEMA_signal_5849}), .clk ( clk ), .r ({Fresh[1133], Fresh[1132], Fresh[1131]}), .c ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, n2433}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2587 ( .a ({new_AGEMA_signal_5517, new_AGEMA_signal_5515, new_AGEMA_signal_5513}), .b ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, n2429}), .clk ( clk ), .r ({Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, n2689}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2591 ( .a ({new_AGEMA_signal_1221, new_AGEMA_signal_1220, n2647}), .b ({new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2492}), .clk ( clk ), .r ({Fresh[1139], Fresh[1138], Fresh[1137]}), .c ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, n2434}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2595 ( .a ({new_AGEMA_signal_1521, new_AGEMA_signal_1520, n2438}), .b ({new_AGEMA_signal_1273, new_AGEMA_signal_1272, n2483}), .clk ( clk ), .r ({Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, n2439}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2598 ( .a ({new_AGEMA_signal_5841, new_AGEMA_signal_5839, new_AGEMA_signal_5837}), .b ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, n2540}), .clk ( clk ), .r ({Fresh[1145], Fresh[1144], Fresh[1143]}), .c ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, n2445}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2600 ( .a ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, n2690}), .b ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, n2443}), .clk ( clk ), .r ({Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, n2444}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2602 ( .a ({new_AGEMA_signal_5589, new_AGEMA_signal_5587, new_AGEMA_signal_5585}), .b ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, n2446}), .clk ( clk ), .r ({Fresh[1151], Fresh[1150], Fresh[1149]}), .c ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, n2447}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2607 ( .a ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, n2761}), .b ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, n2693}), .clk ( clk ), .r ({Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, n2454}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2617 ( .a ({new_AGEMA_signal_5709, new_AGEMA_signal_5707, new_AGEMA_signal_5705}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, n2464}), .clk ( clk ), .r ({Fresh[1157], Fresh[1156], Fresh[1155]}), .c ({new_AGEMA_signal_1579, new_AGEMA_signal_1578, n2465}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2622 ( .a ({new_AGEMA_signal_5721, new_AGEMA_signal_5719, new_AGEMA_signal_5717}), .b ({new_AGEMA_signal_1233, new_AGEMA_signal_1232, n2576}), .clk ( clk ), .r ({Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, n2470}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2626 ( .a ({new_AGEMA_signal_1281, new_AGEMA_signal_1280, n2473}), .b ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, n2472}), .clk ( clk ), .r ({Fresh[1163], Fresh[1162], Fresh[1161]}), .c ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, n2476}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2633 ( .a ({new_AGEMA_signal_5859, new_AGEMA_signal_5857, new_AGEMA_signal_5855}), .b ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, n2480}), .clk ( clk ), .r ({Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, n2481}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2639 ( .a ({new_AGEMA_signal_5865, new_AGEMA_signal_5863, new_AGEMA_signal_5861}), .b ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2817}), .clk ( clk ), .r ({Fresh[1169], Fresh[1168], Fresh[1167]}), .c ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, n2486}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2642 ( .a ({new_AGEMA_signal_5787, new_AGEMA_signal_5785, new_AGEMA_signal_5783}), .b ({new_AGEMA_signal_1287, new_AGEMA_signal_1286, n2488}), .clk ( clk ), .r ({Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({new_AGEMA_signal_1591, new_AGEMA_signal_1590, n2489}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2645 ( .a ({new_AGEMA_signal_5871, new_AGEMA_signal_5869, new_AGEMA_signal_5867}), .b ({new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2492}), .clk ( clk ), .r ({Fresh[1175], Fresh[1174], Fresh[1173]}), .c ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, n2497}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2646 ( .a ({new_AGEMA_signal_5877, new_AGEMA_signal_5875, new_AGEMA_signal_5873}), .b ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2700}), .clk ( clk ), .r ({Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, n2495}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2647 ( .a ({new_AGEMA_signal_5715, new_AGEMA_signal_5713, new_AGEMA_signal_5711}), .b ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, n2625}), .clk ( clk ), .r ({Fresh[1181], Fresh[1180], Fresh[1179]}), .c ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, n2494}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2650 ( .a ({new_AGEMA_signal_1213, new_AGEMA_signal_1212, n2498}), .b ({new_AGEMA_signal_5541, new_AGEMA_signal_5539, new_AGEMA_signal_5537}), .clk ( clk ), .r ({Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, n2499}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2653 ( .a ({new_AGEMA_signal_5541, new_AGEMA_signal_5539, new_AGEMA_signal_5537}), .b ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, n2674}), .clk ( clk ), .r ({Fresh[1187], Fresh[1186], Fresh[1185]}), .c ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, n2503}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) U2655 ( .s ({new_AGEMA_signal_5721, new_AGEMA_signal_5719, new_AGEMA_signal_5717}), .b ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, n2505}), .a ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2651}), .clk ( clk ), .r ({Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, n2506}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2662 ( .a ({new_AGEMA_signal_1341, new_AGEMA_signal_1340, n2662}), .b ({new_AGEMA_signal_5607, new_AGEMA_signal_5605, new_AGEMA_signal_5603}), .clk ( clk ), .r ({Fresh[1193], Fresh[1192], Fresh[1191]}), .c ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, n2518}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2663 ( .a ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, n2720}), .b ({new_AGEMA_signal_5649, new_AGEMA_signal_5647, new_AGEMA_signal_5645}), .clk ( clk ), .r ({Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, n2517}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2666 ( .a ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, n2520}), .b ({new_AGEMA_signal_5751, new_AGEMA_signal_5749, new_AGEMA_signal_5747}), .clk ( clk ), .r ({Fresh[1199], Fresh[1198], Fresh[1197]}), .c ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, n2523}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2668 ( .a ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, n2774}), .b ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, n2521}), .clk ( clk ), .r ({Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, n2522}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2675 ( .a ({new_AGEMA_signal_5607, new_AGEMA_signal_5605, new_AGEMA_signal_5603}), .b ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, n2531}), .clk ( clk ), .r ({Fresh[1205], Fresh[1204], Fresh[1203]}), .c ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, n2532}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2677 ( .a ({new_AGEMA_signal_5511, new_AGEMA_signal_5509, new_AGEMA_signal_5507}), .b ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, n2533}), .clk ( clk ), .r ({Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, n2534}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2681 ( .a ({new_AGEMA_signal_5883, new_AGEMA_signal_5881, new_AGEMA_signal_5879}), .b ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, n2540}), .clk ( clk ), .r ({Fresh[1211], Fresh[1210], Fresh[1209]}), .c ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, n2542}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2683 ( .a ({new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2545}), .b ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, n2544}), .clk ( clk ), .r ({Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, n2546}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2687 ( .a ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, n2673}), .b ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, n2732}), .clk ( clk ), .r ({Fresh[1217], Fresh[1216], Fresh[1215]}), .c ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, n2551}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2690 ( .a ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, n2553}), .b ({new_AGEMA_signal_5889, new_AGEMA_signal_5887, new_AGEMA_signal_5885}), .clk ( clk ), .r ({Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, n2558}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2692 ( .a ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, n2555}), .b ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, n2554}), .clk ( clk ), .r ({Fresh[1223], Fresh[1222], Fresh[1221]}), .c ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, n2556}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2696 ( .a ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, n2561}), .b ({new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2560}), .clk ( clk ), .r ({Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, n2566}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2697 ( .a ({new_AGEMA_signal_5895, new_AGEMA_signal_5893, new_AGEMA_signal_5891}), .b ({new_AGEMA_signal_1431, new_AGEMA_signal_1430, n2562}), .clk ( clk ), .r ({Fresh[1229], Fresh[1228], Fresh[1227]}), .c ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, n2715}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2703 ( .a ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, n2572}), .b ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, n2571}), .clk ( clk ), .r ({Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, n2573}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2705 ( .a ({new_AGEMA_signal_5847, new_AGEMA_signal_5845, new_AGEMA_signal_5843}), .b ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, n2754}), .clk ( clk ), .r ({Fresh[1235], Fresh[1234], Fresh[1233]}), .c ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, n2585}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2706 ( .a ({new_AGEMA_signal_5781, new_AGEMA_signal_5779, new_AGEMA_signal_5777}), .b ({new_AGEMA_signal_1155, new_AGEMA_signal_1154, n2627}), .clk ( clk ), .r ({Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({new_AGEMA_signal_1611, new_AGEMA_signal_1610, n2581}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2707 ( .a ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, n2575}), .b ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2817}), .clk ( clk ), .r ({Fresh[1241], Fresh[1240], Fresh[1239]}), .c ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, n2579}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2708 ( .a ({new_AGEMA_signal_5877, new_AGEMA_signal_5875, new_AGEMA_signal_5873}), .b ({new_AGEMA_signal_1233, new_AGEMA_signal_1232, n2576}), .clk ( clk ), .r ({Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, n2578}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2711 ( .a ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, n2625}), .b ({new_AGEMA_signal_5757, new_AGEMA_signal_5755, new_AGEMA_signal_5753}), .clk ( clk ), .r ({Fresh[1247], Fresh[1246], Fresh[1245]}), .c ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, n2582}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2715 ( .a ({new_AGEMA_signal_5565, new_AGEMA_signal_5563, new_AGEMA_signal_5561}), .b ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, n2586}), .clk ( clk ), .r ({Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, n2588}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2719 ( .a ({new_AGEMA_signal_1269, new_AGEMA_signal_1268, n2594}), .b ({new_AGEMA_signal_5847, new_AGEMA_signal_5845, new_AGEMA_signal_5843}), .clk ( clk ), .r ({Fresh[1253], Fresh[1252], Fresh[1251]}), .c ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, n2607}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2722 ( .a ({new_AGEMA_signal_1293, new_AGEMA_signal_1292, n2597}), .b ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, n2596}), .clk ( clk ), .r ({Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, n2605}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2724 ( .a ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, n2598}), .b ({new_AGEMA_signal_5901, new_AGEMA_signal_5899, new_AGEMA_signal_5897}), .clk ( clk ), .r ({Fresh[1259], Fresh[1258], Fresh[1257]}), .c ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, n2603}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2726 ( .a ({new_AGEMA_signal_1101, new_AGEMA_signal_1100, n2599}), .b ({new_AGEMA_signal_5775, new_AGEMA_signal_5773, new_AGEMA_signal_5771}), .clk ( clk ), .r ({Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, n2601}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2733 ( .a ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, n2610}), .b ({new_AGEMA_signal_5751, new_AGEMA_signal_5749, new_AGEMA_signal_5747}), .clk ( clk ), .r ({Fresh[1265], Fresh[1264], Fresh[1263]}), .c ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, n2620}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2736 ( .a ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, n2614}), .b ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, n2613}), .clk ( clk ), .r ({Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, n2618}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2743 ( .a ({new_AGEMA_signal_5721, new_AGEMA_signal_5719, new_AGEMA_signal_5717}), .b ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, n2625}), .clk ( clk ), .r ({Fresh[1271], Fresh[1270], Fresh[1269]}), .c ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, n2626}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2746 ( .a ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, n2631}), .b ({new_AGEMA_signal_5649, new_AGEMA_signal_5647, new_AGEMA_signal_5645}), .clk ( clk ), .r ({Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, n2632}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2752 ( .a ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, n2784}), .b ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, n2642}), .clk ( clk ), .r ({Fresh[1277], Fresh[1276], Fresh[1275]}), .c ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, n2644}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2754 ( .a ({new_AGEMA_signal_5535, new_AGEMA_signal_5533, new_AGEMA_signal_5531}), .b ({new_AGEMA_signal_1245, new_AGEMA_signal_1244, n2645}), .clk ( clk ), .r ({Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, n2646}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2758 ( .a ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2651}), .b ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, n2650}), .clk ( clk ), .r ({Fresh[1283], Fresh[1282], Fresh[1281]}), .c ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, n2653}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2760 ( .a ({new_AGEMA_signal_5775, new_AGEMA_signal_5773, new_AGEMA_signal_5771}), .b ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, n2654}), .clk ( clk ), .r ({Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, n2655}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2764 ( .a ({new_AGEMA_signal_1341, new_AGEMA_signal_1340, n2662}), .b ({new_AGEMA_signal_5787, new_AGEMA_signal_5785, new_AGEMA_signal_5783}), .clk ( clk ), .r ({Fresh[1289], Fresh[1288], Fresh[1287]}), .c ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, n2663}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2770 ( .a ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, n2673}), .b ({new_AGEMA_signal_5757, new_AGEMA_signal_5755, new_AGEMA_signal_5753}), .clk ( clk ), .r ({Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, n2675}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2772 ( .a ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, n2677}), .b ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, n2676}), .clk ( clk ), .r ({Fresh[1295], Fresh[1294], Fresh[1293]}), .c ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, n2678}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2780 ( .a ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, n2690}), .b ({new_AGEMA_signal_5781, new_AGEMA_signal_5779, new_AGEMA_signal_5777}), .clk ( clk ), .r ({Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, n2691}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2782 ( .a ({new_AGEMA_signal_5799, new_AGEMA_signal_5797, new_AGEMA_signal_5795}), .b ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, n2693}), .clk ( clk ), .r ({Fresh[1301], Fresh[1300], Fresh[1299]}), .c ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, n2695}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2785 ( .a ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2700}), .b ({new_AGEMA_signal_5895, new_AGEMA_signal_5893, new_AGEMA_signal_5891}), .clk ( clk ), .r ({Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, n2701}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2791 ( .a ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, n2711}), .b ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, n2710}), .clk ( clk ), .r ({Fresh[1307], Fresh[1306], Fresh[1305]}), .c ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, n2717}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2796 ( .a ({new_AGEMA_signal_1705, new_AGEMA_signal_1704, n2720}), .b ({new_AGEMA_signal_5721, new_AGEMA_signal_5719, new_AGEMA_signal_5717}), .clk ( clk ), .r ({Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, n2729}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2798 ( .a ({new_AGEMA_signal_5619, new_AGEMA_signal_5617, new_AGEMA_signal_5615}), .b ({new_AGEMA_signal_1305, new_AGEMA_signal_1304, n2722}), .clk ( clk ), .r ({Fresh[1313], Fresh[1312], Fresh[1311]}), .c ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, n2727}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2803 ( .a ({new_AGEMA_signal_1329, new_AGEMA_signal_1328, n2732}), .b ({new_AGEMA_signal_1419, new_AGEMA_signal_1418, n2731}), .clk ( clk ), .r ({Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, n2733}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2807 ( .a ({new_AGEMA_signal_5907, new_AGEMA_signal_5905, new_AGEMA_signal_5903}), .b ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, n2738}), .clk ( clk ), .r ({Fresh[1319], Fresh[1318], Fresh[1317]}), .c ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, n2740}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2812 ( .a ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, n2748}), .b ({new_AGEMA_signal_5511, new_AGEMA_signal_5509, new_AGEMA_signal_5507}), .clk ( clk ), .r ({Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, n2749}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2815 ( .a ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, n2754}), .b ({new_AGEMA_signal_5631, new_AGEMA_signal_5629, new_AGEMA_signal_5627}), .clk ( clk ), .r ({Fresh[1325], Fresh[1324], Fresh[1323]}), .c ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, n2757}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2816 ( .a ({new_AGEMA_signal_1119, new_AGEMA_signal_1118, n2755}), .b ({new_AGEMA_signal_5913, new_AGEMA_signal_5911, new_AGEMA_signal_5909}), .clk ( clk ), .r ({Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, n2756}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2819 ( .a ({new_AGEMA_signal_1347, new_AGEMA_signal_1346, n2761}), .b ({new_AGEMA_signal_5805, new_AGEMA_signal_5803, new_AGEMA_signal_5801}), .clk ( clk ), .r ({Fresh[1331], Fresh[1330], Fresh[1329]}), .c ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, n2762}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2823 ( .a ({new_AGEMA_signal_5511, new_AGEMA_signal_5509, new_AGEMA_signal_5507}), .b ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, n2768}), .clk ( clk ), .r ({Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, n2770}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2825 ( .a ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, n2773}), .b ({new_AGEMA_signal_5913, new_AGEMA_signal_5911, new_AGEMA_signal_5909}), .clk ( clk ), .r ({Fresh[1337], Fresh[1336], Fresh[1335]}), .c ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, n2776}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2826 ( .a ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, n2774}), .b ({new_AGEMA_signal_5517, new_AGEMA_signal_5515, new_AGEMA_signal_5513}), .clk ( clk ), .r ({Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, n2775}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2830 ( .a ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, n2782}), .b ({new_AGEMA_signal_1309, new_AGEMA_signal_1308, n2781}), .clk ( clk ), .r ({Fresh[1343], Fresh[1342], Fresh[1341]}), .c ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, n2783}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2836 ( .a ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, n2794}), .b ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, n2793}), .clk ( clk ), .r ({Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, n2795}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2845 ( .a ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, n2812}), .b ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, n2811}), .clk ( clk ), .r ({Fresh[1349], Fresh[1348], Fresh[1347]}), .c ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, n2814}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2848 ( .a ({new_AGEMA_signal_5583, new_AGEMA_signal_5581, new_AGEMA_signal_5579}), .b ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2817}), .clk ( clk ), .r ({Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, n2819}) ) ;
    buf_clk new_AGEMA_reg_buffer_1426 ( .C ( clk ), .D ( new_AGEMA_signal_5914 ), .Q ( new_AGEMA_signal_5915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1428 ( .C ( clk ), .D ( new_AGEMA_signal_5916 ), .Q ( new_AGEMA_signal_5917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1430 ( .C ( clk ), .D ( new_AGEMA_signal_5918 ), .Q ( new_AGEMA_signal_5919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1432 ( .C ( clk ), .D ( new_AGEMA_signal_5920 ), .Q ( new_AGEMA_signal_5921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1434 ( .C ( clk ), .D ( new_AGEMA_signal_5922 ), .Q ( new_AGEMA_signal_5923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1436 ( .C ( clk ), .D ( new_AGEMA_signal_5924 ), .Q ( new_AGEMA_signal_5925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1440 ( .C ( clk ), .D ( new_AGEMA_signal_5928 ), .Q ( new_AGEMA_signal_5929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1444 ( .C ( clk ), .D ( new_AGEMA_signal_5932 ), .Q ( new_AGEMA_signal_5933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1448 ( .C ( clk ), .D ( new_AGEMA_signal_5936 ), .Q ( new_AGEMA_signal_5937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1450 ( .C ( clk ), .D ( new_AGEMA_signal_5938 ), .Q ( new_AGEMA_signal_5939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1452 ( .C ( clk ), .D ( new_AGEMA_signal_5940 ), .Q ( new_AGEMA_signal_5941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1454 ( .C ( clk ), .D ( new_AGEMA_signal_5942 ), .Q ( new_AGEMA_signal_5943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1456 ( .C ( clk ), .D ( new_AGEMA_signal_5944 ), .Q ( new_AGEMA_signal_5945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1458 ( .C ( clk ), .D ( new_AGEMA_signal_5946 ), .Q ( new_AGEMA_signal_5947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1460 ( .C ( clk ), .D ( new_AGEMA_signal_5948 ), .Q ( new_AGEMA_signal_5949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1462 ( .C ( clk ), .D ( new_AGEMA_signal_5950 ), .Q ( new_AGEMA_signal_5951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1464 ( .C ( clk ), .D ( new_AGEMA_signal_5952 ), .Q ( new_AGEMA_signal_5953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1466 ( .C ( clk ), .D ( new_AGEMA_signal_5954 ), .Q ( new_AGEMA_signal_5955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1468 ( .C ( clk ), .D ( new_AGEMA_signal_5956 ), .Q ( new_AGEMA_signal_5957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1470 ( .C ( clk ), .D ( new_AGEMA_signal_5958 ), .Q ( new_AGEMA_signal_5959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1472 ( .C ( clk ), .D ( new_AGEMA_signal_5960 ), .Q ( new_AGEMA_signal_5961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1474 ( .C ( clk ), .D ( new_AGEMA_signal_5962 ), .Q ( new_AGEMA_signal_5963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1476 ( .C ( clk ), .D ( new_AGEMA_signal_5964 ), .Q ( new_AGEMA_signal_5965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1478 ( .C ( clk ), .D ( new_AGEMA_signal_5966 ), .Q ( new_AGEMA_signal_5967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1480 ( .C ( clk ), .D ( new_AGEMA_signal_5968 ), .Q ( new_AGEMA_signal_5969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1482 ( .C ( clk ), .D ( new_AGEMA_signal_5970 ), .Q ( new_AGEMA_signal_5971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1484 ( .C ( clk ), .D ( new_AGEMA_signal_5972 ), .Q ( new_AGEMA_signal_5973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1486 ( .C ( clk ), .D ( new_AGEMA_signal_5974 ), .Q ( new_AGEMA_signal_5975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1488 ( .C ( clk ), .D ( new_AGEMA_signal_5976 ), .Q ( new_AGEMA_signal_5977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1490 ( .C ( clk ), .D ( new_AGEMA_signal_5978 ), .Q ( new_AGEMA_signal_5979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1492 ( .C ( clk ), .D ( new_AGEMA_signal_5980 ), .Q ( new_AGEMA_signal_5981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1494 ( .C ( clk ), .D ( new_AGEMA_signal_5982 ), .Q ( new_AGEMA_signal_5983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1496 ( .C ( clk ), .D ( new_AGEMA_signal_5984 ), .Q ( new_AGEMA_signal_5985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1498 ( .C ( clk ), .D ( new_AGEMA_signal_5986 ), .Q ( new_AGEMA_signal_5987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1500 ( .C ( clk ), .D ( new_AGEMA_signal_5988 ), .Q ( new_AGEMA_signal_5989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1502 ( .C ( clk ), .D ( new_AGEMA_signal_5990 ), .Q ( new_AGEMA_signal_5991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1504 ( .C ( clk ), .D ( new_AGEMA_signal_5992 ), .Q ( new_AGEMA_signal_5993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1506 ( .C ( clk ), .D ( new_AGEMA_signal_5994 ), .Q ( new_AGEMA_signal_5995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1508 ( .C ( clk ), .D ( new_AGEMA_signal_5996 ), .Q ( new_AGEMA_signal_5997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1510 ( .C ( clk ), .D ( new_AGEMA_signal_5998 ), .Q ( new_AGEMA_signal_5999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1512 ( .C ( clk ), .D ( new_AGEMA_signal_6000 ), .Q ( new_AGEMA_signal_6001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1514 ( .C ( clk ), .D ( new_AGEMA_signal_6002 ), .Q ( new_AGEMA_signal_6003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1518 ( .C ( clk ), .D ( new_AGEMA_signal_6006 ), .Q ( new_AGEMA_signal_6007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1522 ( .C ( clk ), .D ( new_AGEMA_signal_6010 ), .Q ( new_AGEMA_signal_6011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1526 ( .C ( clk ), .D ( new_AGEMA_signal_6014 ), .Q ( new_AGEMA_signal_6015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1528 ( .C ( clk ), .D ( new_AGEMA_signal_6016 ), .Q ( new_AGEMA_signal_6017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1530 ( .C ( clk ), .D ( new_AGEMA_signal_6018 ), .Q ( new_AGEMA_signal_6019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1532 ( .C ( clk ), .D ( new_AGEMA_signal_6020 ), .Q ( new_AGEMA_signal_6021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1534 ( .C ( clk ), .D ( new_AGEMA_signal_6022 ), .Q ( new_AGEMA_signal_6023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1536 ( .C ( clk ), .D ( new_AGEMA_signal_6024 ), .Q ( new_AGEMA_signal_6025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1538 ( .C ( clk ), .D ( new_AGEMA_signal_6026 ), .Q ( new_AGEMA_signal_6027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1540 ( .C ( clk ), .D ( new_AGEMA_signal_6028 ), .Q ( new_AGEMA_signal_6029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1542 ( .C ( clk ), .D ( new_AGEMA_signal_6030 ), .Q ( new_AGEMA_signal_6031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1544 ( .C ( clk ), .D ( new_AGEMA_signal_6032 ), .Q ( new_AGEMA_signal_6033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1546 ( .C ( clk ), .D ( new_AGEMA_signal_6034 ), .Q ( new_AGEMA_signal_6035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1548 ( .C ( clk ), .D ( new_AGEMA_signal_6036 ), .Q ( new_AGEMA_signal_6037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1550 ( .C ( clk ), .D ( new_AGEMA_signal_6038 ), .Q ( new_AGEMA_signal_6039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1552 ( .C ( clk ), .D ( new_AGEMA_signal_6040 ), .Q ( new_AGEMA_signal_6041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1554 ( .C ( clk ), .D ( new_AGEMA_signal_6042 ), .Q ( new_AGEMA_signal_6043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1556 ( .C ( clk ), .D ( new_AGEMA_signal_6044 ), .Q ( new_AGEMA_signal_6045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1558 ( .C ( clk ), .D ( new_AGEMA_signal_6046 ), .Q ( new_AGEMA_signal_6047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1560 ( .C ( clk ), .D ( new_AGEMA_signal_6048 ), .Q ( new_AGEMA_signal_6049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1562 ( .C ( clk ), .D ( new_AGEMA_signal_6050 ), .Q ( new_AGEMA_signal_6051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1564 ( .C ( clk ), .D ( new_AGEMA_signal_6052 ), .Q ( new_AGEMA_signal_6053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1566 ( .C ( clk ), .D ( new_AGEMA_signal_6054 ), .Q ( new_AGEMA_signal_6055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1568 ( .C ( clk ), .D ( new_AGEMA_signal_6056 ), .Q ( new_AGEMA_signal_6057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1572 ( .C ( clk ), .D ( new_AGEMA_signal_6060 ), .Q ( new_AGEMA_signal_6061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1576 ( .C ( clk ), .D ( new_AGEMA_signal_6064 ), .Q ( new_AGEMA_signal_6065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1580 ( .C ( clk ), .D ( new_AGEMA_signal_6068 ), .Q ( new_AGEMA_signal_6069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1582 ( .C ( clk ), .D ( new_AGEMA_signal_6070 ), .Q ( new_AGEMA_signal_6071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1584 ( .C ( clk ), .D ( new_AGEMA_signal_6072 ), .Q ( new_AGEMA_signal_6073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1586 ( .C ( clk ), .D ( new_AGEMA_signal_6074 ), .Q ( new_AGEMA_signal_6075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1588 ( .C ( clk ), .D ( new_AGEMA_signal_6076 ), .Q ( new_AGEMA_signal_6077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1590 ( .C ( clk ), .D ( new_AGEMA_signal_6078 ), .Q ( new_AGEMA_signal_6079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1592 ( .C ( clk ), .D ( new_AGEMA_signal_6080 ), .Q ( new_AGEMA_signal_6081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1594 ( .C ( clk ), .D ( new_AGEMA_signal_6082 ), .Q ( new_AGEMA_signal_6083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1596 ( .C ( clk ), .D ( new_AGEMA_signal_6084 ), .Q ( new_AGEMA_signal_6085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1598 ( .C ( clk ), .D ( new_AGEMA_signal_6086 ), .Q ( new_AGEMA_signal_6087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1600 ( .C ( clk ), .D ( new_AGEMA_signal_6088 ), .Q ( new_AGEMA_signal_6089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1602 ( .C ( clk ), .D ( new_AGEMA_signal_6090 ), .Q ( new_AGEMA_signal_6091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1604 ( .C ( clk ), .D ( new_AGEMA_signal_6092 ), .Q ( new_AGEMA_signal_6093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1606 ( .C ( clk ), .D ( new_AGEMA_signal_6094 ), .Q ( new_AGEMA_signal_6095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1608 ( .C ( clk ), .D ( new_AGEMA_signal_6096 ), .Q ( new_AGEMA_signal_6097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1610 ( .C ( clk ), .D ( new_AGEMA_signal_6098 ), .Q ( new_AGEMA_signal_6099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1614 ( .C ( clk ), .D ( new_AGEMA_signal_6102 ), .Q ( new_AGEMA_signal_6103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1618 ( .C ( clk ), .D ( new_AGEMA_signal_6106 ), .Q ( new_AGEMA_signal_6107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1622 ( .C ( clk ), .D ( new_AGEMA_signal_6110 ), .Q ( new_AGEMA_signal_6111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1624 ( .C ( clk ), .D ( new_AGEMA_signal_6112 ), .Q ( new_AGEMA_signal_6113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1626 ( .C ( clk ), .D ( new_AGEMA_signal_6114 ), .Q ( new_AGEMA_signal_6115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1628 ( .C ( clk ), .D ( new_AGEMA_signal_6116 ), .Q ( new_AGEMA_signal_6117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1630 ( .C ( clk ), .D ( new_AGEMA_signal_6118 ), .Q ( new_AGEMA_signal_6119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1632 ( .C ( clk ), .D ( new_AGEMA_signal_6120 ), .Q ( new_AGEMA_signal_6121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1634 ( .C ( clk ), .D ( new_AGEMA_signal_6122 ), .Q ( new_AGEMA_signal_6123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1636 ( .C ( clk ), .D ( new_AGEMA_signal_6124 ), .Q ( new_AGEMA_signal_6125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1638 ( .C ( clk ), .D ( new_AGEMA_signal_6126 ), .Q ( new_AGEMA_signal_6127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1640 ( .C ( clk ), .D ( new_AGEMA_signal_6128 ), .Q ( new_AGEMA_signal_6129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1644 ( .C ( clk ), .D ( new_AGEMA_signal_6132 ), .Q ( new_AGEMA_signal_6133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1648 ( .C ( clk ), .D ( new_AGEMA_signal_6136 ), .Q ( new_AGEMA_signal_6137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1652 ( .C ( clk ), .D ( new_AGEMA_signal_6140 ), .Q ( new_AGEMA_signal_6141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1654 ( .C ( clk ), .D ( new_AGEMA_signal_6142 ), .Q ( new_AGEMA_signal_6143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1656 ( .C ( clk ), .D ( new_AGEMA_signal_6144 ), .Q ( new_AGEMA_signal_6145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1658 ( .C ( clk ), .D ( new_AGEMA_signal_6146 ), .Q ( new_AGEMA_signal_6147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1660 ( .C ( clk ), .D ( new_AGEMA_signal_6148 ), .Q ( new_AGEMA_signal_6149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1662 ( .C ( clk ), .D ( new_AGEMA_signal_6150 ), .Q ( new_AGEMA_signal_6151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1664 ( .C ( clk ), .D ( new_AGEMA_signal_6152 ), .Q ( new_AGEMA_signal_6153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1666 ( .C ( clk ), .D ( new_AGEMA_signal_6154 ), .Q ( new_AGEMA_signal_6155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1668 ( .C ( clk ), .D ( new_AGEMA_signal_6156 ), .Q ( new_AGEMA_signal_6157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1670 ( .C ( clk ), .D ( new_AGEMA_signal_6158 ), .Q ( new_AGEMA_signal_6159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1674 ( .C ( clk ), .D ( new_AGEMA_signal_6162 ), .Q ( new_AGEMA_signal_6163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1678 ( .C ( clk ), .D ( new_AGEMA_signal_6166 ), .Q ( new_AGEMA_signal_6167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1682 ( .C ( clk ), .D ( new_AGEMA_signal_6170 ), .Q ( new_AGEMA_signal_6171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1684 ( .C ( clk ), .D ( new_AGEMA_signal_6172 ), .Q ( new_AGEMA_signal_6173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1686 ( .C ( clk ), .D ( new_AGEMA_signal_6174 ), .Q ( new_AGEMA_signal_6175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1688 ( .C ( clk ), .D ( new_AGEMA_signal_6176 ), .Q ( new_AGEMA_signal_6177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1690 ( .C ( clk ), .D ( new_AGEMA_signal_6178 ), .Q ( new_AGEMA_signal_6179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1692 ( .C ( clk ), .D ( new_AGEMA_signal_6180 ), .Q ( new_AGEMA_signal_6181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1694 ( .C ( clk ), .D ( new_AGEMA_signal_6182 ), .Q ( new_AGEMA_signal_6183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1696 ( .C ( clk ), .D ( new_AGEMA_signal_6184 ), .Q ( new_AGEMA_signal_6185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1698 ( .C ( clk ), .D ( new_AGEMA_signal_6186 ), .Q ( new_AGEMA_signal_6187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1700 ( .C ( clk ), .D ( new_AGEMA_signal_6188 ), .Q ( new_AGEMA_signal_6189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1702 ( .C ( clk ), .D ( new_AGEMA_signal_6190 ), .Q ( new_AGEMA_signal_6191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1704 ( .C ( clk ), .D ( new_AGEMA_signal_6192 ), .Q ( new_AGEMA_signal_6193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1706 ( .C ( clk ), .D ( new_AGEMA_signal_6194 ), .Q ( new_AGEMA_signal_6195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1708 ( .C ( clk ), .D ( new_AGEMA_signal_6196 ), .Q ( new_AGEMA_signal_6197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1710 ( .C ( clk ), .D ( new_AGEMA_signal_6198 ), .Q ( new_AGEMA_signal_6199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1712 ( .C ( clk ), .D ( new_AGEMA_signal_6200 ), .Q ( new_AGEMA_signal_6201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C ( clk ), .D ( new_AGEMA_signal_6202 ), .Q ( new_AGEMA_signal_6203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C ( clk ), .D ( new_AGEMA_signal_6204 ), .Q ( new_AGEMA_signal_6205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C ( clk ), .D ( new_AGEMA_signal_6206 ), .Q ( new_AGEMA_signal_6207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C ( clk ), .D ( new_AGEMA_signal_6208 ), .Q ( new_AGEMA_signal_6209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C ( clk ), .D ( new_AGEMA_signal_6210 ), .Q ( new_AGEMA_signal_6211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C ( clk ), .D ( new_AGEMA_signal_6212 ), .Q ( new_AGEMA_signal_6213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C ( clk ), .D ( new_AGEMA_signal_6214 ), .Q ( new_AGEMA_signal_6215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C ( clk ), .D ( new_AGEMA_signal_6216 ), .Q ( new_AGEMA_signal_6217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C ( clk ), .D ( new_AGEMA_signal_6218 ), .Q ( new_AGEMA_signal_6219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C ( clk ), .D ( new_AGEMA_signal_6220 ), .Q ( new_AGEMA_signal_6221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C ( clk ), .D ( new_AGEMA_signal_6222 ), .Q ( new_AGEMA_signal_6223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C ( clk ), .D ( new_AGEMA_signal_6224 ), .Q ( new_AGEMA_signal_6225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C ( clk ), .D ( new_AGEMA_signal_6226 ), .Q ( new_AGEMA_signal_6227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C ( clk ), .D ( new_AGEMA_signal_6228 ), .Q ( new_AGEMA_signal_6229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C ( clk ), .D ( new_AGEMA_signal_6230 ), .Q ( new_AGEMA_signal_6231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C ( clk ), .D ( new_AGEMA_signal_6232 ), .Q ( new_AGEMA_signal_6233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C ( clk ), .D ( new_AGEMA_signal_6234 ), .Q ( new_AGEMA_signal_6235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C ( clk ), .D ( new_AGEMA_signal_6236 ), .Q ( new_AGEMA_signal_6237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C ( clk ), .D ( new_AGEMA_signal_6238 ), .Q ( new_AGEMA_signal_6239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C ( clk ), .D ( new_AGEMA_signal_6240 ), .Q ( new_AGEMA_signal_6241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C ( clk ), .D ( new_AGEMA_signal_6242 ), .Q ( new_AGEMA_signal_6243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C ( clk ), .D ( new_AGEMA_signal_6244 ), .Q ( new_AGEMA_signal_6245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C ( clk ), .D ( new_AGEMA_signal_6246 ), .Q ( new_AGEMA_signal_6247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C ( clk ), .D ( new_AGEMA_signal_6248 ), .Q ( new_AGEMA_signal_6249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C ( clk ), .D ( new_AGEMA_signal_6250 ), .Q ( new_AGEMA_signal_6251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C ( clk ), .D ( new_AGEMA_signal_6252 ), .Q ( new_AGEMA_signal_6253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C ( clk ), .D ( new_AGEMA_signal_6254 ), .Q ( new_AGEMA_signal_6255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C ( clk ), .D ( new_AGEMA_signal_6256 ), .Q ( new_AGEMA_signal_6257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C ( clk ), .D ( new_AGEMA_signal_6258 ), .Q ( new_AGEMA_signal_6259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C ( clk ), .D ( new_AGEMA_signal_6260 ), .Q ( new_AGEMA_signal_6261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C ( clk ), .D ( new_AGEMA_signal_6262 ), .Q ( new_AGEMA_signal_6263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C ( clk ), .D ( new_AGEMA_signal_6264 ), .Q ( new_AGEMA_signal_6265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C ( clk ), .D ( new_AGEMA_signal_6266 ), .Q ( new_AGEMA_signal_6267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C ( clk ), .D ( new_AGEMA_signal_6268 ), .Q ( new_AGEMA_signal_6269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C ( clk ), .D ( new_AGEMA_signal_6270 ), .Q ( new_AGEMA_signal_6271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C ( clk ), .D ( new_AGEMA_signal_6272 ), .Q ( new_AGEMA_signal_6273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C ( clk ), .D ( new_AGEMA_signal_6278 ), .Q ( new_AGEMA_signal_6279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C ( clk ), .D ( new_AGEMA_signal_6284 ), .Q ( new_AGEMA_signal_6285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C ( clk ), .D ( new_AGEMA_signal_6290 ), .Q ( new_AGEMA_signal_6291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C ( clk ), .D ( new_AGEMA_signal_6292 ), .Q ( new_AGEMA_signal_6293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C ( clk ), .D ( new_AGEMA_signal_6294 ), .Q ( new_AGEMA_signal_6295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C ( clk ), .D ( new_AGEMA_signal_6296 ), .Q ( new_AGEMA_signal_6297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C ( clk ), .D ( new_AGEMA_signal_6298 ), .Q ( new_AGEMA_signal_6299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C ( clk ), .D ( new_AGEMA_signal_6300 ), .Q ( new_AGEMA_signal_6301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C ( clk ), .D ( new_AGEMA_signal_6302 ), .Q ( new_AGEMA_signal_6303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C ( clk ), .D ( new_AGEMA_signal_6304 ), .Q ( new_AGEMA_signal_6305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C ( clk ), .D ( new_AGEMA_signal_6306 ), .Q ( new_AGEMA_signal_6307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C ( clk ), .D ( new_AGEMA_signal_6308 ), .Q ( new_AGEMA_signal_6309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C ( clk ), .D ( new_AGEMA_signal_6312 ), .Q ( new_AGEMA_signal_6313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C ( clk ), .D ( new_AGEMA_signal_6316 ), .Q ( new_AGEMA_signal_6317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C ( clk ), .D ( new_AGEMA_signal_6320 ), .Q ( new_AGEMA_signal_6321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C ( clk ), .D ( new_AGEMA_signal_6322 ), .Q ( new_AGEMA_signal_6323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C ( clk ), .D ( new_AGEMA_signal_6324 ), .Q ( new_AGEMA_signal_6325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C ( clk ), .D ( new_AGEMA_signal_6326 ), .Q ( new_AGEMA_signal_6327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C ( clk ), .D ( new_AGEMA_signal_6328 ), .Q ( new_AGEMA_signal_6329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C ( clk ), .D ( new_AGEMA_signal_6330 ), .Q ( new_AGEMA_signal_6331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C ( clk ), .D ( new_AGEMA_signal_6332 ), .Q ( new_AGEMA_signal_6333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C ( clk ), .D ( new_AGEMA_signal_6334 ), .Q ( new_AGEMA_signal_6335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C ( clk ), .D ( new_AGEMA_signal_6336 ), .Q ( new_AGEMA_signal_6337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C ( clk ), .D ( new_AGEMA_signal_6338 ), .Q ( new_AGEMA_signal_6339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C ( clk ), .D ( new_AGEMA_signal_6342 ), .Q ( new_AGEMA_signal_6343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C ( clk ), .D ( new_AGEMA_signal_6346 ), .Q ( new_AGEMA_signal_6347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C ( clk ), .D ( new_AGEMA_signal_6350 ), .Q ( new_AGEMA_signal_6351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C ( clk ), .D ( new_AGEMA_signal_6352 ), .Q ( new_AGEMA_signal_6353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C ( clk ), .D ( new_AGEMA_signal_6354 ), .Q ( new_AGEMA_signal_6355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C ( clk ), .D ( new_AGEMA_signal_6356 ), .Q ( new_AGEMA_signal_6357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C ( clk ), .D ( new_AGEMA_signal_6358 ), .Q ( new_AGEMA_signal_6359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C ( clk ), .D ( new_AGEMA_signal_6360 ), .Q ( new_AGEMA_signal_6361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C ( clk ), .D ( new_AGEMA_signal_6362 ), .Q ( new_AGEMA_signal_6363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C ( clk ), .D ( new_AGEMA_signal_6364 ), .Q ( new_AGEMA_signal_6365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C ( clk ), .D ( new_AGEMA_signal_6366 ), .Q ( new_AGEMA_signal_6367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C ( clk ), .D ( new_AGEMA_signal_6368 ), .Q ( new_AGEMA_signal_6369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C ( clk ), .D ( new_AGEMA_signal_6370 ), .Q ( new_AGEMA_signal_6371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C ( clk ), .D ( new_AGEMA_signal_6372 ), .Q ( new_AGEMA_signal_6373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C ( clk ), .D ( new_AGEMA_signal_6374 ), .Q ( new_AGEMA_signal_6375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C ( clk ), .D ( new_AGEMA_signal_6376 ), .Q ( new_AGEMA_signal_6377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C ( clk ), .D ( new_AGEMA_signal_6378 ), .Q ( new_AGEMA_signal_6379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C ( clk ), .D ( new_AGEMA_signal_6380 ), .Q ( new_AGEMA_signal_6381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C ( clk ), .D ( new_AGEMA_signal_6382 ), .Q ( new_AGEMA_signal_6383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C ( clk ), .D ( new_AGEMA_signal_6384 ), .Q ( new_AGEMA_signal_6385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C ( clk ), .D ( new_AGEMA_signal_6386 ), .Q ( new_AGEMA_signal_6387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C ( clk ), .D ( new_AGEMA_signal_6388 ), .Q ( new_AGEMA_signal_6389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1902 ( .C ( clk ), .D ( new_AGEMA_signal_6390 ), .Q ( new_AGEMA_signal_6391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C ( clk ), .D ( new_AGEMA_signal_6392 ), .Q ( new_AGEMA_signal_6393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C ( clk ), .D ( new_AGEMA_signal_6396 ), .Q ( new_AGEMA_signal_6397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C ( clk ), .D ( new_AGEMA_signal_6400 ), .Q ( new_AGEMA_signal_6401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C ( clk ), .D ( new_AGEMA_signal_6404 ), .Q ( new_AGEMA_signal_6405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C ( clk ), .D ( new_AGEMA_signal_6406 ), .Q ( new_AGEMA_signal_6407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C ( clk ), .D ( new_AGEMA_signal_6408 ), .Q ( new_AGEMA_signal_6409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C ( clk ), .D ( new_AGEMA_signal_6410 ), .Q ( new_AGEMA_signal_6411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C ( clk ), .D ( new_AGEMA_signal_6412 ), .Q ( new_AGEMA_signal_6413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C ( clk ), .D ( new_AGEMA_signal_6414 ), .Q ( new_AGEMA_signal_6415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C ( clk ), .D ( new_AGEMA_signal_6416 ), .Q ( new_AGEMA_signal_6417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C ( clk ), .D ( new_AGEMA_signal_6420 ), .Q ( new_AGEMA_signal_6421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C ( clk ), .D ( new_AGEMA_signal_6424 ), .Q ( new_AGEMA_signal_6425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C ( clk ), .D ( new_AGEMA_signal_6428 ), .Q ( new_AGEMA_signal_6429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C ( clk ), .D ( new_AGEMA_signal_6430 ), .Q ( new_AGEMA_signal_6431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C ( clk ), .D ( new_AGEMA_signal_6432 ), .Q ( new_AGEMA_signal_6433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C ( clk ), .D ( new_AGEMA_signal_6434 ), .Q ( new_AGEMA_signal_6435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C ( clk ), .D ( new_AGEMA_signal_6436 ), .Q ( new_AGEMA_signal_6437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C ( clk ), .D ( new_AGEMA_signal_6440 ), .Q ( new_AGEMA_signal_6441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C ( clk ), .D ( new_AGEMA_signal_6444 ), .Q ( new_AGEMA_signal_6445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C ( clk ), .D ( new_AGEMA_signal_6448 ), .Q ( new_AGEMA_signal_6449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C ( clk ), .D ( new_AGEMA_signal_6452 ), .Q ( new_AGEMA_signal_6453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C ( clk ), .D ( new_AGEMA_signal_6456 ), .Q ( new_AGEMA_signal_6457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C ( clk ), .D ( new_AGEMA_signal_6472 ), .Q ( new_AGEMA_signal_6473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C ( clk ), .D ( new_AGEMA_signal_6476 ), .Q ( new_AGEMA_signal_6477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C ( clk ), .D ( new_AGEMA_signal_6480 ), .Q ( new_AGEMA_signal_6481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C ( clk ), .D ( new_AGEMA_signal_6490 ), .Q ( new_AGEMA_signal_6491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C ( clk ), .D ( new_AGEMA_signal_6494 ), .Q ( new_AGEMA_signal_6495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C ( clk ), .D ( new_AGEMA_signal_6498 ), .Q ( new_AGEMA_signal_6499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C ( clk ), .D ( new_AGEMA_signal_6508 ), .Q ( new_AGEMA_signal_6509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C ( clk ), .D ( new_AGEMA_signal_6512 ), .Q ( new_AGEMA_signal_6513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C ( clk ), .D ( new_AGEMA_signal_6516 ), .Q ( new_AGEMA_signal_6517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C ( clk ), .D ( new_AGEMA_signal_6520 ), .Q ( new_AGEMA_signal_6521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C ( clk ), .D ( new_AGEMA_signal_6524 ), .Q ( new_AGEMA_signal_6525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C ( clk ), .D ( new_AGEMA_signal_6528 ), .Q ( new_AGEMA_signal_6529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C ( clk ), .D ( new_AGEMA_signal_6556 ), .Q ( new_AGEMA_signal_6557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C ( clk ), .D ( new_AGEMA_signal_6560 ), .Q ( new_AGEMA_signal_6561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C ( clk ), .D ( new_AGEMA_signal_6564 ), .Q ( new_AGEMA_signal_6565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C ( clk ), .D ( new_AGEMA_signal_6568 ), .Q ( new_AGEMA_signal_6569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C ( clk ), .D ( new_AGEMA_signal_6572 ), .Q ( new_AGEMA_signal_6573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C ( clk ), .D ( new_AGEMA_signal_6576 ), .Q ( new_AGEMA_signal_6577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C ( clk ), .D ( new_AGEMA_signal_6580 ), .Q ( new_AGEMA_signal_6581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C ( clk ), .D ( new_AGEMA_signal_6584 ), .Q ( new_AGEMA_signal_6585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C ( clk ), .D ( new_AGEMA_signal_6588 ), .Q ( new_AGEMA_signal_6589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C ( clk ), .D ( new_AGEMA_signal_6610 ), .Q ( new_AGEMA_signal_6611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C ( clk ), .D ( new_AGEMA_signal_6614 ), .Q ( new_AGEMA_signal_6615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C ( clk ), .D ( new_AGEMA_signal_6618 ), .Q ( new_AGEMA_signal_6619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C ( clk ), .D ( new_AGEMA_signal_6628 ), .Q ( new_AGEMA_signal_6629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2144 ( .C ( clk ), .D ( new_AGEMA_signal_6632 ), .Q ( new_AGEMA_signal_6633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2148 ( .C ( clk ), .D ( new_AGEMA_signal_6636 ), .Q ( new_AGEMA_signal_6637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2154 ( .C ( clk ), .D ( new_AGEMA_signal_6642 ), .Q ( new_AGEMA_signal_6643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C ( clk ), .D ( new_AGEMA_signal_6648 ), .Q ( new_AGEMA_signal_6649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2166 ( .C ( clk ), .D ( new_AGEMA_signal_6654 ), .Q ( new_AGEMA_signal_6655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2170 ( .C ( clk ), .D ( new_AGEMA_signal_6658 ), .Q ( new_AGEMA_signal_6659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2174 ( .C ( clk ), .D ( new_AGEMA_signal_6662 ), .Q ( new_AGEMA_signal_6663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2178 ( .C ( clk ), .D ( new_AGEMA_signal_6666 ), .Q ( new_AGEMA_signal_6667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2182 ( .C ( clk ), .D ( new_AGEMA_signal_6670 ), .Q ( new_AGEMA_signal_6671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2186 ( .C ( clk ), .D ( new_AGEMA_signal_6674 ), .Q ( new_AGEMA_signal_6675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2190 ( .C ( clk ), .D ( new_AGEMA_signal_6678 ), .Q ( new_AGEMA_signal_6679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2218 ( .C ( clk ), .D ( new_AGEMA_signal_6706 ), .Q ( new_AGEMA_signal_6707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2222 ( .C ( clk ), .D ( new_AGEMA_signal_6710 ), .Q ( new_AGEMA_signal_6711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2226 ( .C ( clk ), .D ( new_AGEMA_signal_6714 ), .Q ( new_AGEMA_signal_6715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2232 ( .C ( clk ), .D ( new_AGEMA_signal_6720 ), .Q ( new_AGEMA_signal_6721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2238 ( .C ( clk ), .D ( new_AGEMA_signal_6726 ), .Q ( new_AGEMA_signal_6727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2244 ( .C ( clk ), .D ( new_AGEMA_signal_6732 ), .Q ( new_AGEMA_signal_6733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2248 ( .C ( clk ), .D ( new_AGEMA_signal_6736 ), .Q ( new_AGEMA_signal_6737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2252 ( .C ( clk ), .D ( new_AGEMA_signal_6740 ), .Q ( new_AGEMA_signal_6741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C ( clk ), .D ( new_AGEMA_signal_6744 ), .Q ( new_AGEMA_signal_6745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2278 ( .C ( clk ), .D ( new_AGEMA_signal_6766 ), .Q ( new_AGEMA_signal_6767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2282 ( .C ( clk ), .D ( new_AGEMA_signal_6770 ), .Q ( new_AGEMA_signal_6771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2286 ( .C ( clk ), .D ( new_AGEMA_signal_6774 ), .Q ( new_AGEMA_signal_6775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2302 ( .C ( clk ), .D ( new_AGEMA_signal_6790 ), .Q ( new_AGEMA_signal_6791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2306 ( .C ( clk ), .D ( new_AGEMA_signal_6794 ), .Q ( new_AGEMA_signal_6795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2310 ( .C ( clk ), .D ( new_AGEMA_signal_6798 ), .Q ( new_AGEMA_signal_6799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2314 ( .C ( clk ), .D ( new_AGEMA_signal_6802 ), .Q ( new_AGEMA_signal_6803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2318 ( .C ( clk ), .D ( new_AGEMA_signal_6806 ), .Q ( new_AGEMA_signal_6807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2322 ( .C ( clk ), .D ( new_AGEMA_signal_6810 ), .Q ( new_AGEMA_signal_6811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2326 ( .C ( clk ), .D ( new_AGEMA_signal_6814 ), .Q ( new_AGEMA_signal_6815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2330 ( .C ( clk ), .D ( new_AGEMA_signal_6818 ), .Q ( new_AGEMA_signal_6819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2334 ( .C ( clk ), .D ( new_AGEMA_signal_6822 ), .Q ( new_AGEMA_signal_6823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2338 ( .C ( clk ), .D ( new_AGEMA_signal_6826 ), .Q ( new_AGEMA_signal_6827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2342 ( .C ( clk ), .D ( new_AGEMA_signal_6830 ), .Q ( new_AGEMA_signal_6831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2346 ( .C ( clk ), .D ( new_AGEMA_signal_6834 ), .Q ( new_AGEMA_signal_6835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2350 ( .C ( clk ), .D ( new_AGEMA_signal_6838 ), .Q ( new_AGEMA_signal_6839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2354 ( .C ( clk ), .D ( new_AGEMA_signal_6842 ), .Q ( new_AGEMA_signal_6843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2358 ( .C ( clk ), .D ( new_AGEMA_signal_6846 ), .Q ( new_AGEMA_signal_6847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2386 ( .C ( clk ), .D ( new_AGEMA_signal_6874 ), .Q ( new_AGEMA_signal_6875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2390 ( .C ( clk ), .D ( new_AGEMA_signal_6878 ), .Q ( new_AGEMA_signal_6879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2394 ( .C ( clk ), .D ( new_AGEMA_signal_6882 ), .Q ( new_AGEMA_signal_6883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2398 ( .C ( clk ), .D ( new_AGEMA_signal_6886 ), .Q ( new_AGEMA_signal_6887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2402 ( .C ( clk ), .D ( new_AGEMA_signal_6890 ), .Q ( new_AGEMA_signal_6891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2406 ( .C ( clk ), .D ( new_AGEMA_signal_6894 ), .Q ( new_AGEMA_signal_6895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2464 ( .C ( clk ), .D ( new_AGEMA_signal_6952 ), .Q ( new_AGEMA_signal_6953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2468 ( .C ( clk ), .D ( new_AGEMA_signal_6956 ), .Q ( new_AGEMA_signal_6957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2472 ( .C ( clk ), .D ( new_AGEMA_signal_6960 ), .Q ( new_AGEMA_signal_6961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2506 ( .C ( clk ), .D ( new_AGEMA_signal_6994 ), .Q ( new_AGEMA_signal_6995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2510 ( .C ( clk ), .D ( new_AGEMA_signal_6998 ), .Q ( new_AGEMA_signal_6999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2514 ( .C ( clk ), .D ( new_AGEMA_signal_7002 ), .Q ( new_AGEMA_signal_7003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2518 ( .C ( clk ), .D ( new_AGEMA_signal_7006 ), .Q ( new_AGEMA_signal_7007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2522 ( .C ( clk ), .D ( new_AGEMA_signal_7010 ), .Q ( new_AGEMA_signal_7011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2526 ( .C ( clk ), .D ( new_AGEMA_signal_7014 ), .Q ( new_AGEMA_signal_7015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2530 ( .C ( clk ), .D ( new_AGEMA_signal_7018 ), .Q ( new_AGEMA_signal_7019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2534 ( .C ( clk ), .D ( new_AGEMA_signal_7022 ), .Q ( new_AGEMA_signal_7023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2538 ( .C ( clk ), .D ( new_AGEMA_signal_7026 ), .Q ( new_AGEMA_signal_7027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2542 ( .C ( clk ), .D ( new_AGEMA_signal_7030 ), .Q ( new_AGEMA_signal_7031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2546 ( .C ( clk ), .D ( new_AGEMA_signal_7034 ), .Q ( new_AGEMA_signal_7035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2550 ( .C ( clk ), .D ( new_AGEMA_signal_7038 ), .Q ( new_AGEMA_signal_7039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2580 ( .C ( clk ), .D ( new_AGEMA_signal_7068 ), .Q ( new_AGEMA_signal_7069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2588 ( .C ( clk ), .D ( new_AGEMA_signal_7076 ), .Q ( new_AGEMA_signal_7077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2596 ( .C ( clk ), .D ( new_AGEMA_signal_7084 ), .Q ( new_AGEMA_signal_7085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2610 ( .C ( clk ), .D ( new_AGEMA_signal_7098 ), .Q ( new_AGEMA_signal_7099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2618 ( .C ( clk ), .D ( new_AGEMA_signal_7106 ), .Q ( new_AGEMA_signal_7107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2626 ( .C ( clk ), .D ( new_AGEMA_signal_7114 ), .Q ( new_AGEMA_signal_7115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2632 ( .C ( clk ), .D ( new_AGEMA_signal_7120 ), .Q ( new_AGEMA_signal_7121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2638 ( .C ( clk ), .D ( new_AGEMA_signal_7126 ), .Q ( new_AGEMA_signal_7127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2644 ( .C ( clk ), .D ( new_AGEMA_signal_7132 ), .Q ( new_AGEMA_signal_7133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2662 ( .C ( clk ), .D ( new_AGEMA_signal_7150 ), .Q ( new_AGEMA_signal_7151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2668 ( .C ( clk ), .D ( new_AGEMA_signal_7156 ), .Q ( new_AGEMA_signal_7157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2674 ( .C ( clk ), .D ( new_AGEMA_signal_7162 ), .Q ( new_AGEMA_signal_7163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2686 ( .C ( clk ), .D ( new_AGEMA_signal_7174 ), .Q ( new_AGEMA_signal_7175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2692 ( .C ( clk ), .D ( new_AGEMA_signal_7180 ), .Q ( new_AGEMA_signal_7181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2698 ( .C ( clk ), .D ( new_AGEMA_signal_7186 ), .Q ( new_AGEMA_signal_7187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2704 ( .C ( clk ), .D ( new_AGEMA_signal_7192 ), .Q ( new_AGEMA_signal_7193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2710 ( .C ( clk ), .D ( new_AGEMA_signal_7198 ), .Q ( new_AGEMA_signal_7199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2716 ( .C ( clk ), .D ( new_AGEMA_signal_7204 ), .Q ( new_AGEMA_signal_7205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2740 ( .C ( clk ), .D ( new_AGEMA_signal_7228 ), .Q ( new_AGEMA_signal_7229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2746 ( .C ( clk ), .D ( new_AGEMA_signal_7234 ), .Q ( new_AGEMA_signal_7235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2752 ( .C ( clk ), .D ( new_AGEMA_signal_7240 ), .Q ( new_AGEMA_signal_7241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2758 ( .C ( clk ), .D ( new_AGEMA_signal_7246 ), .Q ( new_AGEMA_signal_7247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2764 ( .C ( clk ), .D ( new_AGEMA_signal_7252 ), .Q ( new_AGEMA_signal_7253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2770 ( .C ( clk ), .D ( new_AGEMA_signal_7258 ), .Q ( new_AGEMA_signal_7259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2782 ( .C ( clk ), .D ( new_AGEMA_signal_7270 ), .Q ( new_AGEMA_signal_7271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2788 ( .C ( clk ), .D ( new_AGEMA_signal_7276 ), .Q ( new_AGEMA_signal_7277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2794 ( .C ( clk ), .D ( new_AGEMA_signal_7282 ), .Q ( new_AGEMA_signal_7283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2838 ( .C ( clk ), .D ( new_AGEMA_signal_7326 ), .Q ( new_AGEMA_signal_7327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2846 ( .C ( clk ), .D ( new_AGEMA_signal_7334 ), .Q ( new_AGEMA_signal_7335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2854 ( .C ( clk ), .D ( new_AGEMA_signal_7342 ), .Q ( new_AGEMA_signal_7343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2860 ( .C ( clk ), .D ( new_AGEMA_signal_7348 ), .Q ( new_AGEMA_signal_7349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2866 ( .C ( clk ), .D ( new_AGEMA_signal_7354 ), .Q ( new_AGEMA_signal_7355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2872 ( .C ( clk ), .D ( new_AGEMA_signal_7360 ), .Q ( new_AGEMA_signal_7361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2944 ( .C ( clk ), .D ( new_AGEMA_signal_7432 ), .Q ( new_AGEMA_signal_7433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2950 ( .C ( clk ), .D ( new_AGEMA_signal_7438 ), .Q ( new_AGEMA_signal_7439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2956 ( .C ( clk ), .D ( new_AGEMA_signal_7444 ), .Q ( new_AGEMA_signal_7445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3040 ( .C ( clk ), .D ( new_AGEMA_signal_7528 ), .Q ( new_AGEMA_signal_7529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3046 ( .C ( clk ), .D ( new_AGEMA_signal_7534 ), .Q ( new_AGEMA_signal_7535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3052 ( .C ( clk ), .D ( new_AGEMA_signal_7540 ), .Q ( new_AGEMA_signal_7541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3058 ( .C ( clk ), .D ( new_AGEMA_signal_7546 ), .Q ( new_AGEMA_signal_7547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3064 ( .C ( clk ), .D ( new_AGEMA_signal_7552 ), .Q ( new_AGEMA_signal_7553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3070 ( .C ( clk ), .D ( new_AGEMA_signal_7558 ), .Q ( new_AGEMA_signal_7559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3096 ( .C ( clk ), .D ( new_AGEMA_signal_7584 ), .Q ( new_AGEMA_signal_7585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3104 ( .C ( clk ), .D ( new_AGEMA_signal_7592 ), .Q ( new_AGEMA_signal_7593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3112 ( .C ( clk ), .D ( new_AGEMA_signal_7600 ), .Q ( new_AGEMA_signal_7601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3186 ( .C ( clk ), .D ( new_AGEMA_signal_7674 ), .Q ( new_AGEMA_signal_7675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3194 ( .C ( clk ), .D ( new_AGEMA_signal_7682 ), .Q ( new_AGEMA_signal_7683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3202 ( .C ( clk ), .D ( new_AGEMA_signal_7690 ), .Q ( new_AGEMA_signal_7691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3232 ( .C ( clk ), .D ( new_AGEMA_signal_7720 ), .Q ( new_AGEMA_signal_7721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3238 ( .C ( clk ), .D ( new_AGEMA_signal_7726 ), .Q ( new_AGEMA_signal_7727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3244 ( .C ( clk ), .D ( new_AGEMA_signal_7732 ), .Q ( new_AGEMA_signal_7733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3256 ( .C ( clk ), .D ( new_AGEMA_signal_7744 ), .Q ( new_AGEMA_signal_7745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3264 ( .C ( clk ), .D ( new_AGEMA_signal_7752 ), .Q ( new_AGEMA_signal_7753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3272 ( .C ( clk ), .D ( new_AGEMA_signal_7760 ), .Q ( new_AGEMA_signal_7761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3298 ( .C ( clk ), .D ( new_AGEMA_signal_7786 ), .Q ( new_AGEMA_signal_7787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3306 ( .C ( clk ), .D ( new_AGEMA_signal_7794 ), .Q ( new_AGEMA_signal_7795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3314 ( .C ( clk ), .D ( new_AGEMA_signal_7802 ), .Q ( new_AGEMA_signal_7803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3358 ( .C ( clk ), .D ( new_AGEMA_signal_7846 ), .Q ( new_AGEMA_signal_7847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3366 ( .C ( clk ), .D ( new_AGEMA_signal_7854 ), .Q ( new_AGEMA_signal_7855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3374 ( .C ( clk ), .D ( new_AGEMA_signal_7862 ), .Q ( new_AGEMA_signal_7863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3496 ( .C ( clk ), .D ( new_AGEMA_signal_7984 ), .Q ( new_AGEMA_signal_7985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3504 ( .C ( clk ), .D ( new_AGEMA_signal_7992 ), .Q ( new_AGEMA_signal_7993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3512 ( .C ( clk ), .D ( new_AGEMA_signal_8000 ), .Q ( new_AGEMA_signal_8001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3550 ( .C ( clk ), .D ( new_AGEMA_signal_8038 ), .Q ( new_AGEMA_signal_8039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3558 ( .C ( clk ), .D ( new_AGEMA_signal_8046 ), .Q ( new_AGEMA_signal_8047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3566 ( .C ( clk ), .D ( new_AGEMA_signal_8054 ), .Q ( new_AGEMA_signal_8055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3646 ( .C ( clk ), .D ( new_AGEMA_signal_8134 ), .Q ( new_AGEMA_signal_8135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3654 ( .C ( clk ), .D ( new_AGEMA_signal_8142 ), .Q ( new_AGEMA_signal_8143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3662 ( .C ( clk ), .D ( new_AGEMA_signal_8150 ), .Q ( new_AGEMA_signal_8151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3670 ( .C ( clk ), .D ( new_AGEMA_signal_8158 ), .Q ( new_AGEMA_signal_8159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3678 ( .C ( clk ), .D ( new_AGEMA_signal_8166 ), .Q ( new_AGEMA_signal_8167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3686 ( .C ( clk ), .D ( new_AGEMA_signal_8174 ), .Q ( new_AGEMA_signal_8175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3928 ( .C ( clk ), .D ( new_AGEMA_signal_8416 ), .Q ( new_AGEMA_signal_8417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3938 ( .C ( clk ), .D ( new_AGEMA_signal_8426 ), .Q ( new_AGEMA_signal_8427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3948 ( .C ( clk ), .D ( new_AGEMA_signal_8436 ), .Q ( new_AGEMA_signal_8437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4078 ( .C ( clk ), .D ( new_AGEMA_signal_8566 ), .Q ( new_AGEMA_signal_8567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4088 ( .C ( clk ), .D ( new_AGEMA_signal_8576 ), .Q ( new_AGEMA_signal_8577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4098 ( .C ( clk ), .D ( new_AGEMA_signal_8586 ), .Q ( new_AGEMA_signal_8587 ) ) ;

    /* cells in depth 7 */
    buf_clk new_AGEMA_reg_buffer_1949 ( .C ( clk ), .D ( new_AGEMA_signal_6437 ), .Q ( new_AGEMA_signal_6438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C ( clk ), .D ( new_AGEMA_signal_6441 ), .Q ( new_AGEMA_signal_6442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C ( clk ), .D ( new_AGEMA_signal_6445 ), .Q ( new_AGEMA_signal_6446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C ( clk ), .D ( new_AGEMA_signal_6449 ), .Q ( new_AGEMA_signal_6450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C ( clk ), .D ( new_AGEMA_signal_6453 ), .Q ( new_AGEMA_signal_6454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C ( clk ), .D ( new_AGEMA_signal_6457 ), .Q ( new_AGEMA_signal_6458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C ( clk ), .D ( new_AGEMA_signal_6323 ), .Q ( new_AGEMA_signal_6460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C ( clk ), .D ( new_AGEMA_signal_6325 ), .Q ( new_AGEMA_signal_6462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C ( clk ), .D ( new_AGEMA_signal_6327 ), .Q ( new_AGEMA_signal_6464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C ( clk ), .D ( n1966 ), .Q ( new_AGEMA_signal_6466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C ( clk ), .D ( new_AGEMA_signal_1700 ), .Q ( new_AGEMA_signal_6468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C ( clk ), .D ( new_AGEMA_signal_1701 ), .Q ( new_AGEMA_signal_6470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C ( clk ), .D ( new_AGEMA_signal_6473 ), .Q ( new_AGEMA_signal_6474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C ( clk ), .D ( new_AGEMA_signal_6477 ), .Q ( new_AGEMA_signal_6478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C ( clk ), .D ( new_AGEMA_signal_6481 ), .Q ( new_AGEMA_signal_6482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C ( clk ), .D ( new_AGEMA_signal_6215 ), .Q ( new_AGEMA_signal_6484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C ( clk ), .D ( new_AGEMA_signal_6217 ), .Q ( new_AGEMA_signal_6486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C ( clk ), .D ( new_AGEMA_signal_6219 ), .Q ( new_AGEMA_signal_6488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C ( clk ), .D ( new_AGEMA_signal_6491 ), .Q ( new_AGEMA_signal_6492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C ( clk ), .D ( new_AGEMA_signal_6495 ), .Q ( new_AGEMA_signal_6496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C ( clk ), .D ( new_AGEMA_signal_6499 ), .Q ( new_AGEMA_signal_6500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2013 ( .C ( clk ), .D ( n1996 ), .Q ( new_AGEMA_signal_6502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C ( clk ), .D ( new_AGEMA_signal_1720 ), .Q ( new_AGEMA_signal_6504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C ( clk ), .D ( new_AGEMA_signal_1721 ), .Q ( new_AGEMA_signal_6506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C ( clk ), .D ( new_AGEMA_signal_6509 ), .Q ( new_AGEMA_signal_6510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C ( clk ), .D ( new_AGEMA_signal_6513 ), .Q ( new_AGEMA_signal_6514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C ( clk ), .D ( new_AGEMA_signal_6517 ), .Q ( new_AGEMA_signal_6518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C ( clk ), .D ( new_AGEMA_signal_6521 ), .Q ( new_AGEMA_signal_6522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C ( clk ), .D ( new_AGEMA_signal_6525 ), .Q ( new_AGEMA_signal_6526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2041 ( .C ( clk ), .D ( new_AGEMA_signal_6529 ), .Q ( new_AGEMA_signal_6530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C ( clk ), .D ( n2033 ), .Q ( new_AGEMA_signal_6532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C ( clk ), .D ( new_AGEMA_signal_1732 ), .Q ( new_AGEMA_signal_6534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C ( clk ), .D ( new_AGEMA_signal_1733 ), .Q ( new_AGEMA_signal_6536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C ( clk ), .D ( new_AGEMA_signal_6083 ), .Q ( new_AGEMA_signal_6538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C ( clk ), .D ( new_AGEMA_signal_6085 ), .Q ( new_AGEMA_signal_6540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C ( clk ), .D ( new_AGEMA_signal_6087 ), .Q ( new_AGEMA_signal_6542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C ( clk ), .D ( new_AGEMA_signal_6113 ), .Q ( new_AGEMA_signal_6544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C ( clk ), .D ( new_AGEMA_signal_6115 ), .Q ( new_AGEMA_signal_6546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C ( clk ), .D ( new_AGEMA_signal_6117 ), .Q ( new_AGEMA_signal_6548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C ( clk ), .D ( new_AGEMA_signal_6197 ), .Q ( new_AGEMA_signal_6550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C ( clk ), .D ( new_AGEMA_signal_6199 ), .Q ( new_AGEMA_signal_6552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C ( clk ), .D ( new_AGEMA_signal_6201 ), .Q ( new_AGEMA_signal_6554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C ( clk ), .D ( new_AGEMA_signal_6557 ), .Q ( new_AGEMA_signal_6558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C ( clk ), .D ( new_AGEMA_signal_6561 ), .Q ( new_AGEMA_signal_6562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C ( clk ), .D ( new_AGEMA_signal_6565 ), .Q ( new_AGEMA_signal_6566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C ( clk ), .D ( new_AGEMA_signal_6569 ), .Q ( new_AGEMA_signal_6570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C ( clk ), .D ( new_AGEMA_signal_6573 ), .Q ( new_AGEMA_signal_6574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C ( clk ), .D ( new_AGEMA_signal_6577 ), .Q ( new_AGEMA_signal_6578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C ( clk ), .D ( new_AGEMA_signal_6581 ), .Q ( new_AGEMA_signal_6582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C ( clk ), .D ( new_AGEMA_signal_6585 ), .Q ( new_AGEMA_signal_6586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C ( clk ), .D ( new_AGEMA_signal_6589 ), .Q ( new_AGEMA_signal_6590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C ( clk ), .D ( n2089 ), .Q ( new_AGEMA_signal_6592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C ( clk ), .D ( new_AGEMA_signal_1762 ), .Q ( new_AGEMA_signal_6594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C ( clk ), .D ( new_AGEMA_signal_1763 ), .Q ( new_AGEMA_signal_6596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C ( clk ), .D ( n2092 ), .Q ( new_AGEMA_signal_6598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C ( clk ), .D ( new_AGEMA_signal_1766 ), .Q ( new_AGEMA_signal_6600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C ( clk ), .D ( new_AGEMA_signal_1767 ), .Q ( new_AGEMA_signal_6602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C ( clk ), .D ( n2115 ), .Q ( new_AGEMA_signal_6604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C ( clk ), .D ( new_AGEMA_signal_1438 ), .Q ( new_AGEMA_signal_6606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C ( clk ), .D ( new_AGEMA_signal_1439 ), .Q ( new_AGEMA_signal_6608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C ( clk ), .D ( new_AGEMA_signal_6611 ), .Q ( new_AGEMA_signal_6612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C ( clk ), .D ( new_AGEMA_signal_6615 ), .Q ( new_AGEMA_signal_6616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C ( clk ), .D ( new_AGEMA_signal_6619 ), .Q ( new_AGEMA_signal_6620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C ( clk ), .D ( n2687 ), .Q ( new_AGEMA_signal_6622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C ( clk ), .D ( new_AGEMA_signal_1698 ), .Q ( new_AGEMA_signal_6624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C ( clk ), .D ( new_AGEMA_signal_1699 ), .Q ( new_AGEMA_signal_6626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C ( clk ), .D ( new_AGEMA_signal_6629 ), .Q ( new_AGEMA_signal_6630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2145 ( .C ( clk ), .D ( new_AGEMA_signal_6633 ), .Q ( new_AGEMA_signal_6634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2149 ( .C ( clk ), .D ( new_AGEMA_signal_6637 ), .Q ( new_AGEMA_signal_6638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2155 ( .C ( clk ), .D ( new_AGEMA_signal_6643 ), .Q ( new_AGEMA_signal_6644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2161 ( .C ( clk ), .D ( new_AGEMA_signal_6649 ), .Q ( new_AGEMA_signal_6650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2167 ( .C ( clk ), .D ( new_AGEMA_signal_6655 ), .Q ( new_AGEMA_signal_6656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2171 ( .C ( clk ), .D ( new_AGEMA_signal_6659 ), .Q ( new_AGEMA_signal_6660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2175 ( .C ( clk ), .D ( new_AGEMA_signal_6663 ), .Q ( new_AGEMA_signal_6664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2179 ( .C ( clk ), .D ( new_AGEMA_signal_6667 ), .Q ( new_AGEMA_signal_6668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2183 ( .C ( clk ), .D ( new_AGEMA_signal_6671 ), .Q ( new_AGEMA_signal_6672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2187 ( .C ( clk ), .D ( new_AGEMA_signal_6675 ), .Q ( new_AGEMA_signal_6676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2191 ( .C ( clk ), .D ( new_AGEMA_signal_6679 ), .Q ( new_AGEMA_signal_6680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2193 ( .C ( clk ), .D ( n2193 ), .Q ( new_AGEMA_signal_6682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2195 ( .C ( clk ), .D ( new_AGEMA_signal_1802 ), .Q ( new_AGEMA_signal_6684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2197 ( .C ( clk ), .D ( new_AGEMA_signal_1803 ), .Q ( new_AGEMA_signal_6686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2199 ( .C ( clk ), .D ( n2202 ), .Q ( new_AGEMA_signal_6688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2201 ( .C ( clk ), .D ( new_AGEMA_signal_2090 ), .Q ( new_AGEMA_signal_6690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2203 ( .C ( clk ), .D ( new_AGEMA_signal_2091 ), .Q ( new_AGEMA_signal_6692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C ( clk ), .D ( n2228 ), .Q ( new_AGEMA_signal_6694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C ( clk ), .D ( new_AGEMA_signal_1486 ), .Q ( new_AGEMA_signal_6696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2209 ( .C ( clk ), .D ( new_AGEMA_signal_1487 ), .Q ( new_AGEMA_signal_6698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2211 ( .C ( clk ), .D ( n2235 ), .Q ( new_AGEMA_signal_6700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2213 ( .C ( clk ), .D ( new_AGEMA_signal_1688 ), .Q ( new_AGEMA_signal_6702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2215 ( .C ( clk ), .D ( new_AGEMA_signal_1689 ), .Q ( new_AGEMA_signal_6704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2219 ( .C ( clk ), .D ( new_AGEMA_signal_6707 ), .Q ( new_AGEMA_signal_6708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2223 ( .C ( clk ), .D ( new_AGEMA_signal_6711 ), .Q ( new_AGEMA_signal_6712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2227 ( .C ( clk ), .D ( new_AGEMA_signal_6715 ), .Q ( new_AGEMA_signal_6716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2233 ( .C ( clk ), .D ( new_AGEMA_signal_6721 ), .Q ( new_AGEMA_signal_6722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2239 ( .C ( clk ), .D ( new_AGEMA_signal_6727 ), .Q ( new_AGEMA_signal_6728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2245 ( .C ( clk ), .D ( new_AGEMA_signal_6733 ), .Q ( new_AGEMA_signal_6734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2249 ( .C ( clk ), .D ( new_AGEMA_signal_6737 ), .Q ( new_AGEMA_signal_6738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C ( clk ), .D ( new_AGEMA_signal_6741 ), .Q ( new_AGEMA_signal_6742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2257 ( .C ( clk ), .D ( new_AGEMA_signal_6745 ), .Q ( new_AGEMA_signal_6746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2259 ( .C ( clk ), .D ( n2752 ), .Q ( new_AGEMA_signal_6748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2261 ( .C ( clk ), .D ( new_AGEMA_signal_2108 ), .Q ( new_AGEMA_signal_6750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2263 ( .C ( clk ), .D ( new_AGEMA_signal_2109 ), .Q ( new_AGEMA_signal_6752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2265 ( .C ( clk ), .D ( new_AGEMA_signal_6279 ), .Q ( new_AGEMA_signal_6754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2267 ( .C ( clk ), .D ( new_AGEMA_signal_6285 ), .Q ( new_AGEMA_signal_6756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2269 ( .C ( clk ), .D ( new_AGEMA_signal_6291 ), .Q ( new_AGEMA_signal_6758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2271 ( .C ( clk ), .D ( n2293 ), .Q ( new_AGEMA_signal_6760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2273 ( .C ( clk ), .D ( new_AGEMA_signal_1844 ), .Q ( new_AGEMA_signal_6762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2275 ( .C ( clk ), .D ( new_AGEMA_signal_1845 ), .Q ( new_AGEMA_signal_6764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2279 ( .C ( clk ), .D ( new_AGEMA_signal_6767 ), .Q ( new_AGEMA_signal_6768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2283 ( .C ( clk ), .D ( new_AGEMA_signal_6771 ), .Q ( new_AGEMA_signal_6772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2287 ( .C ( clk ), .D ( new_AGEMA_signal_6775 ), .Q ( new_AGEMA_signal_6776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2289 ( .C ( clk ), .D ( n2357 ), .Q ( new_AGEMA_signal_6778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2291 ( .C ( clk ), .D ( new_AGEMA_signal_1862 ), .Q ( new_AGEMA_signal_6780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2293 ( .C ( clk ), .D ( new_AGEMA_signal_1863 ), .Q ( new_AGEMA_signal_6782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2295 ( .C ( clk ), .D ( n2386 ), .Q ( new_AGEMA_signal_6784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2297 ( .C ( clk ), .D ( new_AGEMA_signal_1872 ), .Q ( new_AGEMA_signal_6786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2299 ( .C ( clk ), .D ( new_AGEMA_signal_1873 ), .Q ( new_AGEMA_signal_6788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2303 ( .C ( clk ), .D ( new_AGEMA_signal_6791 ), .Q ( new_AGEMA_signal_6792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2307 ( .C ( clk ), .D ( new_AGEMA_signal_6795 ), .Q ( new_AGEMA_signal_6796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2311 ( .C ( clk ), .D ( new_AGEMA_signal_6799 ), .Q ( new_AGEMA_signal_6800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2315 ( .C ( clk ), .D ( new_AGEMA_signal_6803 ), .Q ( new_AGEMA_signal_6804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2319 ( .C ( clk ), .D ( new_AGEMA_signal_6807 ), .Q ( new_AGEMA_signal_6808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2323 ( .C ( clk ), .D ( new_AGEMA_signal_6811 ), .Q ( new_AGEMA_signal_6812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2327 ( .C ( clk ), .D ( new_AGEMA_signal_6815 ), .Q ( new_AGEMA_signal_6816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2331 ( .C ( clk ), .D ( new_AGEMA_signal_6819 ), .Q ( new_AGEMA_signal_6820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2335 ( .C ( clk ), .D ( new_AGEMA_signal_6823 ), .Q ( new_AGEMA_signal_6824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2339 ( .C ( clk ), .D ( new_AGEMA_signal_6827 ), .Q ( new_AGEMA_signal_6828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2343 ( .C ( clk ), .D ( new_AGEMA_signal_6831 ), .Q ( new_AGEMA_signal_6832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2347 ( .C ( clk ), .D ( new_AGEMA_signal_6835 ), .Q ( new_AGEMA_signal_6836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2351 ( .C ( clk ), .D ( new_AGEMA_signal_6839 ), .Q ( new_AGEMA_signal_6840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2355 ( .C ( clk ), .D ( new_AGEMA_signal_6843 ), .Q ( new_AGEMA_signal_6844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2359 ( .C ( clk ), .D ( new_AGEMA_signal_6847 ), .Q ( new_AGEMA_signal_6848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2361 ( .C ( clk ), .D ( n2433 ), .Q ( new_AGEMA_signal_6850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2363 ( .C ( clk ), .D ( new_AGEMA_signal_1886 ), .Q ( new_AGEMA_signal_6852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2365 ( .C ( clk ), .D ( new_AGEMA_signal_1887 ), .Q ( new_AGEMA_signal_6854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2367 ( .C ( clk ), .D ( new_AGEMA_signal_6103 ), .Q ( new_AGEMA_signal_6856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2369 ( .C ( clk ), .D ( new_AGEMA_signal_6107 ), .Q ( new_AGEMA_signal_6858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2371 ( .C ( clk ), .D ( new_AGEMA_signal_6111 ), .Q ( new_AGEMA_signal_6860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2373 ( .C ( clk ), .D ( n2459 ), .Q ( new_AGEMA_signal_6862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2375 ( .C ( clk ), .D ( new_AGEMA_signal_1838 ), .Q ( new_AGEMA_signal_6864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2377 ( .C ( clk ), .D ( new_AGEMA_signal_1839 ), .Q ( new_AGEMA_signal_6866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2379 ( .C ( clk ), .D ( n2467 ), .Q ( new_AGEMA_signal_6868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2381 ( .C ( clk ), .D ( new_AGEMA_signal_1550 ), .Q ( new_AGEMA_signal_6870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2383 ( .C ( clk ), .D ( new_AGEMA_signal_1551 ), .Q ( new_AGEMA_signal_6872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2387 ( .C ( clk ), .D ( new_AGEMA_signal_6875 ), .Q ( new_AGEMA_signal_6876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2391 ( .C ( clk ), .D ( new_AGEMA_signal_6879 ), .Q ( new_AGEMA_signal_6880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2395 ( .C ( clk ), .D ( new_AGEMA_signal_6883 ), .Q ( new_AGEMA_signal_6884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2399 ( .C ( clk ), .D ( new_AGEMA_signal_6887 ), .Q ( new_AGEMA_signal_6888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2403 ( .C ( clk ), .D ( new_AGEMA_signal_6891 ), .Q ( new_AGEMA_signal_6892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2407 ( .C ( clk ), .D ( new_AGEMA_signal_6895 ), .Q ( new_AGEMA_signal_6896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2409 ( .C ( clk ), .D ( n2489 ), .Q ( new_AGEMA_signal_6898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2411 ( .C ( clk ), .D ( new_AGEMA_signal_1590 ), .Q ( new_AGEMA_signal_6900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2413 ( .C ( clk ), .D ( new_AGEMA_signal_1591 ), .Q ( new_AGEMA_signal_6902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2415 ( .C ( clk ), .D ( n2497 ), .Q ( new_AGEMA_signal_6904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2417 ( .C ( clk ), .D ( new_AGEMA_signal_1592 ), .Q ( new_AGEMA_signal_6906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2419 ( .C ( clk ), .D ( new_AGEMA_signal_1593 ), .Q ( new_AGEMA_signal_6908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2421 ( .C ( clk ), .D ( n2506 ), .Q ( new_AGEMA_signal_6910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2423 ( .C ( clk ), .D ( new_AGEMA_signal_1912 ), .Q ( new_AGEMA_signal_6912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2425 ( .C ( clk ), .D ( new_AGEMA_signal_1913 ), .Q ( new_AGEMA_signal_6914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2427 ( .C ( clk ), .D ( n2542 ), .Q ( new_AGEMA_signal_6916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2429 ( .C ( clk ), .D ( new_AGEMA_signal_1924 ), .Q ( new_AGEMA_signal_6918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2431 ( .C ( clk ), .D ( new_AGEMA_signal_1925 ), .Q ( new_AGEMA_signal_6920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2433 ( .C ( clk ), .D ( n2558 ), .Q ( new_AGEMA_signal_6922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2435 ( .C ( clk ), .D ( new_AGEMA_signal_1930 ), .Q ( new_AGEMA_signal_6924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2437 ( .C ( clk ), .D ( new_AGEMA_signal_1931 ), .Q ( new_AGEMA_signal_6926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2439 ( .C ( clk ), .D ( n2566 ), .Q ( new_AGEMA_signal_6928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2441 ( .C ( clk ), .D ( new_AGEMA_signal_1934 ), .Q ( new_AGEMA_signal_6930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2443 ( .C ( clk ), .D ( new_AGEMA_signal_1935 ), .Q ( new_AGEMA_signal_6932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2445 ( .C ( clk ), .D ( n2581 ), .Q ( new_AGEMA_signal_6934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2447 ( .C ( clk ), .D ( new_AGEMA_signal_1610 ), .Q ( new_AGEMA_signal_6936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2449 ( .C ( clk ), .D ( new_AGEMA_signal_1611 ), .Q ( new_AGEMA_signal_6938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2451 ( .C ( clk ), .D ( n2603 ), .Q ( new_AGEMA_signal_6940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2453 ( .C ( clk ), .D ( new_AGEMA_signal_1950 ), .Q ( new_AGEMA_signal_6942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2455 ( .C ( clk ), .D ( new_AGEMA_signal_1951 ), .Q ( new_AGEMA_signal_6944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2457 ( .C ( clk ), .D ( n2620 ), .Q ( new_AGEMA_signal_6946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2459 ( .C ( clk ), .D ( new_AGEMA_signal_1952 ), .Q ( new_AGEMA_signal_6948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2461 ( .C ( clk ), .D ( new_AGEMA_signal_1953 ), .Q ( new_AGEMA_signal_6950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2465 ( .C ( clk ), .D ( new_AGEMA_signal_6953 ), .Q ( new_AGEMA_signal_6954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2469 ( .C ( clk ), .D ( new_AGEMA_signal_6957 ), .Q ( new_AGEMA_signal_6958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2473 ( .C ( clk ), .D ( new_AGEMA_signal_6961 ), .Q ( new_AGEMA_signal_6962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2475 ( .C ( clk ), .D ( n2653 ), .Q ( new_AGEMA_signal_6964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2477 ( .C ( clk ), .D ( new_AGEMA_signal_1636 ), .Q ( new_AGEMA_signal_6966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2479 ( .C ( clk ), .D ( new_AGEMA_signal_1637 ), .Q ( new_AGEMA_signal_6968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2481 ( .C ( clk ), .D ( n2665 ), .Q ( new_AGEMA_signal_6970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2483 ( .C ( clk ), .D ( new_AGEMA_signal_1684 ), .Q ( new_AGEMA_signal_6972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2485 ( .C ( clk ), .D ( new_AGEMA_signal_1685 ), .Q ( new_AGEMA_signal_6974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2487 ( .C ( clk ), .D ( n2691 ), .Q ( new_AGEMA_signal_6976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2489 ( .C ( clk ), .D ( new_AGEMA_signal_1642 ), .Q ( new_AGEMA_signal_6978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2491 ( .C ( clk ), .D ( new_AGEMA_signal_1643 ), .Q ( new_AGEMA_signal_6980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2493 ( .C ( clk ), .D ( n2717 ), .Q ( new_AGEMA_signal_6982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2495 ( .C ( clk ), .D ( new_AGEMA_signal_1970 ), .Q ( new_AGEMA_signal_6984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2497 ( .C ( clk ), .D ( new_AGEMA_signal_1971 ), .Q ( new_AGEMA_signal_6986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2499 ( .C ( clk ), .D ( n2729 ), .Q ( new_AGEMA_signal_6988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2501 ( .C ( clk ), .D ( new_AGEMA_signal_2210 ), .Q ( new_AGEMA_signal_6990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2503 ( .C ( clk ), .D ( new_AGEMA_signal_2211 ), .Q ( new_AGEMA_signal_6992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2507 ( .C ( clk ), .D ( new_AGEMA_signal_6995 ), .Q ( new_AGEMA_signal_6996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2511 ( .C ( clk ), .D ( new_AGEMA_signal_6999 ), .Q ( new_AGEMA_signal_7000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2515 ( .C ( clk ), .D ( new_AGEMA_signal_7003 ), .Q ( new_AGEMA_signal_7004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2519 ( .C ( clk ), .D ( new_AGEMA_signal_7007 ), .Q ( new_AGEMA_signal_7008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2523 ( .C ( clk ), .D ( new_AGEMA_signal_7011 ), .Q ( new_AGEMA_signal_7012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2527 ( .C ( clk ), .D ( new_AGEMA_signal_7015 ), .Q ( new_AGEMA_signal_7016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2531 ( .C ( clk ), .D ( new_AGEMA_signal_7019 ), .Q ( new_AGEMA_signal_7020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2535 ( .C ( clk ), .D ( new_AGEMA_signal_7023 ), .Q ( new_AGEMA_signal_7024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2539 ( .C ( clk ), .D ( new_AGEMA_signal_7027 ), .Q ( new_AGEMA_signal_7028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2543 ( .C ( clk ), .D ( new_AGEMA_signal_7031 ), .Q ( new_AGEMA_signal_7032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2547 ( .C ( clk ), .D ( new_AGEMA_signal_7035 ), .Q ( new_AGEMA_signal_7036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2551 ( .C ( clk ), .D ( new_AGEMA_signal_7039 ), .Q ( new_AGEMA_signal_7040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2553 ( .C ( clk ), .D ( new_AGEMA_signal_6239 ), .Q ( new_AGEMA_signal_7042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2557 ( .C ( clk ), .D ( new_AGEMA_signal_6241 ), .Q ( new_AGEMA_signal_7046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2561 ( .C ( clk ), .D ( new_AGEMA_signal_6243 ), .Q ( new_AGEMA_signal_7050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2565 ( .C ( clk ), .D ( n1956 ), .Q ( new_AGEMA_signal_7054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2569 ( .C ( clk ), .D ( new_AGEMA_signal_1692 ), .Q ( new_AGEMA_signal_7058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2573 ( .C ( clk ), .D ( new_AGEMA_signal_1693 ), .Q ( new_AGEMA_signal_7062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2581 ( .C ( clk ), .D ( new_AGEMA_signal_7069 ), .Q ( new_AGEMA_signal_7070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2589 ( .C ( clk ), .D ( new_AGEMA_signal_7077 ), .Q ( new_AGEMA_signal_7078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2597 ( .C ( clk ), .D ( new_AGEMA_signal_7085 ), .Q ( new_AGEMA_signal_7086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2611 ( .C ( clk ), .D ( new_AGEMA_signal_7099 ), .Q ( new_AGEMA_signal_7100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2619 ( .C ( clk ), .D ( new_AGEMA_signal_7107 ), .Q ( new_AGEMA_signal_7108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2627 ( .C ( clk ), .D ( new_AGEMA_signal_7115 ), .Q ( new_AGEMA_signal_7116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2633 ( .C ( clk ), .D ( new_AGEMA_signal_7121 ), .Q ( new_AGEMA_signal_7122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2639 ( .C ( clk ), .D ( new_AGEMA_signal_7127 ), .Q ( new_AGEMA_signal_7128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2645 ( .C ( clk ), .D ( new_AGEMA_signal_7133 ), .Q ( new_AGEMA_signal_7134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2649 ( .C ( clk ), .D ( n2023 ), .Q ( new_AGEMA_signal_7138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2653 ( .C ( clk ), .D ( new_AGEMA_signal_1390 ), .Q ( new_AGEMA_signal_7142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2657 ( .C ( clk ), .D ( new_AGEMA_signal_1391 ), .Q ( new_AGEMA_signal_7146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2663 ( .C ( clk ), .D ( new_AGEMA_signal_7151 ), .Q ( new_AGEMA_signal_7152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2669 ( .C ( clk ), .D ( new_AGEMA_signal_7157 ), .Q ( new_AGEMA_signal_7158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2675 ( .C ( clk ), .D ( new_AGEMA_signal_7163 ), .Q ( new_AGEMA_signal_7164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2687 ( .C ( clk ), .D ( new_AGEMA_signal_7175 ), .Q ( new_AGEMA_signal_7176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2693 ( .C ( clk ), .D ( new_AGEMA_signal_7181 ), .Q ( new_AGEMA_signal_7182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2699 ( .C ( clk ), .D ( new_AGEMA_signal_7187 ), .Q ( new_AGEMA_signal_7188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2705 ( .C ( clk ), .D ( new_AGEMA_signal_7193 ), .Q ( new_AGEMA_signal_7194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2711 ( .C ( clk ), .D ( new_AGEMA_signal_7199 ), .Q ( new_AGEMA_signal_7200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2717 ( .C ( clk ), .D ( new_AGEMA_signal_7205 ), .Q ( new_AGEMA_signal_7206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2727 ( .C ( clk ), .D ( n2094 ), .Q ( new_AGEMA_signal_7216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2731 ( .C ( clk ), .D ( new_AGEMA_signal_1768 ), .Q ( new_AGEMA_signal_7220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2735 ( .C ( clk ), .D ( new_AGEMA_signal_1769 ), .Q ( new_AGEMA_signal_7224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2741 ( .C ( clk ), .D ( new_AGEMA_signal_7229 ), .Q ( new_AGEMA_signal_7230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2747 ( .C ( clk ), .D ( new_AGEMA_signal_7235 ), .Q ( new_AGEMA_signal_7236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2753 ( .C ( clk ), .D ( new_AGEMA_signal_7241 ), .Q ( new_AGEMA_signal_7242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2759 ( .C ( clk ), .D ( new_AGEMA_signal_7247 ), .Q ( new_AGEMA_signal_7248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2765 ( .C ( clk ), .D ( new_AGEMA_signal_7253 ), .Q ( new_AGEMA_signal_7254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2771 ( .C ( clk ), .D ( new_AGEMA_signal_7259 ), .Q ( new_AGEMA_signal_7260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2783 ( .C ( clk ), .D ( new_AGEMA_signal_7271 ), .Q ( new_AGEMA_signal_7272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2789 ( .C ( clk ), .D ( new_AGEMA_signal_7277 ), .Q ( new_AGEMA_signal_7278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2795 ( .C ( clk ), .D ( new_AGEMA_signal_7283 ), .Q ( new_AGEMA_signal_7284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2805 ( .C ( clk ), .D ( n2181 ), .Q ( new_AGEMA_signal_7294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2809 ( .C ( clk ), .D ( new_AGEMA_signal_1796 ), .Q ( new_AGEMA_signal_7298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2813 ( .C ( clk ), .D ( new_AGEMA_signal_1797 ), .Q ( new_AGEMA_signal_7302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2817 ( .C ( clk ), .D ( n2195 ), .Q ( new_AGEMA_signal_7306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2821 ( .C ( clk ), .D ( new_AGEMA_signal_1800 ), .Q ( new_AGEMA_signal_7310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2825 ( .C ( clk ), .D ( new_AGEMA_signal_1801 ), .Q ( new_AGEMA_signal_7314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2839 ( .C ( clk ), .D ( new_AGEMA_signal_7327 ), .Q ( new_AGEMA_signal_7328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2847 ( .C ( clk ), .D ( new_AGEMA_signal_7335 ), .Q ( new_AGEMA_signal_7336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2855 ( .C ( clk ), .D ( new_AGEMA_signal_7343 ), .Q ( new_AGEMA_signal_7344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2861 ( .C ( clk ), .D ( new_AGEMA_signal_7349 ), .Q ( new_AGEMA_signal_7350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2867 ( .C ( clk ), .D ( new_AGEMA_signal_7355 ), .Q ( new_AGEMA_signal_7356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2873 ( .C ( clk ), .D ( new_AGEMA_signal_7361 ), .Q ( new_AGEMA_signal_7362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2877 ( .C ( clk ), .D ( n2237 ), .Q ( new_AGEMA_signal_7366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2881 ( .C ( clk ), .D ( new_AGEMA_signal_1488 ), .Q ( new_AGEMA_signal_7370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2885 ( .C ( clk ), .D ( new_AGEMA_signal_1489 ), .Q ( new_AGEMA_signal_7374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2889 ( .C ( clk ), .D ( n2248 ), .Q ( new_AGEMA_signal_7378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2893 ( .C ( clk ), .D ( new_AGEMA_signal_1818 ), .Q ( new_AGEMA_signal_7382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2897 ( .C ( clk ), .D ( new_AGEMA_signal_1819 ), .Q ( new_AGEMA_signal_7386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2913 ( .C ( clk ), .D ( n2294 ), .Q ( new_AGEMA_signal_7402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2917 ( .C ( clk ), .D ( new_AGEMA_signal_1518 ), .Q ( new_AGEMA_signal_7406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2921 ( .C ( clk ), .D ( new_AGEMA_signal_1519 ), .Q ( new_AGEMA_signal_7410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2925 ( .C ( clk ), .D ( n2323 ), .Q ( new_AGEMA_signal_7414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2929 ( .C ( clk ), .D ( new_AGEMA_signal_1848 ), .Q ( new_AGEMA_signal_7418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2933 ( .C ( clk ), .D ( new_AGEMA_signal_1849 ), .Q ( new_AGEMA_signal_7422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2945 ( .C ( clk ), .D ( new_AGEMA_signal_7433 ), .Q ( new_AGEMA_signal_7434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2951 ( .C ( clk ), .D ( new_AGEMA_signal_7439 ), .Q ( new_AGEMA_signal_7440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2957 ( .C ( clk ), .D ( new_AGEMA_signal_7445 ), .Q ( new_AGEMA_signal_7446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2961 ( .C ( clk ), .D ( n2360 ), .Q ( new_AGEMA_signal_7450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2965 ( .C ( clk ), .D ( new_AGEMA_signal_1864 ), .Q ( new_AGEMA_signal_7454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2969 ( .C ( clk ), .D ( new_AGEMA_signal_1865 ), .Q ( new_AGEMA_signal_7458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2979 ( .C ( clk ), .D ( n2394 ), .Q ( new_AGEMA_signal_7468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2983 ( .C ( clk ), .D ( new_AGEMA_signal_1556 ), .Q ( new_AGEMA_signal_7472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2987 ( .C ( clk ), .D ( new_AGEMA_signal_1557 ), .Q ( new_AGEMA_signal_7476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2991 ( .C ( clk ), .D ( n2406 ), .Q ( new_AGEMA_signal_7480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2995 ( .C ( clk ), .D ( new_AGEMA_signal_1876 ), .Q ( new_AGEMA_signal_7484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2999 ( .C ( clk ), .D ( new_AGEMA_signal_1877 ), .Q ( new_AGEMA_signal_7488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3003 ( .C ( clk ), .D ( new_AGEMA_signal_5939 ), .Q ( new_AGEMA_signal_7492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3007 ( .C ( clk ), .D ( new_AGEMA_signal_5941 ), .Q ( new_AGEMA_signal_7496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3011 ( .C ( clk ), .D ( new_AGEMA_signal_5943 ), .Q ( new_AGEMA_signal_7500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3021 ( .C ( clk ), .D ( new_AGEMA_signal_5945 ), .Q ( new_AGEMA_signal_7510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3025 ( .C ( clk ), .D ( new_AGEMA_signal_5947 ), .Q ( new_AGEMA_signal_7514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3029 ( .C ( clk ), .D ( new_AGEMA_signal_5949 ), .Q ( new_AGEMA_signal_7518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3041 ( .C ( clk ), .D ( new_AGEMA_signal_7529 ), .Q ( new_AGEMA_signal_7530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3047 ( .C ( clk ), .D ( new_AGEMA_signal_7535 ), .Q ( new_AGEMA_signal_7536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3053 ( .C ( clk ), .D ( new_AGEMA_signal_7541 ), .Q ( new_AGEMA_signal_7542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3059 ( .C ( clk ), .D ( new_AGEMA_signal_7547 ), .Q ( new_AGEMA_signal_7548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3065 ( .C ( clk ), .D ( new_AGEMA_signal_7553 ), .Q ( new_AGEMA_signal_7554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3071 ( .C ( clk ), .D ( new_AGEMA_signal_7559 ), .Q ( new_AGEMA_signal_7560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3075 ( .C ( clk ), .D ( n2499 ), .Q ( new_AGEMA_signal_7564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3079 ( .C ( clk ), .D ( new_AGEMA_signal_1596 ), .Q ( new_AGEMA_signal_7568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3083 ( .C ( clk ), .D ( new_AGEMA_signal_1597 ), .Q ( new_AGEMA_signal_7572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3097 ( .C ( clk ), .D ( new_AGEMA_signal_7585 ), .Q ( new_AGEMA_signal_7586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3105 ( .C ( clk ), .D ( new_AGEMA_signal_7593 ), .Q ( new_AGEMA_signal_7594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3113 ( .C ( clk ), .D ( new_AGEMA_signal_7601 ), .Q ( new_AGEMA_signal_7602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3123 ( .C ( clk ), .D ( n2582 ), .Q ( new_AGEMA_signal_7612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3127 ( .C ( clk ), .D ( new_AGEMA_signal_1944 ), .Q ( new_AGEMA_signal_7616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3131 ( .C ( clk ), .D ( new_AGEMA_signal_1945 ), .Q ( new_AGEMA_signal_7620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3135 ( .C ( clk ), .D ( n2605 ), .Q ( new_AGEMA_signal_7624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3139 ( .C ( clk ), .D ( new_AGEMA_signal_1948 ), .Q ( new_AGEMA_signal_7628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3143 ( .C ( clk ), .D ( new_AGEMA_signal_1949 ), .Q ( new_AGEMA_signal_7632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3147 ( .C ( clk ), .D ( n2632 ), .Q ( new_AGEMA_signal_7636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3151 ( .C ( clk ), .D ( new_AGEMA_signal_1630 ), .Q ( new_AGEMA_signal_7640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3155 ( .C ( clk ), .D ( new_AGEMA_signal_1631 ), .Q ( new_AGEMA_signal_7644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3159 ( .C ( clk ), .D ( n2655 ), .Q ( new_AGEMA_signal_7648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3163 ( .C ( clk ), .D ( new_AGEMA_signal_1962 ), .Q ( new_AGEMA_signal_7652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3167 ( .C ( clk ), .D ( new_AGEMA_signal_1963 ), .Q ( new_AGEMA_signal_7656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3171 ( .C ( clk ), .D ( n2695 ), .Q ( new_AGEMA_signal_7660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3175 ( .C ( clk ), .D ( new_AGEMA_signal_1968 ), .Q ( new_AGEMA_signal_7664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3179 ( .C ( clk ), .D ( new_AGEMA_signal_1969 ), .Q ( new_AGEMA_signal_7668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3187 ( .C ( clk ), .D ( new_AGEMA_signal_7675 ), .Q ( new_AGEMA_signal_7676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3195 ( .C ( clk ), .D ( new_AGEMA_signal_7683 ), .Q ( new_AGEMA_signal_7684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3203 ( .C ( clk ), .D ( new_AGEMA_signal_7691 ), .Q ( new_AGEMA_signal_7692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3213 ( .C ( clk ), .D ( n2770 ), .Q ( new_AGEMA_signal_7702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3217 ( .C ( clk ), .D ( new_AGEMA_signal_1984 ), .Q ( new_AGEMA_signal_7706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3221 ( .C ( clk ), .D ( new_AGEMA_signal_1985 ), .Q ( new_AGEMA_signal_7710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3233 ( .C ( clk ), .D ( new_AGEMA_signal_7721 ), .Q ( new_AGEMA_signal_7722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3239 ( .C ( clk ), .D ( new_AGEMA_signal_7727 ), .Q ( new_AGEMA_signal_7728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3245 ( .C ( clk ), .D ( new_AGEMA_signal_7733 ), .Q ( new_AGEMA_signal_7734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3257 ( .C ( clk ), .D ( new_AGEMA_signal_7745 ), .Q ( new_AGEMA_signal_7746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3265 ( .C ( clk ), .D ( new_AGEMA_signal_7753 ), .Q ( new_AGEMA_signal_7754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3273 ( .C ( clk ), .D ( new_AGEMA_signal_7761 ), .Q ( new_AGEMA_signal_7762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3299 ( .C ( clk ), .D ( new_AGEMA_signal_7787 ), .Q ( new_AGEMA_signal_7788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3307 ( .C ( clk ), .D ( new_AGEMA_signal_7795 ), .Q ( new_AGEMA_signal_7796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3315 ( .C ( clk ), .D ( new_AGEMA_signal_7803 ), .Q ( new_AGEMA_signal_7804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3327 ( .C ( clk ), .D ( n2050 ), .Q ( new_AGEMA_signal_7816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3333 ( .C ( clk ), .D ( new_AGEMA_signal_1400 ), .Q ( new_AGEMA_signal_7822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3339 ( .C ( clk ), .D ( new_AGEMA_signal_1401 ), .Q ( new_AGEMA_signal_7828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3359 ( .C ( clk ), .D ( new_AGEMA_signal_7847 ), .Q ( new_AGEMA_signal_7848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3367 ( .C ( clk ), .D ( new_AGEMA_signal_7855 ), .Q ( new_AGEMA_signal_7856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3375 ( .C ( clk ), .D ( new_AGEMA_signal_7863 ), .Q ( new_AGEMA_signal_7864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3393 ( .C ( clk ), .D ( n2183 ), .Q ( new_AGEMA_signal_7882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3399 ( .C ( clk ), .D ( new_AGEMA_signal_1230 ), .Q ( new_AGEMA_signal_7888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3405 ( .C ( clk ), .D ( new_AGEMA_signal_1231 ), .Q ( new_AGEMA_signal_7894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3411 ( .C ( clk ), .D ( n2196 ), .Q ( new_AGEMA_signal_7900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3417 ( .C ( clk ), .D ( new_AGEMA_signal_1476 ), .Q ( new_AGEMA_signal_7906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3423 ( .C ( clk ), .D ( new_AGEMA_signal_1477 ), .Q ( new_AGEMA_signal_7912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3429 ( .C ( clk ), .D ( n2238 ), .Q ( new_AGEMA_signal_7918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3435 ( .C ( clk ), .D ( new_AGEMA_signal_1490 ), .Q ( new_AGEMA_signal_7924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3441 ( .C ( clk ), .D ( new_AGEMA_signal_1491 ), .Q ( new_AGEMA_signal_7930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3447 ( .C ( clk ), .D ( n2249 ), .Q ( new_AGEMA_signal_7936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3453 ( .C ( clk ), .D ( new_AGEMA_signal_1822 ), .Q ( new_AGEMA_signal_7942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3459 ( .C ( clk ), .D ( new_AGEMA_signal_1823 ), .Q ( new_AGEMA_signal_7948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3465 ( .C ( clk ), .D ( n2273 ), .Q ( new_AGEMA_signal_7954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3471 ( .C ( clk ), .D ( new_AGEMA_signal_2106 ), .Q ( new_AGEMA_signal_7960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3477 ( .C ( clk ), .D ( new_AGEMA_signal_2107 ), .Q ( new_AGEMA_signal_7966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3497 ( .C ( clk ), .D ( new_AGEMA_signal_7985 ), .Q ( new_AGEMA_signal_7986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3505 ( .C ( clk ), .D ( new_AGEMA_signal_7993 ), .Q ( new_AGEMA_signal_7994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3513 ( .C ( clk ), .D ( new_AGEMA_signal_8001 ), .Q ( new_AGEMA_signal_8002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3531 ( .C ( clk ), .D ( n2349 ), .Q ( new_AGEMA_signal_8020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3537 ( .C ( clk ), .D ( new_AGEMA_signal_1538 ), .Q ( new_AGEMA_signal_8026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3543 ( .C ( clk ), .D ( new_AGEMA_signal_1539 ), .Q ( new_AGEMA_signal_8032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3551 ( .C ( clk ), .D ( new_AGEMA_signal_8039 ), .Q ( new_AGEMA_signal_8040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3559 ( .C ( clk ), .D ( new_AGEMA_signal_8047 ), .Q ( new_AGEMA_signal_8048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3567 ( .C ( clk ), .D ( new_AGEMA_signal_8055 ), .Q ( new_AGEMA_signal_8056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3579 ( .C ( clk ), .D ( n2396 ), .Q ( new_AGEMA_signal_8068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3585 ( .C ( clk ), .D ( new_AGEMA_signal_1560 ), .Q ( new_AGEMA_signal_8074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3591 ( .C ( clk ), .D ( new_AGEMA_signal_1561 ), .Q ( new_AGEMA_signal_8080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3609 ( .C ( clk ), .D ( n2439 ), .Q ( new_AGEMA_signal_8098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3615 ( .C ( clk ), .D ( new_AGEMA_signal_1892 ), .Q ( new_AGEMA_signal_8104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3621 ( .C ( clk ), .D ( new_AGEMA_signal_1893 ), .Q ( new_AGEMA_signal_8110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3627 ( .C ( clk ), .D ( n2470 ), .Q ( new_AGEMA_signal_8116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3633 ( .C ( clk ), .D ( new_AGEMA_signal_1580 ), .Q ( new_AGEMA_signal_8122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3639 ( .C ( clk ), .D ( new_AGEMA_signal_1581 ), .Q ( new_AGEMA_signal_8128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3647 ( .C ( clk ), .D ( new_AGEMA_signal_8135 ), .Q ( new_AGEMA_signal_8136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3655 ( .C ( clk ), .D ( new_AGEMA_signal_8143 ), .Q ( new_AGEMA_signal_8144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3663 ( .C ( clk ), .D ( new_AGEMA_signal_8151 ), .Q ( new_AGEMA_signal_8152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3671 ( .C ( clk ), .D ( new_AGEMA_signal_8159 ), .Q ( new_AGEMA_signal_8160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3679 ( .C ( clk ), .D ( new_AGEMA_signal_8167 ), .Q ( new_AGEMA_signal_8168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3687 ( .C ( clk ), .D ( new_AGEMA_signal_8175 ), .Q ( new_AGEMA_signal_8176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3693 ( .C ( clk ), .D ( n2585 ), .Q ( new_AGEMA_signal_8182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3699 ( .C ( clk ), .D ( new_AGEMA_signal_1940 ), .Q ( new_AGEMA_signal_8188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3705 ( .C ( clk ), .D ( new_AGEMA_signal_1941 ), .Q ( new_AGEMA_signal_8194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3711 ( .C ( clk ), .D ( n2607 ), .Q ( new_AGEMA_signal_8200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3717 ( .C ( clk ), .D ( new_AGEMA_signal_1616 ), .Q ( new_AGEMA_signal_8206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3723 ( .C ( clk ), .D ( new_AGEMA_signal_1617 ), .Q ( new_AGEMA_signal_8212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3813 ( .C ( clk ), .D ( n2013 ), .Q ( new_AGEMA_signal_8302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3821 ( .C ( clk ), .D ( new_AGEMA_signal_1728 ), .Q ( new_AGEMA_signal_8310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3829 ( .C ( clk ), .D ( new_AGEMA_signal_1729 ), .Q ( new_AGEMA_signal_8318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3837 ( .C ( clk ), .D ( n2028 ), .Q ( new_AGEMA_signal_8326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3845 ( .C ( clk ), .D ( new_AGEMA_signal_1200 ), .Q ( new_AGEMA_signal_8334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3853 ( .C ( clk ), .D ( new_AGEMA_signal_1201 ), .Q ( new_AGEMA_signal_8342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3861 ( .C ( clk ), .D ( n2051 ), .Q ( new_AGEMA_signal_8350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3869 ( .C ( clk ), .D ( new_AGEMA_signal_1740 ), .Q ( new_AGEMA_signal_8358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3877 ( .C ( clk ), .D ( new_AGEMA_signal_1741 ), .Q ( new_AGEMA_signal_8366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3885 ( .C ( clk ), .D ( n2069 ), .Q ( new_AGEMA_signal_8374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3893 ( .C ( clk ), .D ( new_AGEMA_signal_1750 ), .Q ( new_AGEMA_signal_8382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3901 ( .C ( clk ), .D ( new_AGEMA_signal_1751 ), .Q ( new_AGEMA_signal_8390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3929 ( .C ( clk ), .D ( new_AGEMA_signal_8417 ), .Q ( new_AGEMA_signal_8418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3939 ( .C ( clk ), .D ( new_AGEMA_signal_8427 ), .Q ( new_AGEMA_signal_8428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3949 ( .C ( clk ), .D ( new_AGEMA_signal_8437 ), .Q ( new_AGEMA_signal_8438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3957 ( .C ( clk ), .D ( n2144 ), .Q ( new_AGEMA_signal_8446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3965 ( .C ( clk ), .D ( new_AGEMA_signal_1784 ), .Q ( new_AGEMA_signal_8454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3973 ( .C ( clk ), .D ( new_AGEMA_signal_1785 ), .Q ( new_AGEMA_signal_8462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3981 ( .C ( clk ), .D ( n2170 ), .Q ( new_AGEMA_signal_8470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3989 ( .C ( clk ), .D ( new_AGEMA_signal_1788 ), .Q ( new_AGEMA_signal_8478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3997 ( .C ( clk ), .D ( new_AGEMA_signal_1789 ), .Q ( new_AGEMA_signal_8486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4005 ( .C ( clk ), .D ( n2186 ), .Q ( new_AGEMA_signal_8494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4013 ( .C ( clk ), .D ( new_AGEMA_signal_1226 ), .Q ( new_AGEMA_signal_8502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4021 ( .C ( clk ), .D ( new_AGEMA_signal_1227 ), .Q ( new_AGEMA_signal_8510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4079 ( .C ( clk ), .D ( new_AGEMA_signal_8567 ), .Q ( new_AGEMA_signal_8568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4089 ( .C ( clk ), .D ( new_AGEMA_signal_8577 ), .Q ( new_AGEMA_signal_8578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4099 ( .C ( clk ), .D ( new_AGEMA_signal_8587 ), .Q ( new_AGEMA_signal_8588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4107 ( .C ( clk ), .D ( new_AGEMA_signal_6329 ), .Q ( new_AGEMA_signal_8596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4115 ( .C ( clk ), .D ( new_AGEMA_signal_6331 ), .Q ( new_AGEMA_signal_8604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4123 ( .C ( clk ), .D ( new_AGEMA_signal_6333 ), .Q ( new_AGEMA_signal_8612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4149 ( .C ( clk ), .D ( n2551 ), .Q ( new_AGEMA_signal_8638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4157 ( .C ( clk ), .D ( new_AGEMA_signal_1928 ), .Q ( new_AGEMA_signal_8646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4165 ( .C ( clk ), .D ( new_AGEMA_signal_1929 ), .Q ( new_AGEMA_signal_8654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4173 ( .C ( clk ), .D ( n2588 ), .Q ( new_AGEMA_signal_8662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4181 ( .C ( clk ), .D ( new_AGEMA_signal_1946 ), .Q ( new_AGEMA_signal_8670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4189 ( .C ( clk ), .D ( new_AGEMA_signal_1947 ), .Q ( new_AGEMA_signal_8678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4227 ( .C ( clk ), .D ( n2701 ), .Q ( new_AGEMA_signal_8716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4235 ( .C ( clk ), .D ( new_AGEMA_signal_1644 ), .Q ( new_AGEMA_signal_8724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4243 ( .C ( clk ), .D ( new_AGEMA_signal_1645 ), .Q ( new_AGEMA_signal_8732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4425 ( .C ( clk ), .D ( n2172 ), .Q ( new_AGEMA_signal_8914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4435 ( .C ( clk ), .D ( new_AGEMA_signal_1794 ), .Q ( new_AGEMA_signal_8924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4445 ( .C ( clk ), .D ( new_AGEMA_signal_1795 ), .Q ( new_AGEMA_signal_8934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5013 ( .C ( clk ), .D ( n2150 ), .Q ( new_AGEMA_signal_9502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5027 ( .C ( clk ), .D ( new_AGEMA_signal_1452 ), .Q ( new_AGEMA_signal_9516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5041 ( .C ( clk ), .D ( new_AGEMA_signal_1453 ), .Q ( new_AGEMA_signal_9530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5079 ( .C ( clk ), .D ( n2369 ), .Q ( new_AGEMA_signal_9568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5093 ( .C ( clk ), .D ( new_AGEMA_signal_2138 ), .Q ( new_AGEMA_signal_9582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5107 ( .C ( clk ), .D ( new_AGEMA_signal_2139 ), .Q ( new_AGEMA_signal_9596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5187 ( .C ( clk ), .D ( n2152 ), .Q ( new_AGEMA_signal_9676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5203 ( .C ( clk ), .D ( new_AGEMA_signal_1786 ), .Q ( new_AGEMA_signal_9692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5219 ( .C ( clk ), .D ( new_AGEMA_signal_1787 ), .Q ( new_AGEMA_signal_9708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5253 ( .C ( clk ), .D ( n2372 ), .Q ( new_AGEMA_signal_9742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5269 ( .C ( clk ), .D ( new_AGEMA_signal_1866 ), .Q ( new_AGEMA_signal_9758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5285 ( .C ( clk ), .D ( new_AGEMA_signal_1867 ), .Q ( new_AGEMA_signal_9774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5481 ( .C ( clk ), .D ( n2375 ), .Q ( new_AGEMA_signal_9970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5499 ( .C ( clk ), .D ( new_AGEMA_signal_1540 ), .Q ( new_AGEMA_signal_9988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5517 ( .C ( clk ), .D ( new_AGEMA_signal_1541 ), .Q ( new_AGEMA_signal_10006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5631 ( .C ( clk ), .D ( n2377 ), .Q ( new_AGEMA_signal_10120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5651 ( .C ( clk ), .D ( new_AGEMA_signal_1868 ), .Q ( new_AGEMA_signal_10140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5671 ( .C ( clk ), .D ( new_AGEMA_signal_1869 ), .Q ( new_AGEMA_signal_10160 ) ) ;

    /* cells in depth 8 */
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1968 ( .a ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, n1924}), .b ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, n1923}), .clk ( clk ), .r ({Fresh[1355], Fresh[1354], Fresh[1353]}), .c ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, n1936}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1982 ( .a ({new_AGEMA_signal_5919, new_AGEMA_signal_5917, new_AGEMA_signal_5915}), .b ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, n1927}), .clk ( clk ), .r ({Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, n1928}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U1994 ( .a ({new_AGEMA_signal_5925, new_AGEMA_signal_5923, new_AGEMA_signal_5921}), .b ({new_AGEMA_signal_1683, new_AGEMA_signal_1682, n1929}), .clk ( clk ), .r ({Fresh[1361], Fresh[1360], Fresh[1359]}), .c ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, n1931}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2012 ( .a ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, n2665}), .b ({new_AGEMA_signal_1687, new_AGEMA_signal_1686, n1938}), .clk ( clk ), .r ({Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, n1939}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2024 ( .a ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, n2235}), .b ({new_AGEMA_signal_1333, new_AGEMA_signal_1332, n1943}), .clk ( clk ), .r ({Fresh[1367], Fresh[1366], Fresh[1365]}), .c ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, n1948}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2032 ( .a ({new_AGEMA_signal_1335, new_AGEMA_signal_1334, n1946}), .b ({new_AGEMA_signal_1691, new_AGEMA_signal_1690, n1945}), .clk ( clk ), .r ({Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, n1947}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2041 ( .a ({new_AGEMA_signal_5937, new_AGEMA_signal_5933, new_AGEMA_signal_5929}), .b ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, n1951}), .clk ( clk ), .r ({Fresh[1373], Fresh[1372], Fresh[1371]}), .c ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, n1954}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2049 ( .a ({new_AGEMA_signal_5943, new_AGEMA_signal_5941, new_AGEMA_signal_5939}), .b ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, n1952}), .clk ( clk ), .r ({Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, n1953}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2058 ( .a ({new_AGEMA_signal_5949, new_AGEMA_signal_5947, new_AGEMA_signal_5945}), .b ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, n2687}), .clk ( clk ), .r ({Fresh[1379], Fresh[1378], Fresh[1377]}), .c ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, n2658}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2065 ( .a ({new_AGEMA_signal_5955, new_AGEMA_signal_5953, new_AGEMA_signal_5951}), .b ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, n1963}), .clk ( clk ), .r ({Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, n1965}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2078 ( .a ({new_AGEMA_signal_5961, new_AGEMA_signal_5959, new_AGEMA_signal_5957}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, n1968}), .clk ( clk ), .r ({Fresh[1385], Fresh[1384], Fresh[1383]}), .c ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, n1970}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2084 ( .a ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, n2684}), .b ({new_AGEMA_signal_5967, new_AGEMA_signal_5965, new_AGEMA_signal_5963}), .clk ( clk ), .r ({Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, n1969}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2093 ( .a ({new_AGEMA_signal_1711, new_AGEMA_signal_1710, n1972}), .b ({new_AGEMA_signal_1357, new_AGEMA_signal_1356, n1971}), .clk ( clk ), .r ({Fresh[1391], Fresh[1390], Fresh[1389]}), .c ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, n1978}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2102 ( .a ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, n1974}), .b ({new_AGEMA_signal_5973, new_AGEMA_signal_5971, new_AGEMA_signal_5969}), .clk ( clk ), .r ({Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, n1975}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2107 ( .a ({new_AGEMA_signal_5979, new_AGEMA_signal_5977, new_AGEMA_signal_5975}), .b ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, n1979}), .clk ( clk ), .r ({Fresh[1397], Fresh[1396], Fresh[1395]}), .c ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, n1980}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2114 ( .a ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, n1985}), .b ({new_AGEMA_signal_5985, new_AGEMA_signal_5983, new_AGEMA_signal_5981}), .clk ( clk ), .r ({Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, n1986}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2124 ( .a ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, n1994}), .b ({new_AGEMA_signal_5991, new_AGEMA_signal_5989, new_AGEMA_signal_5987}), .clk ( clk ), .r ({Fresh[1403], Fresh[1402], Fresh[1401]}), .c ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, n1997}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2137 ( .a ({new_AGEMA_signal_5997, new_AGEMA_signal_5995, new_AGEMA_signal_5993}), .b ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, n2137}), .clk ( clk ), .r ({Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, n2012}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2145 ( .a ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, n2006}), .b ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, n2005}), .clk ( clk ), .r ({Fresh[1409], Fresh[1408], Fresh[1407]}), .c ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, n2007}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) U2161 ( .s ({new_AGEMA_signal_6003, new_AGEMA_signal_6001, new_AGEMA_signal_5999}), .b ({new_AGEMA_signal_1389, new_AGEMA_signal_1388, n2020}), .a ({new_AGEMA_signal_6015, new_AGEMA_signal_6011, new_AGEMA_signal_6007}), .clk ( clk ), .r ({Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, n2021}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2176 ( .a ({new_AGEMA_signal_6021, new_AGEMA_signal_6019, new_AGEMA_signal_6017}), .b ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, n2031}), .clk ( clk ), .r ({Fresh[1415], Fresh[1414], Fresh[1413]}), .c ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, n2032}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2185 ( .a ({new_AGEMA_signal_6027, new_AGEMA_signal_6025, new_AGEMA_signal_6023}), .b ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, n2040}), .clk ( clk ), .r ({Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, n2041}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2189 ( .a ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, n2665}), .b ({new_AGEMA_signal_6033, new_AGEMA_signal_6031, new_AGEMA_signal_6029}), .clk ( clk ), .r ({Fresh[1421], Fresh[1420], Fresh[1419]}), .c ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, n2043}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2194 ( .a ({new_AGEMA_signal_6039, new_AGEMA_signal_6037, new_AGEMA_signal_6035}), .b ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, n2045}), .clk ( clk ), .r ({Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, n2046}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) U2204 ( .s ({new_AGEMA_signal_6003, new_AGEMA_signal_6001, new_AGEMA_signal_5999}), .b ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, n2056}), .a ({new_AGEMA_signal_6045, new_AGEMA_signal_6043, new_AGEMA_signal_6041}), .clk ( clk ), .r ({Fresh[1427], Fresh[1426], Fresh[1425]}), .c ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, n2058}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2210 ( .a ({new_AGEMA_signal_6051, new_AGEMA_signal_6049, new_AGEMA_signal_6047}), .b ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, n2060}), .clk ( clk ), .r ({Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, n2063}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2218 ( .a ({new_AGEMA_signal_1747, new_AGEMA_signal_1746, n2066}), .b ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, n2065}), .clk ( clk ), .r ({Fresh[1433], Fresh[1432], Fresh[1431]}), .c ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, n2652}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2227 ( .a ({new_AGEMA_signal_6057, new_AGEMA_signal_6055, new_AGEMA_signal_6053}), .b ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, n2074}), .clk ( clk ), .r ({Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, n2076}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2236 ( .a ({new_AGEMA_signal_6069, new_AGEMA_signal_6065, new_AGEMA_signal_6061}), .b ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, n2082}), .clk ( clk ), .r ({Fresh[1439], Fresh[1438], Fresh[1437]}), .c ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, n2105}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2241 ( .a ({new_AGEMA_signal_6075, new_AGEMA_signal_6073, new_AGEMA_signal_6071}), .b ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, n2084}), .clk ( clk ), .r ({Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, n2099}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2243 ( .a ({new_AGEMA_signal_1759, new_AGEMA_signal_1758, n2085}), .b ({new_AGEMA_signal_6081, new_AGEMA_signal_6079, new_AGEMA_signal_6077}), .clk ( clk ), .r ({Fresh[1445], Fresh[1444], Fresh[1443]}), .c ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, n2091}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) U2246 ( .a ({new_AGEMA_signal_6087, new_AGEMA_signal_6085, new_AGEMA_signal_6083}), .b ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, n2131}), .clk ( clk ), .r ({Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, n2090}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2253 ( .a ({new_AGEMA_signal_6093, new_AGEMA_signal_6091, new_AGEMA_signal_6089}), .b ({new_AGEMA_signal_1765, new_AGEMA_signal_1764, n2330}), .clk ( clk ), .r ({Fresh[1451], Fresh[1450], Fresh[1449]}), .c ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, n2093}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2262 ( .a ({new_AGEMA_signal_6099, new_AGEMA_signal_6097, new_AGEMA_signal_6095}), .b ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, n2160}), .clk ( clk ), .r ({Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, n2102}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2266 ( .a ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, n2504}), .b ({new_AGEMA_signal_6111, new_AGEMA_signal_6107, new_AGEMA_signal_6103}), .clk ( clk ), .r ({Fresh[1457], Fresh[1456], Fresh[1455]}), .c ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, n2106}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2272 ( .a ({new_AGEMA_signal_6117, new_AGEMA_signal_6115, new_AGEMA_signal_6113}), .b ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, n2114}), .clk ( clk ), .r ({Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, n2116}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2282 ( .a ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, n2291}), .b ({new_AGEMA_signal_1443, new_AGEMA_signal_1442, n2119}), .clk ( clk ), .r ({Fresh[1463], Fresh[1462], Fresh[1461]}), .c ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, n2120}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2293 ( .a ({new_AGEMA_signal_1449, new_AGEMA_signal_1448, n2130}), .b ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, n2129}), .clk ( clk ), .r ({Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({new_AGEMA_signal_1777, new_AGEMA_signal_1776, n2155}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2296 ( .a ({new_AGEMA_signal_6123, new_AGEMA_signal_6121, new_AGEMA_signal_6119}), .b ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, n2131}), .clk ( clk ), .r ({Fresh[1469], Fresh[1468], Fresh[1467]}), .c ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, n2543}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2299 ( .a ({new_AGEMA_signal_1455, new_AGEMA_signal_1454, n2133}), .b ({new_AGEMA_signal_6129, new_AGEMA_signal_6127, new_AGEMA_signal_6125}), .clk ( clk ), .r ({Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, n2134}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2303 ( .a ({new_AGEMA_signal_1723, new_AGEMA_signal_1722, n2137}), .b ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, n2136}), .clk ( clk ), .r ({Fresh[1475], Fresh[1474], Fresh[1473]}), .c ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, n2143}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2308 ( .a ({new_AGEMA_signal_1783, new_AGEMA_signal_1782, n2139}), .b ({new_AGEMA_signal_6141, new_AGEMA_signal_6137, new_AGEMA_signal_6133}), .clk ( clk ), .r ({Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, n2140}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2324 ( .a ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, n2157}), .b ({new_AGEMA_signal_6147, new_AGEMA_signal_6145, new_AGEMA_signal_6143}), .clk ( clk ), .r ({Fresh[1481], Fresh[1480], Fresh[1479]}), .c ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, n2159}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2326 ( .a ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, n2160}), .b ({new_AGEMA_signal_6153, new_AGEMA_signal_6151, new_AGEMA_signal_6149}), .clk ( clk ), .r ({Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, n2161}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2330 ( .a ({new_AGEMA_signal_5937, new_AGEMA_signal_5933, new_AGEMA_signal_5929}), .b ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, n2163}), .clk ( clk ), .r ({Fresh[1487], Fresh[1486], Fresh[1485]}), .c ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, n2164}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2345 ( .a ({new_AGEMA_signal_6159, new_AGEMA_signal_6157, new_AGEMA_signal_6155}), .b ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, n2177}), .clk ( clk ), .r ({Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, n2179}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2359 ( .a ({new_AGEMA_signal_6171, new_AGEMA_signal_6167, new_AGEMA_signal_6163}), .b ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, n2191}), .clk ( clk ), .r ({Fresh[1493], Fresh[1492], Fresh[1491]}), .c ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, n2192}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2370 ( .a ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, n2201}), .b ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2200}), .clk ( clk ), .r ({Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, n2203}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2382 ( .a ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, n2217}), .b ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, n2216}), .clk ( clk ), .r ({Fresh[1499], Fresh[1498], Fresh[1497]}), .c ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, n2224}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2388 ( .a ({new_AGEMA_signal_1813, new_AGEMA_signal_1812, n2222}), .b ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, n2221}), .clk ( clk ), .r ({Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, n2223}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2392 ( .a ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, n2504}), .b ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, n2226}), .clk ( clk ), .r ({Fresh[1505], Fresh[1504], Fresh[1503]}), .c ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, n2229}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2399 ( .a ({new_AGEMA_signal_5943, new_AGEMA_signal_5941, new_AGEMA_signal_5939}), .b ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, n2233}), .clk ( clk ), .r ({Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, n2234}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2410 ( .a ({new_AGEMA_signal_5949, new_AGEMA_signal_5947, new_AGEMA_signal_5945}), .b ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, n2244}), .clk ( clk ), .r ({Fresh[1511], Fresh[1510], Fresh[1509]}), .c ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, n2246}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2418 ( .a ({new_AGEMA_signal_6177, new_AGEMA_signal_6175, new_AGEMA_signal_6173}), .b ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, n2253}), .clk ( clk ), .r ({Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, n2254}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2425 ( .a ({new_AGEMA_signal_6183, new_AGEMA_signal_6181, new_AGEMA_signal_6179}), .b ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, n2260}), .clk ( clk ), .r ({Fresh[1517], Fresh[1516], Fresh[1515]}), .c ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, n2263}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2434 ( .a ({new_AGEMA_signal_6189, new_AGEMA_signal_6187, new_AGEMA_signal_6185}), .b ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, n2265}), .clk ( clk ), .r ({Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, n2267}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2438 ( .a ({new_AGEMA_signal_5943, new_AGEMA_signal_5941, new_AGEMA_signal_5939}), .b ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, n2269}), .clk ( clk ), .r ({Fresh[1523], Fresh[1522], Fresh[1521]}), .c ({new_AGEMA_signal_1831, new_AGEMA_signal_1830, n2270}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2445 ( .a ({new_AGEMA_signal_6195, new_AGEMA_signal_6193, new_AGEMA_signal_6191}), .b ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, n2277}), .clk ( clk ), .r ({Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, n2279}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2450 ( .a ({new_AGEMA_signal_6015, new_AGEMA_signal_6011, new_AGEMA_signal_6007}), .b ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, n2282}), .clk ( clk ), .r ({Fresh[1529], Fresh[1528], Fresh[1527]}), .c ({new_AGEMA_signal_1835, new_AGEMA_signal_1834, n2283}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2453 ( .a ({new_AGEMA_signal_6075, new_AGEMA_signal_6073, new_AGEMA_signal_6071}), .b ({new_AGEMA_signal_1837, new_AGEMA_signal_1836, n2284}), .clk ( clk ), .r ({Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, n2285}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2457 ( .a ({new_AGEMA_signal_5937, new_AGEMA_signal_5933, new_AGEMA_signal_5929}), .b ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, n2459}), .clk ( clk ), .r ({Fresh[1535], Fresh[1534], Fresh[1533]}), .c ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, n2686}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2460 ( .a ({new_AGEMA_signal_5949, new_AGEMA_signal_5947, new_AGEMA_signal_5945}), .b ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, n2288}), .clk ( clk ), .r ({Fresh[1538], Fresh[1537], Fresh[1536]}), .c ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, n2289}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2463 ( .a ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, n2458}), .b ({new_AGEMA_signal_6201, new_AGEMA_signal_6199, new_AGEMA_signal_6197}), .clk ( clk ), .r ({Fresh[1541], Fresh[1540], Fresh[1539]}), .c ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, n2297}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2465 ( .a ({new_AGEMA_signal_6207, new_AGEMA_signal_6205, new_AGEMA_signal_6203}), .b ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, n2291}), .clk ( clk ), .r ({Fresh[1544], Fresh[1543], Fresh[1542]}), .c ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, n2292}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2473 ( .a ({new_AGEMA_signal_6213, new_AGEMA_signal_6211, new_AGEMA_signal_6209}), .b ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, n2300}), .clk ( clk ), .r ({Fresh[1547], Fresh[1546], Fresh[1545]}), .c ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, n2301}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2483 ( .a ({new_AGEMA_signal_6219, new_AGEMA_signal_6217, new_AGEMA_signal_6215}), .b ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, n2314}), .clk ( clk ), .r ({Fresh[1550], Fresh[1549], Fresh[1548]}), .c ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, n2321}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2487 ( .a ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, n2319}), .b ({new_AGEMA_signal_6225, new_AGEMA_signal_6223, new_AGEMA_signal_6221}), .clk ( clk ), .r ({Fresh[1553], Fresh[1552], Fresh[1551]}), .c ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, n2320}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2493 ( .a ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, n2326}), .b ({new_AGEMA_signal_6231, new_AGEMA_signal_6229, new_AGEMA_signal_6227}), .clk ( clk ), .r ({Fresh[1556], Fresh[1555], Fresh[1554]}), .c ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, n2334}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2497 ( .a ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, n2329}), .b ({new_AGEMA_signal_6015, new_AGEMA_signal_6011, new_AGEMA_signal_6007}), .clk ( clk ), .r ({Fresh[1559], Fresh[1558], Fresh[1557]}), .c ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, n2332}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2498 ( .a ({new_AGEMA_signal_6237, new_AGEMA_signal_6235, new_AGEMA_signal_6233}), .b ({new_AGEMA_signal_1765, new_AGEMA_signal_1764, n2330}), .clk ( clk ), .r ({Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, n2331}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2502 ( .a ({new_AGEMA_signal_6243, new_AGEMA_signal_6241, new_AGEMA_signal_6239}), .b ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, n2335}), .clk ( clk ), .r ({Fresh[1565], Fresh[1564], Fresh[1563]}), .c ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, n2336}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2508 ( .a ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, n2341}), .b ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, n2340}), .clk ( clk ), .r ({Fresh[1568], Fresh[1567], Fresh[1566]}), .c ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, n2342}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2519 ( .a ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, n2352}), .b ({new_AGEMA_signal_6249, new_AGEMA_signal_6247, new_AGEMA_signal_6245}), .clk ( clk ), .r ({Fresh[1571], Fresh[1570], Fresh[1569]}), .c ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, n2367}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2523 ( .a ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, n2354}), .b ({new_AGEMA_signal_6255, new_AGEMA_signal_6253, new_AGEMA_signal_6251}), .clk ( clk ), .r ({Fresh[1574], Fresh[1573], Fresh[1572]}), .c ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, n2358}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2547 ( .a ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, n2385}), .b ({new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2384}), .clk ( clk ), .r ({Fresh[1577], Fresh[1576], Fresh[1575]}), .c ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, n2387}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2555 ( .a ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, n2391}), .b ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, n2390}), .clk ( clk ), .r ({Fresh[1580], Fresh[1579], Fresh[1578]}), .c ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, n2392}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2566 ( .a ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, n2403}), .b ({new_AGEMA_signal_6261, new_AGEMA_signal_6259, new_AGEMA_signal_6257}), .clk ( clk ), .r ({Fresh[1583], Fresh[1582], Fresh[1581]}), .c ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, n2404}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2570 ( .a ({new_AGEMA_signal_6051, new_AGEMA_signal_6049, new_AGEMA_signal_6047}), .b ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, n2408}), .clk ( clk ), .r ({Fresh[1586], Fresh[1585], Fresh[1584]}), .c ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, n2409}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2575 ( .a ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, n2574}), .b ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, n2413}), .clk ( clk ), .r ({Fresh[1589], Fresh[1588], Fresh[1587]}), .c ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, n2414}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2578 ( .a ({new_AGEMA_signal_6267, new_AGEMA_signal_6265, new_AGEMA_signal_6263}), .b ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, n2416}), .clk ( clk ), .r ({Fresh[1592], Fresh[1591], Fresh[1590]}), .c ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, n2418}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2589 ( .a ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, n2689}), .b ({new_AGEMA_signal_6273, new_AGEMA_signal_6271, new_AGEMA_signal_6269}), .clk ( clk ), .r ({Fresh[1595], Fresh[1594], Fresh[1593]}), .c ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, n2432}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2592 ( .a ({new_AGEMA_signal_6291, new_AGEMA_signal_6285, new_AGEMA_signal_6279}), .b ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, n2434}), .clk ( clk ), .r ({Fresh[1598], Fresh[1597], Fresh[1596]}), .c ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, n2435}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2601 ( .a ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, n2445}), .b ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, n2444}), .clk ( clk ), .r ({Fresh[1601], Fresh[1600], Fresh[1599]}), .c ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, n2449}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2603 ( .a ({new_AGEMA_signal_6219, new_AGEMA_signal_6217, new_AGEMA_signal_6215}), .b ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, n2447}), .clk ( clk ), .r ({Fresh[1604], Fresh[1603], Fresh[1602]}), .c ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, n2448}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2609 ( .a ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, n2454}), .b ({new_AGEMA_signal_6297, new_AGEMA_signal_6295, new_AGEMA_signal_6293}), .clk ( clk ), .r ({Fresh[1607], Fresh[1606], Fresh[1605]}), .c ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, n2455}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2612 ( .a ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, n2687}), .b ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, n2458}), .clk ( clk ), .r ({Fresh[1610], Fresh[1609], Fresh[1608]}), .c ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, n2460}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2618 ( .a ({new_AGEMA_signal_6207, new_AGEMA_signal_6205, new_AGEMA_signal_6203}), .b ({new_AGEMA_signal_1579, new_AGEMA_signal_1578, n2465}), .clk ( clk ), .r ({Fresh[1613], Fresh[1612], Fresh[1611]}), .c ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, n2466}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2629 ( .a ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, n2476}), .b ({new_AGEMA_signal_6303, new_AGEMA_signal_6301, new_AGEMA_signal_6299}), .clk ( clk ), .r ({Fresh[1616], Fresh[1615], Fresh[1614]}), .c ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, n2477}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2634 ( .a ({new_AGEMA_signal_6045, new_AGEMA_signal_6043, new_AGEMA_signal_6041}), .b ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, n2481}), .clk ( clk ), .r ({Fresh[1619], Fresh[1618], Fresh[1617]}), .c ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, n2482}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2640 ( .a ({new_AGEMA_signal_6309, new_AGEMA_signal_6307, new_AGEMA_signal_6305}), .b ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, n2486}), .clk ( clk ), .r ({Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, n2490}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2648 ( .a ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, n2495}), .b ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, n2494}), .clk ( clk ), .r ({Fresh[1625], Fresh[1624], Fresh[1623]}), .c ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, n2496}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2654 ( .a ({new_AGEMA_signal_1437, new_AGEMA_signal_1436, n2504}), .b ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, n2503}), .clk ( clk ), .r ({Fresh[1628], Fresh[1627], Fresh[1626]}), .c ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, n2507}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2664 ( .a ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, n2518}), .b ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, n2517}), .clk ( clk ), .r ({Fresh[1631], Fresh[1630], Fresh[1629]}), .c ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, n2525}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2669 ( .a ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, n2523}), .b ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, n2522}), .clk ( clk ), .r ({Fresh[1634], Fresh[1633], Fresh[1632]}), .c ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, n2524}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2676 ( .a ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, n2532}), .b ({new_AGEMA_signal_6321, new_AGEMA_signal_6317, new_AGEMA_signal_6313}), .clk ( clk ), .r ({Fresh[1637], Fresh[1636], Fresh[1635]}), .c ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, n2537}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2678 ( .a ({new_AGEMA_signal_6051, new_AGEMA_signal_6049, new_AGEMA_signal_6047}), .b ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, n2534}), .clk ( clk ), .r ({Fresh[1640], Fresh[1639], Fresh[1638]}), .c ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, n2536}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2684 ( .a ({new_AGEMA_signal_6327, new_AGEMA_signal_6325, new_AGEMA_signal_6323}), .b ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, n2546}), .clk ( clk ), .r ({Fresh[1643], Fresh[1642], Fresh[1641]}), .c ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, n2547}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2693 ( .a ({new_AGEMA_signal_6333, new_AGEMA_signal_6331, new_AGEMA_signal_6329}), .b ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, n2556}), .clk ( clk ), .r ({Fresh[1646], Fresh[1645], Fresh[1644]}), .c ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, n2557}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2699 ( .a ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, n2715}), .b ({new_AGEMA_signal_6339, new_AGEMA_signal_6337, new_AGEMA_signal_6335}), .clk ( clk ), .r ({Fresh[1649], Fresh[1648], Fresh[1647]}), .c ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, n2565}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2704 ( .a ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, n2574}), .b ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, n2573}), .clk ( clk ), .r ({Fresh[1652], Fresh[1651], Fresh[1650]}), .c ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, n2591}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2709 ( .a ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, n2579}), .b ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, n2578}), .clk ( clk ), .r ({Fresh[1655], Fresh[1654], Fresh[1653]}), .c ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, n2580}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2727 ( .a ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, n2601}), .b ({new_AGEMA_signal_6351, new_AGEMA_signal_6347, new_AGEMA_signal_6343}), .clk ( clk ), .r ({Fresh[1658], Fresh[1657], Fresh[1656]}), .c ({new_AGEMA_signal_1623, new_AGEMA_signal_1622, n2602}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2738 ( .a ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, n2618}), .b ({new_AGEMA_signal_6357, new_AGEMA_signal_6355, new_AGEMA_signal_6353}), .clk ( clk ), .r ({Fresh[1661], Fresh[1660], Fresh[1659]}), .c ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, n2619}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2744 ( .a ({new_AGEMA_signal_6081, new_AGEMA_signal_6079, new_AGEMA_signal_6077}), .b ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, n2626}), .clk ( clk ), .r ({Fresh[1664], Fresh[1663], Fresh[1662]}), .c ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, n2628}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2753 ( .a ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, n2644}), .b ({new_AGEMA_signal_6123, new_AGEMA_signal_6121, new_AGEMA_signal_6119}), .clk ( clk ), .r ({Fresh[1667], Fresh[1666], Fresh[1665]}), .c ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, n2649}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2755 ( .a ({new_AGEMA_signal_6363, new_AGEMA_signal_6361, new_AGEMA_signal_6359}), .b ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, n2646}), .clk ( clk ), .r ({Fresh[1670], Fresh[1669], Fresh[1668]}), .c ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, n2648}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2765 ( .a ({new_AGEMA_signal_5949, new_AGEMA_signal_5947, new_AGEMA_signal_5945}), .b ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, n2663}), .clk ( clk ), .r ({Fresh[1673], Fresh[1672], Fresh[1671]}), .c ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, n2664}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2771 ( .a ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, n2675}), .b ({new_AGEMA_signal_6369, new_AGEMA_signal_6367, new_AGEMA_signal_6365}), .clk ( clk ), .r ({Fresh[1676], Fresh[1675], Fresh[1674]}), .c ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, n2681}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2773 ( .a ({new_AGEMA_signal_6147, new_AGEMA_signal_6145, new_AGEMA_signal_6143}), .b ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, n2678}), .clk ( clk ), .r ({Fresh[1679], Fresh[1678], Fresh[1677]}), .c ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, n2680}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2776 ( .a ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, n2684}), .b ({new_AGEMA_signal_6375, new_AGEMA_signal_6373, new_AGEMA_signal_6371}), .clk ( clk ), .r ({Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, n2685}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2778 ( .a ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, n2687}), .b ({new_AGEMA_signal_6327, new_AGEMA_signal_6325, new_AGEMA_signal_6323}), .clk ( clk ), .r ({Fresh[1685], Fresh[1684], Fresh[1683]}), .c ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, n2698}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2779 ( .a ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, n2689}), .b ({new_AGEMA_signal_6333, new_AGEMA_signal_6331, new_AGEMA_signal_6329}), .clk ( clk ), .r ({Fresh[1688], Fresh[1687], Fresh[1686]}), .c ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, n2692}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2793 ( .a ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, n2715}), .b ({new_AGEMA_signal_6381, new_AGEMA_signal_6379, new_AGEMA_signal_6377}), .clk ( clk ), .r ({Fresh[1691], Fresh[1690], Fresh[1689]}), .c ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, n2716}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2800 ( .a ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, n2727}), .b ({new_AGEMA_signal_6387, new_AGEMA_signal_6385, new_AGEMA_signal_6383}), .clk ( clk ), .r ({Fresh[1694], Fresh[1693], Fresh[1692]}), .c ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, n2728}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2804 ( .a ({new_AGEMA_signal_6393, new_AGEMA_signal_6391, new_AGEMA_signal_6389}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, n2733}), .clk ( clk ), .r ({Fresh[1697], Fresh[1696], Fresh[1695]}), .c ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, n2735}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2808 ( .a ({new_AGEMA_signal_5985, new_AGEMA_signal_5983, new_AGEMA_signal_5981}), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, n2740}), .clk ( clk ), .r ({Fresh[1700], Fresh[1699], Fresh[1698]}), .c ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, n2743}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2813 ( .a ({new_AGEMA_signal_6405, new_AGEMA_signal_6401, new_AGEMA_signal_6397}), .b ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, n2749}), .clk ( clk ), .r ({Fresh[1703], Fresh[1702], Fresh[1701]}), .c ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, n2751}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2817 ( .a ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, n2757}), .b ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, n2756}), .clk ( clk ), .r ({Fresh[1706], Fresh[1705], Fresh[1704]}), .c ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, n2758}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2820 ( .a ({new_AGEMA_signal_6411, new_AGEMA_signal_6409, new_AGEMA_signal_6407}), .b ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, n2762}), .clk ( clk ), .r ({Fresh[1709], Fresh[1708], Fresh[1707]}), .c ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, n2764}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2827 ( .a ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, n2776}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, n2775}), .clk ( clk ), .r ({Fresh[1712], Fresh[1711], Fresh[1710]}), .c ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, n2800}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2831 ( .a ({new_AGEMA_signal_6417, new_AGEMA_signal_6415, new_AGEMA_signal_6413}), .b ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, n2783}), .clk ( clk ), .r ({Fresh[1715], Fresh[1714], Fresh[1713]}), .c ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, n2788}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2837 ( .a ({new_AGEMA_signal_6429, new_AGEMA_signal_6425, new_AGEMA_signal_6421}), .b ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, n2795}), .clk ( clk ), .r ({Fresh[1718], Fresh[1717], Fresh[1716]}), .c ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, n2797}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2846 ( .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, n2814}), .b ({new_AGEMA_signal_6003, new_AGEMA_signal_6001, new_AGEMA_signal_5999}), .clk ( clk ), .r ({Fresh[1721], Fresh[1720], Fresh[1719]}), .c ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, n2822}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2849 ( .a ({new_AGEMA_signal_6435, new_AGEMA_signal_6433, new_AGEMA_signal_6431}), .b ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, n2819}), .clk ( clk ), .r ({Fresh[1724], Fresh[1723], Fresh[1722]}), .c ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, n2821}) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C ( clk ), .D ( new_AGEMA_signal_6438 ), .Q ( new_AGEMA_signal_6439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C ( clk ), .D ( new_AGEMA_signal_6442 ), .Q ( new_AGEMA_signal_6443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C ( clk ), .D ( new_AGEMA_signal_6446 ), .Q ( new_AGEMA_signal_6447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C ( clk ), .D ( new_AGEMA_signal_6450 ), .Q ( new_AGEMA_signal_6451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C ( clk ), .D ( new_AGEMA_signal_6454 ), .Q ( new_AGEMA_signal_6455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C ( clk ), .D ( new_AGEMA_signal_6458 ), .Q ( new_AGEMA_signal_6459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C ( clk ), .D ( new_AGEMA_signal_6460 ), .Q ( new_AGEMA_signal_6461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C ( clk ), .D ( new_AGEMA_signal_6462 ), .Q ( new_AGEMA_signal_6463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C ( clk ), .D ( new_AGEMA_signal_6464 ), .Q ( new_AGEMA_signal_6465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C ( clk ), .D ( new_AGEMA_signal_6466 ), .Q ( new_AGEMA_signal_6467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C ( clk ), .D ( new_AGEMA_signal_6468 ), .Q ( new_AGEMA_signal_6469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C ( clk ), .D ( new_AGEMA_signal_6470 ), .Q ( new_AGEMA_signal_6471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C ( clk ), .D ( new_AGEMA_signal_6474 ), .Q ( new_AGEMA_signal_6475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C ( clk ), .D ( new_AGEMA_signal_6478 ), .Q ( new_AGEMA_signal_6479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C ( clk ), .D ( new_AGEMA_signal_6482 ), .Q ( new_AGEMA_signal_6483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C ( clk ), .D ( new_AGEMA_signal_6484 ), .Q ( new_AGEMA_signal_6485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C ( clk ), .D ( new_AGEMA_signal_6486 ), .Q ( new_AGEMA_signal_6487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C ( clk ), .D ( new_AGEMA_signal_6488 ), .Q ( new_AGEMA_signal_6489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C ( clk ), .D ( new_AGEMA_signal_6492 ), .Q ( new_AGEMA_signal_6493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C ( clk ), .D ( new_AGEMA_signal_6496 ), .Q ( new_AGEMA_signal_6497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C ( clk ), .D ( new_AGEMA_signal_6500 ), .Q ( new_AGEMA_signal_6501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C ( clk ), .D ( new_AGEMA_signal_6502 ), .Q ( new_AGEMA_signal_6503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C ( clk ), .D ( new_AGEMA_signal_6504 ), .Q ( new_AGEMA_signal_6505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C ( clk ), .D ( new_AGEMA_signal_6506 ), .Q ( new_AGEMA_signal_6507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C ( clk ), .D ( new_AGEMA_signal_6510 ), .Q ( new_AGEMA_signal_6511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C ( clk ), .D ( new_AGEMA_signal_6514 ), .Q ( new_AGEMA_signal_6515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C ( clk ), .D ( new_AGEMA_signal_6518 ), .Q ( new_AGEMA_signal_6519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C ( clk ), .D ( new_AGEMA_signal_6522 ), .Q ( new_AGEMA_signal_6523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C ( clk ), .D ( new_AGEMA_signal_6526 ), .Q ( new_AGEMA_signal_6527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C ( clk ), .D ( new_AGEMA_signal_6530 ), .Q ( new_AGEMA_signal_6531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C ( clk ), .D ( new_AGEMA_signal_6532 ), .Q ( new_AGEMA_signal_6533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C ( clk ), .D ( new_AGEMA_signal_6534 ), .Q ( new_AGEMA_signal_6535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C ( clk ), .D ( new_AGEMA_signal_6536 ), .Q ( new_AGEMA_signal_6537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C ( clk ), .D ( new_AGEMA_signal_6538 ), .Q ( new_AGEMA_signal_6539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C ( clk ), .D ( new_AGEMA_signal_6540 ), .Q ( new_AGEMA_signal_6541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C ( clk ), .D ( new_AGEMA_signal_6542 ), .Q ( new_AGEMA_signal_6543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C ( clk ), .D ( new_AGEMA_signal_6544 ), .Q ( new_AGEMA_signal_6545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C ( clk ), .D ( new_AGEMA_signal_6546 ), .Q ( new_AGEMA_signal_6547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C ( clk ), .D ( new_AGEMA_signal_6548 ), .Q ( new_AGEMA_signal_6549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C ( clk ), .D ( new_AGEMA_signal_6550 ), .Q ( new_AGEMA_signal_6551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C ( clk ), .D ( new_AGEMA_signal_6552 ), .Q ( new_AGEMA_signal_6553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C ( clk ), .D ( new_AGEMA_signal_6554 ), .Q ( new_AGEMA_signal_6555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C ( clk ), .D ( new_AGEMA_signal_6558 ), .Q ( new_AGEMA_signal_6559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C ( clk ), .D ( new_AGEMA_signal_6562 ), .Q ( new_AGEMA_signal_6563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C ( clk ), .D ( new_AGEMA_signal_6566 ), .Q ( new_AGEMA_signal_6567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C ( clk ), .D ( new_AGEMA_signal_6570 ), .Q ( new_AGEMA_signal_6571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C ( clk ), .D ( new_AGEMA_signal_6574 ), .Q ( new_AGEMA_signal_6575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C ( clk ), .D ( new_AGEMA_signal_6578 ), .Q ( new_AGEMA_signal_6579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C ( clk ), .D ( new_AGEMA_signal_6582 ), .Q ( new_AGEMA_signal_6583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C ( clk ), .D ( new_AGEMA_signal_6586 ), .Q ( new_AGEMA_signal_6587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C ( clk ), .D ( new_AGEMA_signal_6590 ), .Q ( new_AGEMA_signal_6591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C ( clk ), .D ( new_AGEMA_signal_6592 ), .Q ( new_AGEMA_signal_6593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C ( clk ), .D ( new_AGEMA_signal_6594 ), .Q ( new_AGEMA_signal_6595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C ( clk ), .D ( new_AGEMA_signal_6596 ), .Q ( new_AGEMA_signal_6597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C ( clk ), .D ( new_AGEMA_signal_6598 ), .Q ( new_AGEMA_signal_6599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C ( clk ), .D ( new_AGEMA_signal_6600 ), .Q ( new_AGEMA_signal_6601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C ( clk ), .D ( new_AGEMA_signal_6602 ), .Q ( new_AGEMA_signal_6603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C ( clk ), .D ( new_AGEMA_signal_6604 ), .Q ( new_AGEMA_signal_6605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C ( clk ), .D ( new_AGEMA_signal_6606 ), .Q ( new_AGEMA_signal_6607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C ( clk ), .D ( new_AGEMA_signal_6608 ), .Q ( new_AGEMA_signal_6609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C ( clk ), .D ( new_AGEMA_signal_6612 ), .Q ( new_AGEMA_signal_6613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C ( clk ), .D ( new_AGEMA_signal_6616 ), .Q ( new_AGEMA_signal_6617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C ( clk ), .D ( new_AGEMA_signal_6620 ), .Q ( new_AGEMA_signal_6621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C ( clk ), .D ( new_AGEMA_signal_6622 ), .Q ( new_AGEMA_signal_6623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C ( clk ), .D ( new_AGEMA_signal_6624 ), .Q ( new_AGEMA_signal_6625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C ( clk ), .D ( new_AGEMA_signal_6626 ), .Q ( new_AGEMA_signal_6627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C ( clk ), .D ( new_AGEMA_signal_6630 ), .Q ( new_AGEMA_signal_6631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2146 ( .C ( clk ), .D ( new_AGEMA_signal_6634 ), .Q ( new_AGEMA_signal_6635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2150 ( .C ( clk ), .D ( new_AGEMA_signal_6638 ), .Q ( new_AGEMA_signal_6639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2156 ( .C ( clk ), .D ( new_AGEMA_signal_6644 ), .Q ( new_AGEMA_signal_6645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2162 ( .C ( clk ), .D ( new_AGEMA_signal_6650 ), .Q ( new_AGEMA_signal_6651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2168 ( .C ( clk ), .D ( new_AGEMA_signal_6656 ), .Q ( new_AGEMA_signal_6657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2172 ( .C ( clk ), .D ( new_AGEMA_signal_6660 ), .Q ( new_AGEMA_signal_6661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2176 ( .C ( clk ), .D ( new_AGEMA_signal_6664 ), .Q ( new_AGEMA_signal_6665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2180 ( .C ( clk ), .D ( new_AGEMA_signal_6668 ), .Q ( new_AGEMA_signal_6669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2184 ( .C ( clk ), .D ( new_AGEMA_signal_6672 ), .Q ( new_AGEMA_signal_6673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2188 ( .C ( clk ), .D ( new_AGEMA_signal_6676 ), .Q ( new_AGEMA_signal_6677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2192 ( .C ( clk ), .D ( new_AGEMA_signal_6680 ), .Q ( new_AGEMA_signal_6681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2194 ( .C ( clk ), .D ( new_AGEMA_signal_6682 ), .Q ( new_AGEMA_signal_6683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2196 ( .C ( clk ), .D ( new_AGEMA_signal_6684 ), .Q ( new_AGEMA_signal_6685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2198 ( .C ( clk ), .D ( new_AGEMA_signal_6686 ), .Q ( new_AGEMA_signal_6687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2200 ( .C ( clk ), .D ( new_AGEMA_signal_6688 ), .Q ( new_AGEMA_signal_6689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2202 ( .C ( clk ), .D ( new_AGEMA_signal_6690 ), .Q ( new_AGEMA_signal_6691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2204 ( .C ( clk ), .D ( new_AGEMA_signal_6692 ), .Q ( new_AGEMA_signal_6693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C ( clk ), .D ( new_AGEMA_signal_6694 ), .Q ( new_AGEMA_signal_6695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C ( clk ), .D ( new_AGEMA_signal_6696 ), .Q ( new_AGEMA_signal_6697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2210 ( .C ( clk ), .D ( new_AGEMA_signal_6698 ), .Q ( new_AGEMA_signal_6699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2212 ( .C ( clk ), .D ( new_AGEMA_signal_6700 ), .Q ( new_AGEMA_signal_6701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2214 ( .C ( clk ), .D ( new_AGEMA_signal_6702 ), .Q ( new_AGEMA_signal_6703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2216 ( .C ( clk ), .D ( new_AGEMA_signal_6704 ), .Q ( new_AGEMA_signal_6705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2220 ( .C ( clk ), .D ( new_AGEMA_signal_6708 ), .Q ( new_AGEMA_signal_6709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2224 ( .C ( clk ), .D ( new_AGEMA_signal_6712 ), .Q ( new_AGEMA_signal_6713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2228 ( .C ( clk ), .D ( new_AGEMA_signal_6716 ), .Q ( new_AGEMA_signal_6717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2234 ( .C ( clk ), .D ( new_AGEMA_signal_6722 ), .Q ( new_AGEMA_signal_6723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2240 ( .C ( clk ), .D ( new_AGEMA_signal_6728 ), .Q ( new_AGEMA_signal_6729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2246 ( .C ( clk ), .D ( new_AGEMA_signal_6734 ), .Q ( new_AGEMA_signal_6735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2250 ( .C ( clk ), .D ( new_AGEMA_signal_6738 ), .Q ( new_AGEMA_signal_6739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C ( clk ), .D ( new_AGEMA_signal_6742 ), .Q ( new_AGEMA_signal_6743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2258 ( .C ( clk ), .D ( new_AGEMA_signal_6746 ), .Q ( new_AGEMA_signal_6747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2260 ( .C ( clk ), .D ( new_AGEMA_signal_6748 ), .Q ( new_AGEMA_signal_6749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2262 ( .C ( clk ), .D ( new_AGEMA_signal_6750 ), .Q ( new_AGEMA_signal_6751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2264 ( .C ( clk ), .D ( new_AGEMA_signal_6752 ), .Q ( new_AGEMA_signal_6753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2266 ( .C ( clk ), .D ( new_AGEMA_signal_6754 ), .Q ( new_AGEMA_signal_6755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2268 ( .C ( clk ), .D ( new_AGEMA_signal_6756 ), .Q ( new_AGEMA_signal_6757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2270 ( .C ( clk ), .D ( new_AGEMA_signal_6758 ), .Q ( new_AGEMA_signal_6759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2272 ( .C ( clk ), .D ( new_AGEMA_signal_6760 ), .Q ( new_AGEMA_signal_6761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2274 ( .C ( clk ), .D ( new_AGEMA_signal_6762 ), .Q ( new_AGEMA_signal_6763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2276 ( .C ( clk ), .D ( new_AGEMA_signal_6764 ), .Q ( new_AGEMA_signal_6765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2280 ( .C ( clk ), .D ( new_AGEMA_signal_6768 ), .Q ( new_AGEMA_signal_6769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2284 ( .C ( clk ), .D ( new_AGEMA_signal_6772 ), .Q ( new_AGEMA_signal_6773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2288 ( .C ( clk ), .D ( new_AGEMA_signal_6776 ), .Q ( new_AGEMA_signal_6777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2290 ( .C ( clk ), .D ( new_AGEMA_signal_6778 ), .Q ( new_AGEMA_signal_6779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2292 ( .C ( clk ), .D ( new_AGEMA_signal_6780 ), .Q ( new_AGEMA_signal_6781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2294 ( .C ( clk ), .D ( new_AGEMA_signal_6782 ), .Q ( new_AGEMA_signal_6783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2296 ( .C ( clk ), .D ( new_AGEMA_signal_6784 ), .Q ( new_AGEMA_signal_6785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2298 ( .C ( clk ), .D ( new_AGEMA_signal_6786 ), .Q ( new_AGEMA_signal_6787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2300 ( .C ( clk ), .D ( new_AGEMA_signal_6788 ), .Q ( new_AGEMA_signal_6789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2304 ( .C ( clk ), .D ( new_AGEMA_signal_6792 ), .Q ( new_AGEMA_signal_6793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2308 ( .C ( clk ), .D ( new_AGEMA_signal_6796 ), .Q ( new_AGEMA_signal_6797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2312 ( .C ( clk ), .D ( new_AGEMA_signal_6800 ), .Q ( new_AGEMA_signal_6801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2316 ( .C ( clk ), .D ( new_AGEMA_signal_6804 ), .Q ( new_AGEMA_signal_6805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2320 ( .C ( clk ), .D ( new_AGEMA_signal_6808 ), .Q ( new_AGEMA_signal_6809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2324 ( .C ( clk ), .D ( new_AGEMA_signal_6812 ), .Q ( new_AGEMA_signal_6813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2328 ( .C ( clk ), .D ( new_AGEMA_signal_6816 ), .Q ( new_AGEMA_signal_6817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2332 ( .C ( clk ), .D ( new_AGEMA_signal_6820 ), .Q ( new_AGEMA_signal_6821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2336 ( .C ( clk ), .D ( new_AGEMA_signal_6824 ), .Q ( new_AGEMA_signal_6825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2340 ( .C ( clk ), .D ( new_AGEMA_signal_6828 ), .Q ( new_AGEMA_signal_6829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2344 ( .C ( clk ), .D ( new_AGEMA_signal_6832 ), .Q ( new_AGEMA_signal_6833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2348 ( .C ( clk ), .D ( new_AGEMA_signal_6836 ), .Q ( new_AGEMA_signal_6837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2352 ( .C ( clk ), .D ( new_AGEMA_signal_6840 ), .Q ( new_AGEMA_signal_6841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2356 ( .C ( clk ), .D ( new_AGEMA_signal_6844 ), .Q ( new_AGEMA_signal_6845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2360 ( .C ( clk ), .D ( new_AGEMA_signal_6848 ), .Q ( new_AGEMA_signal_6849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2362 ( .C ( clk ), .D ( new_AGEMA_signal_6850 ), .Q ( new_AGEMA_signal_6851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2364 ( .C ( clk ), .D ( new_AGEMA_signal_6852 ), .Q ( new_AGEMA_signal_6853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2366 ( .C ( clk ), .D ( new_AGEMA_signal_6854 ), .Q ( new_AGEMA_signal_6855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2368 ( .C ( clk ), .D ( new_AGEMA_signal_6856 ), .Q ( new_AGEMA_signal_6857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2370 ( .C ( clk ), .D ( new_AGEMA_signal_6858 ), .Q ( new_AGEMA_signal_6859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2372 ( .C ( clk ), .D ( new_AGEMA_signal_6860 ), .Q ( new_AGEMA_signal_6861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2374 ( .C ( clk ), .D ( new_AGEMA_signal_6862 ), .Q ( new_AGEMA_signal_6863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2376 ( .C ( clk ), .D ( new_AGEMA_signal_6864 ), .Q ( new_AGEMA_signal_6865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2378 ( .C ( clk ), .D ( new_AGEMA_signal_6866 ), .Q ( new_AGEMA_signal_6867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2380 ( .C ( clk ), .D ( new_AGEMA_signal_6868 ), .Q ( new_AGEMA_signal_6869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2382 ( .C ( clk ), .D ( new_AGEMA_signal_6870 ), .Q ( new_AGEMA_signal_6871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2384 ( .C ( clk ), .D ( new_AGEMA_signal_6872 ), .Q ( new_AGEMA_signal_6873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2388 ( .C ( clk ), .D ( new_AGEMA_signal_6876 ), .Q ( new_AGEMA_signal_6877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2392 ( .C ( clk ), .D ( new_AGEMA_signal_6880 ), .Q ( new_AGEMA_signal_6881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2396 ( .C ( clk ), .D ( new_AGEMA_signal_6884 ), .Q ( new_AGEMA_signal_6885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2400 ( .C ( clk ), .D ( new_AGEMA_signal_6888 ), .Q ( new_AGEMA_signal_6889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2404 ( .C ( clk ), .D ( new_AGEMA_signal_6892 ), .Q ( new_AGEMA_signal_6893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2408 ( .C ( clk ), .D ( new_AGEMA_signal_6896 ), .Q ( new_AGEMA_signal_6897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2410 ( .C ( clk ), .D ( new_AGEMA_signal_6898 ), .Q ( new_AGEMA_signal_6899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2412 ( .C ( clk ), .D ( new_AGEMA_signal_6900 ), .Q ( new_AGEMA_signal_6901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2414 ( .C ( clk ), .D ( new_AGEMA_signal_6902 ), .Q ( new_AGEMA_signal_6903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2416 ( .C ( clk ), .D ( new_AGEMA_signal_6904 ), .Q ( new_AGEMA_signal_6905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2418 ( .C ( clk ), .D ( new_AGEMA_signal_6906 ), .Q ( new_AGEMA_signal_6907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2420 ( .C ( clk ), .D ( new_AGEMA_signal_6908 ), .Q ( new_AGEMA_signal_6909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2422 ( .C ( clk ), .D ( new_AGEMA_signal_6910 ), .Q ( new_AGEMA_signal_6911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2424 ( .C ( clk ), .D ( new_AGEMA_signal_6912 ), .Q ( new_AGEMA_signal_6913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2426 ( .C ( clk ), .D ( new_AGEMA_signal_6914 ), .Q ( new_AGEMA_signal_6915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2428 ( .C ( clk ), .D ( new_AGEMA_signal_6916 ), .Q ( new_AGEMA_signal_6917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2430 ( .C ( clk ), .D ( new_AGEMA_signal_6918 ), .Q ( new_AGEMA_signal_6919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2432 ( .C ( clk ), .D ( new_AGEMA_signal_6920 ), .Q ( new_AGEMA_signal_6921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2434 ( .C ( clk ), .D ( new_AGEMA_signal_6922 ), .Q ( new_AGEMA_signal_6923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2436 ( .C ( clk ), .D ( new_AGEMA_signal_6924 ), .Q ( new_AGEMA_signal_6925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2438 ( .C ( clk ), .D ( new_AGEMA_signal_6926 ), .Q ( new_AGEMA_signal_6927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2440 ( .C ( clk ), .D ( new_AGEMA_signal_6928 ), .Q ( new_AGEMA_signal_6929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2442 ( .C ( clk ), .D ( new_AGEMA_signal_6930 ), .Q ( new_AGEMA_signal_6931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2444 ( .C ( clk ), .D ( new_AGEMA_signal_6932 ), .Q ( new_AGEMA_signal_6933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2446 ( .C ( clk ), .D ( new_AGEMA_signal_6934 ), .Q ( new_AGEMA_signal_6935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2448 ( .C ( clk ), .D ( new_AGEMA_signal_6936 ), .Q ( new_AGEMA_signal_6937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2450 ( .C ( clk ), .D ( new_AGEMA_signal_6938 ), .Q ( new_AGEMA_signal_6939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2452 ( .C ( clk ), .D ( new_AGEMA_signal_6940 ), .Q ( new_AGEMA_signal_6941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2454 ( .C ( clk ), .D ( new_AGEMA_signal_6942 ), .Q ( new_AGEMA_signal_6943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2456 ( .C ( clk ), .D ( new_AGEMA_signal_6944 ), .Q ( new_AGEMA_signal_6945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2458 ( .C ( clk ), .D ( new_AGEMA_signal_6946 ), .Q ( new_AGEMA_signal_6947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2460 ( .C ( clk ), .D ( new_AGEMA_signal_6948 ), .Q ( new_AGEMA_signal_6949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2462 ( .C ( clk ), .D ( new_AGEMA_signal_6950 ), .Q ( new_AGEMA_signal_6951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2466 ( .C ( clk ), .D ( new_AGEMA_signal_6954 ), .Q ( new_AGEMA_signal_6955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2470 ( .C ( clk ), .D ( new_AGEMA_signal_6958 ), .Q ( new_AGEMA_signal_6959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2474 ( .C ( clk ), .D ( new_AGEMA_signal_6962 ), .Q ( new_AGEMA_signal_6963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2476 ( .C ( clk ), .D ( new_AGEMA_signal_6964 ), .Q ( new_AGEMA_signal_6965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2478 ( .C ( clk ), .D ( new_AGEMA_signal_6966 ), .Q ( new_AGEMA_signal_6967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2480 ( .C ( clk ), .D ( new_AGEMA_signal_6968 ), .Q ( new_AGEMA_signal_6969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2482 ( .C ( clk ), .D ( new_AGEMA_signal_6970 ), .Q ( new_AGEMA_signal_6971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2484 ( .C ( clk ), .D ( new_AGEMA_signal_6972 ), .Q ( new_AGEMA_signal_6973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2486 ( .C ( clk ), .D ( new_AGEMA_signal_6974 ), .Q ( new_AGEMA_signal_6975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2488 ( .C ( clk ), .D ( new_AGEMA_signal_6976 ), .Q ( new_AGEMA_signal_6977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2490 ( .C ( clk ), .D ( new_AGEMA_signal_6978 ), .Q ( new_AGEMA_signal_6979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2492 ( .C ( clk ), .D ( new_AGEMA_signal_6980 ), .Q ( new_AGEMA_signal_6981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2494 ( .C ( clk ), .D ( new_AGEMA_signal_6982 ), .Q ( new_AGEMA_signal_6983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2496 ( .C ( clk ), .D ( new_AGEMA_signal_6984 ), .Q ( new_AGEMA_signal_6985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2498 ( .C ( clk ), .D ( new_AGEMA_signal_6986 ), .Q ( new_AGEMA_signal_6987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2500 ( .C ( clk ), .D ( new_AGEMA_signal_6988 ), .Q ( new_AGEMA_signal_6989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2502 ( .C ( clk ), .D ( new_AGEMA_signal_6990 ), .Q ( new_AGEMA_signal_6991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2504 ( .C ( clk ), .D ( new_AGEMA_signal_6992 ), .Q ( new_AGEMA_signal_6993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2508 ( .C ( clk ), .D ( new_AGEMA_signal_6996 ), .Q ( new_AGEMA_signal_6997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2512 ( .C ( clk ), .D ( new_AGEMA_signal_7000 ), .Q ( new_AGEMA_signal_7001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2516 ( .C ( clk ), .D ( new_AGEMA_signal_7004 ), .Q ( new_AGEMA_signal_7005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2520 ( .C ( clk ), .D ( new_AGEMA_signal_7008 ), .Q ( new_AGEMA_signal_7009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2524 ( .C ( clk ), .D ( new_AGEMA_signal_7012 ), .Q ( new_AGEMA_signal_7013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2528 ( .C ( clk ), .D ( new_AGEMA_signal_7016 ), .Q ( new_AGEMA_signal_7017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2532 ( .C ( clk ), .D ( new_AGEMA_signal_7020 ), .Q ( new_AGEMA_signal_7021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2536 ( .C ( clk ), .D ( new_AGEMA_signal_7024 ), .Q ( new_AGEMA_signal_7025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2540 ( .C ( clk ), .D ( new_AGEMA_signal_7028 ), .Q ( new_AGEMA_signal_7029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2544 ( .C ( clk ), .D ( new_AGEMA_signal_7032 ), .Q ( new_AGEMA_signal_7033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2548 ( .C ( clk ), .D ( new_AGEMA_signal_7036 ), .Q ( new_AGEMA_signal_7037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2552 ( .C ( clk ), .D ( new_AGEMA_signal_7040 ), .Q ( new_AGEMA_signal_7041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2554 ( .C ( clk ), .D ( new_AGEMA_signal_7042 ), .Q ( new_AGEMA_signal_7043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2558 ( .C ( clk ), .D ( new_AGEMA_signal_7046 ), .Q ( new_AGEMA_signal_7047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2562 ( .C ( clk ), .D ( new_AGEMA_signal_7050 ), .Q ( new_AGEMA_signal_7051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2566 ( .C ( clk ), .D ( new_AGEMA_signal_7054 ), .Q ( new_AGEMA_signal_7055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2570 ( .C ( clk ), .D ( new_AGEMA_signal_7058 ), .Q ( new_AGEMA_signal_7059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2574 ( .C ( clk ), .D ( new_AGEMA_signal_7062 ), .Q ( new_AGEMA_signal_7063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2582 ( .C ( clk ), .D ( new_AGEMA_signal_7070 ), .Q ( new_AGEMA_signal_7071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2590 ( .C ( clk ), .D ( new_AGEMA_signal_7078 ), .Q ( new_AGEMA_signal_7079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2598 ( .C ( clk ), .D ( new_AGEMA_signal_7086 ), .Q ( new_AGEMA_signal_7087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2612 ( .C ( clk ), .D ( new_AGEMA_signal_7100 ), .Q ( new_AGEMA_signal_7101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2620 ( .C ( clk ), .D ( new_AGEMA_signal_7108 ), .Q ( new_AGEMA_signal_7109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2628 ( .C ( clk ), .D ( new_AGEMA_signal_7116 ), .Q ( new_AGEMA_signal_7117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2634 ( .C ( clk ), .D ( new_AGEMA_signal_7122 ), .Q ( new_AGEMA_signal_7123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2640 ( .C ( clk ), .D ( new_AGEMA_signal_7128 ), .Q ( new_AGEMA_signal_7129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2646 ( .C ( clk ), .D ( new_AGEMA_signal_7134 ), .Q ( new_AGEMA_signal_7135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2650 ( .C ( clk ), .D ( new_AGEMA_signal_7138 ), .Q ( new_AGEMA_signal_7139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2654 ( .C ( clk ), .D ( new_AGEMA_signal_7142 ), .Q ( new_AGEMA_signal_7143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2658 ( .C ( clk ), .D ( new_AGEMA_signal_7146 ), .Q ( new_AGEMA_signal_7147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2664 ( .C ( clk ), .D ( new_AGEMA_signal_7152 ), .Q ( new_AGEMA_signal_7153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2670 ( .C ( clk ), .D ( new_AGEMA_signal_7158 ), .Q ( new_AGEMA_signal_7159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2676 ( .C ( clk ), .D ( new_AGEMA_signal_7164 ), .Q ( new_AGEMA_signal_7165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2688 ( .C ( clk ), .D ( new_AGEMA_signal_7176 ), .Q ( new_AGEMA_signal_7177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2694 ( .C ( clk ), .D ( new_AGEMA_signal_7182 ), .Q ( new_AGEMA_signal_7183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2700 ( .C ( clk ), .D ( new_AGEMA_signal_7188 ), .Q ( new_AGEMA_signal_7189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2706 ( .C ( clk ), .D ( new_AGEMA_signal_7194 ), .Q ( new_AGEMA_signal_7195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2712 ( .C ( clk ), .D ( new_AGEMA_signal_7200 ), .Q ( new_AGEMA_signal_7201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2718 ( .C ( clk ), .D ( new_AGEMA_signal_7206 ), .Q ( new_AGEMA_signal_7207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2728 ( .C ( clk ), .D ( new_AGEMA_signal_7216 ), .Q ( new_AGEMA_signal_7217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2732 ( .C ( clk ), .D ( new_AGEMA_signal_7220 ), .Q ( new_AGEMA_signal_7221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2736 ( .C ( clk ), .D ( new_AGEMA_signal_7224 ), .Q ( new_AGEMA_signal_7225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2742 ( .C ( clk ), .D ( new_AGEMA_signal_7230 ), .Q ( new_AGEMA_signal_7231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2748 ( .C ( clk ), .D ( new_AGEMA_signal_7236 ), .Q ( new_AGEMA_signal_7237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2754 ( .C ( clk ), .D ( new_AGEMA_signal_7242 ), .Q ( new_AGEMA_signal_7243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2760 ( .C ( clk ), .D ( new_AGEMA_signal_7248 ), .Q ( new_AGEMA_signal_7249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2766 ( .C ( clk ), .D ( new_AGEMA_signal_7254 ), .Q ( new_AGEMA_signal_7255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2772 ( .C ( clk ), .D ( new_AGEMA_signal_7260 ), .Q ( new_AGEMA_signal_7261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2784 ( .C ( clk ), .D ( new_AGEMA_signal_7272 ), .Q ( new_AGEMA_signal_7273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2790 ( .C ( clk ), .D ( new_AGEMA_signal_7278 ), .Q ( new_AGEMA_signal_7279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2796 ( .C ( clk ), .D ( new_AGEMA_signal_7284 ), .Q ( new_AGEMA_signal_7285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2806 ( .C ( clk ), .D ( new_AGEMA_signal_7294 ), .Q ( new_AGEMA_signal_7295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2810 ( .C ( clk ), .D ( new_AGEMA_signal_7298 ), .Q ( new_AGEMA_signal_7299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2814 ( .C ( clk ), .D ( new_AGEMA_signal_7302 ), .Q ( new_AGEMA_signal_7303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2818 ( .C ( clk ), .D ( new_AGEMA_signal_7306 ), .Q ( new_AGEMA_signal_7307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2822 ( .C ( clk ), .D ( new_AGEMA_signal_7310 ), .Q ( new_AGEMA_signal_7311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2826 ( .C ( clk ), .D ( new_AGEMA_signal_7314 ), .Q ( new_AGEMA_signal_7315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2840 ( .C ( clk ), .D ( new_AGEMA_signal_7328 ), .Q ( new_AGEMA_signal_7329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2848 ( .C ( clk ), .D ( new_AGEMA_signal_7336 ), .Q ( new_AGEMA_signal_7337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2856 ( .C ( clk ), .D ( new_AGEMA_signal_7344 ), .Q ( new_AGEMA_signal_7345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2862 ( .C ( clk ), .D ( new_AGEMA_signal_7350 ), .Q ( new_AGEMA_signal_7351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2868 ( .C ( clk ), .D ( new_AGEMA_signal_7356 ), .Q ( new_AGEMA_signal_7357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2874 ( .C ( clk ), .D ( new_AGEMA_signal_7362 ), .Q ( new_AGEMA_signal_7363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2878 ( .C ( clk ), .D ( new_AGEMA_signal_7366 ), .Q ( new_AGEMA_signal_7367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2882 ( .C ( clk ), .D ( new_AGEMA_signal_7370 ), .Q ( new_AGEMA_signal_7371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2886 ( .C ( clk ), .D ( new_AGEMA_signal_7374 ), .Q ( new_AGEMA_signal_7375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2890 ( .C ( clk ), .D ( new_AGEMA_signal_7378 ), .Q ( new_AGEMA_signal_7379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2894 ( .C ( clk ), .D ( new_AGEMA_signal_7382 ), .Q ( new_AGEMA_signal_7383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2898 ( .C ( clk ), .D ( new_AGEMA_signal_7386 ), .Q ( new_AGEMA_signal_7387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2914 ( .C ( clk ), .D ( new_AGEMA_signal_7402 ), .Q ( new_AGEMA_signal_7403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2918 ( .C ( clk ), .D ( new_AGEMA_signal_7406 ), .Q ( new_AGEMA_signal_7407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2922 ( .C ( clk ), .D ( new_AGEMA_signal_7410 ), .Q ( new_AGEMA_signal_7411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2926 ( .C ( clk ), .D ( new_AGEMA_signal_7414 ), .Q ( new_AGEMA_signal_7415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2930 ( .C ( clk ), .D ( new_AGEMA_signal_7418 ), .Q ( new_AGEMA_signal_7419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2934 ( .C ( clk ), .D ( new_AGEMA_signal_7422 ), .Q ( new_AGEMA_signal_7423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2946 ( .C ( clk ), .D ( new_AGEMA_signal_7434 ), .Q ( new_AGEMA_signal_7435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2952 ( .C ( clk ), .D ( new_AGEMA_signal_7440 ), .Q ( new_AGEMA_signal_7441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2958 ( .C ( clk ), .D ( new_AGEMA_signal_7446 ), .Q ( new_AGEMA_signal_7447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2962 ( .C ( clk ), .D ( new_AGEMA_signal_7450 ), .Q ( new_AGEMA_signal_7451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2966 ( .C ( clk ), .D ( new_AGEMA_signal_7454 ), .Q ( new_AGEMA_signal_7455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2970 ( .C ( clk ), .D ( new_AGEMA_signal_7458 ), .Q ( new_AGEMA_signal_7459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2980 ( .C ( clk ), .D ( new_AGEMA_signal_7468 ), .Q ( new_AGEMA_signal_7469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2984 ( .C ( clk ), .D ( new_AGEMA_signal_7472 ), .Q ( new_AGEMA_signal_7473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2988 ( .C ( clk ), .D ( new_AGEMA_signal_7476 ), .Q ( new_AGEMA_signal_7477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2992 ( .C ( clk ), .D ( new_AGEMA_signal_7480 ), .Q ( new_AGEMA_signal_7481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2996 ( .C ( clk ), .D ( new_AGEMA_signal_7484 ), .Q ( new_AGEMA_signal_7485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3000 ( .C ( clk ), .D ( new_AGEMA_signal_7488 ), .Q ( new_AGEMA_signal_7489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3004 ( .C ( clk ), .D ( new_AGEMA_signal_7492 ), .Q ( new_AGEMA_signal_7493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3008 ( .C ( clk ), .D ( new_AGEMA_signal_7496 ), .Q ( new_AGEMA_signal_7497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3012 ( .C ( clk ), .D ( new_AGEMA_signal_7500 ), .Q ( new_AGEMA_signal_7501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3022 ( .C ( clk ), .D ( new_AGEMA_signal_7510 ), .Q ( new_AGEMA_signal_7511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3026 ( .C ( clk ), .D ( new_AGEMA_signal_7514 ), .Q ( new_AGEMA_signal_7515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3030 ( .C ( clk ), .D ( new_AGEMA_signal_7518 ), .Q ( new_AGEMA_signal_7519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3042 ( .C ( clk ), .D ( new_AGEMA_signal_7530 ), .Q ( new_AGEMA_signal_7531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3048 ( .C ( clk ), .D ( new_AGEMA_signal_7536 ), .Q ( new_AGEMA_signal_7537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3054 ( .C ( clk ), .D ( new_AGEMA_signal_7542 ), .Q ( new_AGEMA_signal_7543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3060 ( .C ( clk ), .D ( new_AGEMA_signal_7548 ), .Q ( new_AGEMA_signal_7549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3066 ( .C ( clk ), .D ( new_AGEMA_signal_7554 ), .Q ( new_AGEMA_signal_7555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3072 ( .C ( clk ), .D ( new_AGEMA_signal_7560 ), .Q ( new_AGEMA_signal_7561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3076 ( .C ( clk ), .D ( new_AGEMA_signal_7564 ), .Q ( new_AGEMA_signal_7565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3080 ( .C ( clk ), .D ( new_AGEMA_signal_7568 ), .Q ( new_AGEMA_signal_7569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3084 ( .C ( clk ), .D ( new_AGEMA_signal_7572 ), .Q ( new_AGEMA_signal_7573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3098 ( .C ( clk ), .D ( new_AGEMA_signal_7586 ), .Q ( new_AGEMA_signal_7587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3106 ( .C ( clk ), .D ( new_AGEMA_signal_7594 ), .Q ( new_AGEMA_signal_7595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3114 ( .C ( clk ), .D ( new_AGEMA_signal_7602 ), .Q ( new_AGEMA_signal_7603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3124 ( .C ( clk ), .D ( new_AGEMA_signal_7612 ), .Q ( new_AGEMA_signal_7613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3128 ( .C ( clk ), .D ( new_AGEMA_signal_7616 ), .Q ( new_AGEMA_signal_7617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3132 ( .C ( clk ), .D ( new_AGEMA_signal_7620 ), .Q ( new_AGEMA_signal_7621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3136 ( .C ( clk ), .D ( new_AGEMA_signal_7624 ), .Q ( new_AGEMA_signal_7625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3140 ( .C ( clk ), .D ( new_AGEMA_signal_7628 ), .Q ( new_AGEMA_signal_7629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3144 ( .C ( clk ), .D ( new_AGEMA_signal_7632 ), .Q ( new_AGEMA_signal_7633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3148 ( .C ( clk ), .D ( new_AGEMA_signal_7636 ), .Q ( new_AGEMA_signal_7637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3152 ( .C ( clk ), .D ( new_AGEMA_signal_7640 ), .Q ( new_AGEMA_signal_7641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3156 ( .C ( clk ), .D ( new_AGEMA_signal_7644 ), .Q ( new_AGEMA_signal_7645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3160 ( .C ( clk ), .D ( new_AGEMA_signal_7648 ), .Q ( new_AGEMA_signal_7649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3164 ( .C ( clk ), .D ( new_AGEMA_signal_7652 ), .Q ( new_AGEMA_signal_7653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3168 ( .C ( clk ), .D ( new_AGEMA_signal_7656 ), .Q ( new_AGEMA_signal_7657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3172 ( .C ( clk ), .D ( new_AGEMA_signal_7660 ), .Q ( new_AGEMA_signal_7661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3176 ( .C ( clk ), .D ( new_AGEMA_signal_7664 ), .Q ( new_AGEMA_signal_7665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3180 ( .C ( clk ), .D ( new_AGEMA_signal_7668 ), .Q ( new_AGEMA_signal_7669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3188 ( .C ( clk ), .D ( new_AGEMA_signal_7676 ), .Q ( new_AGEMA_signal_7677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3196 ( .C ( clk ), .D ( new_AGEMA_signal_7684 ), .Q ( new_AGEMA_signal_7685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3204 ( .C ( clk ), .D ( new_AGEMA_signal_7692 ), .Q ( new_AGEMA_signal_7693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3214 ( .C ( clk ), .D ( new_AGEMA_signal_7702 ), .Q ( new_AGEMA_signal_7703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3218 ( .C ( clk ), .D ( new_AGEMA_signal_7706 ), .Q ( new_AGEMA_signal_7707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3222 ( .C ( clk ), .D ( new_AGEMA_signal_7710 ), .Q ( new_AGEMA_signal_7711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3234 ( .C ( clk ), .D ( new_AGEMA_signal_7722 ), .Q ( new_AGEMA_signal_7723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3240 ( .C ( clk ), .D ( new_AGEMA_signal_7728 ), .Q ( new_AGEMA_signal_7729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3246 ( .C ( clk ), .D ( new_AGEMA_signal_7734 ), .Q ( new_AGEMA_signal_7735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3258 ( .C ( clk ), .D ( new_AGEMA_signal_7746 ), .Q ( new_AGEMA_signal_7747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3266 ( .C ( clk ), .D ( new_AGEMA_signal_7754 ), .Q ( new_AGEMA_signal_7755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3274 ( .C ( clk ), .D ( new_AGEMA_signal_7762 ), .Q ( new_AGEMA_signal_7763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3300 ( .C ( clk ), .D ( new_AGEMA_signal_7788 ), .Q ( new_AGEMA_signal_7789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3308 ( .C ( clk ), .D ( new_AGEMA_signal_7796 ), .Q ( new_AGEMA_signal_7797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3316 ( .C ( clk ), .D ( new_AGEMA_signal_7804 ), .Q ( new_AGEMA_signal_7805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3328 ( .C ( clk ), .D ( new_AGEMA_signal_7816 ), .Q ( new_AGEMA_signal_7817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3334 ( .C ( clk ), .D ( new_AGEMA_signal_7822 ), .Q ( new_AGEMA_signal_7823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3340 ( .C ( clk ), .D ( new_AGEMA_signal_7828 ), .Q ( new_AGEMA_signal_7829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3360 ( .C ( clk ), .D ( new_AGEMA_signal_7848 ), .Q ( new_AGEMA_signal_7849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3368 ( .C ( clk ), .D ( new_AGEMA_signal_7856 ), .Q ( new_AGEMA_signal_7857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3376 ( .C ( clk ), .D ( new_AGEMA_signal_7864 ), .Q ( new_AGEMA_signal_7865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3394 ( .C ( clk ), .D ( new_AGEMA_signal_7882 ), .Q ( new_AGEMA_signal_7883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3400 ( .C ( clk ), .D ( new_AGEMA_signal_7888 ), .Q ( new_AGEMA_signal_7889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3406 ( .C ( clk ), .D ( new_AGEMA_signal_7894 ), .Q ( new_AGEMA_signal_7895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3412 ( .C ( clk ), .D ( new_AGEMA_signal_7900 ), .Q ( new_AGEMA_signal_7901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3418 ( .C ( clk ), .D ( new_AGEMA_signal_7906 ), .Q ( new_AGEMA_signal_7907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3424 ( .C ( clk ), .D ( new_AGEMA_signal_7912 ), .Q ( new_AGEMA_signal_7913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3430 ( .C ( clk ), .D ( new_AGEMA_signal_7918 ), .Q ( new_AGEMA_signal_7919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3436 ( .C ( clk ), .D ( new_AGEMA_signal_7924 ), .Q ( new_AGEMA_signal_7925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3442 ( .C ( clk ), .D ( new_AGEMA_signal_7930 ), .Q ( new_AGEMA_signal_7931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3448 ( .C ( clk ), .D ( new_AGEMA_signal_7936 ), .Q ( new_AGEMA_signal_7937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3454 ( .C ( clk ), .D ( new_AGEMA_signal_7942 ), .Q ( new_AGEMA_signal_7943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3460 ( .C ( clk ), .D ( new_AGEMA_signal_7948 ), .Q ( new_AGEMA_signal_7949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3466 ( .C ( clk ), .D ( new_AGEMA_signal_7954 ), .Q ( new_AGEMA_signal_7955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3472 ( .C ( clk ), .D ( new_AGEMA_signal_7960 ), .Q ( new_AGEMA_signal_7961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3478 ( .C ( clk ), .D ( new_AGEMA_signal_7966 ), .Q ( new_AGEMA_signal_7967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3498 ( .C ( clk ), .D ( new_AGEMA_signal_7986 ), .Q ( new_AGEMA_signal_7987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3506 ( .C ( clk ), .D ( new_AGEMA_signal_7994 ), .Q ( new_AGEMA_signal_7995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3514 ( .C ( clk ), .D ( new_AGEMA_signal_8002 ), .Q ( new_AGEMA_signal_8003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3532 ( .C ( clk ), .D ( new_AGEMA_signal_8020 ), .Q ( new_AGEMA_signal_8021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3538 ( .C ( clk ), .D ( new_AGEMA_signal_8026 ), .Q ( new_AGEMA_signal_8027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3544 ( .C ( clk ), .D ( new_AGEMA_signal_8032 ), .Q ( new_AGEMA_signal_8033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3552 ( .C ( clk ), .D ( new_AGEMA_signal_8040 ), .Q ( new_AGEMA_signal_8041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3560 ( .C ( clk ), .D ( new_AGEMA_signal_8048 ), .Q ( new_AGEMA_signal_8049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3568 ( .C ( clk ), .D ( new_AGEMA_signal_8056 ), .Q ( new_AGEMA_signal_8057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3580 ( .C ( clk ), .D ( new_AGEMA_signal_8068 ), .Q ( new_AGEMA_signal_8069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3586 ( .C ( clk ), .D ( new_AGEMA_signal_8074 ), .Q ( new_AGEMA_signal_8075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3592 ( .C ( clk ), .D ( new_AGEMA_signal_8080 ), .Q ( new_AGEMA_signal_8081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3610 ( .C ( clk ), .D ( new_AGEMA_signal_8098 ), .Q ( new_AGEMA_signal_8099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3616 ( .C ( clk ), .D ( new_AGEMA_signal_8104 ), .Q ( new_AGEMA_signal_8105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3622 ( .C ( clk ), .D ( new_AGEMA_signal_8110 ), .Q ( new_AGEMA_signal_8111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3628 ( .C ( clk ), .D ( new_AGEMA_signal_8116 ), .Q ( new_AGEMA_signal_8117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3634 ( .C ( clk ), .D ( new_AGEMA_signal_8122 ), .Q ( new_AGEMA_signal_8123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3640 ( .C ( clk ), .D ( new_AGEMA_signal_8128 ), .Q ( new_AGEMA_signal_8129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3648 ( .C ( clk ), .D ( new_AGEMA_signal_8136 ), .Q ( new_AGEMA_signal_8137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3656 ( .C ( clk ), .D ( new_AGEMA_signal_8144 ), .Q ( new_AGEMA_signal_8145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3664 ( .C ( clk ), .D ( new_AGEMA_signal_8152 ), .Q ( new_AGEMA_signal_8153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3672 ( .C ( clk ), .D ( new_AGEMA_signal_8160 ), .Q ( new_AGEMA_signal_8161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3680 ( .C ( clk ), .D ( new_AGEMA_signal_8168 ), .Q ( new_AGEMA_signal_8169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3688 ( .C ( clk ), .D ( new_AGEMA_signal_8176 ), .Q ( new_AGEMA_signal_8177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3694 ( .C ( clk ), .D ( new_AGEMA_signal_8182 ), .Q ( new_AGEMA_signal_8183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3700 ( .C ( clk ), .D ( new_AGEMA_signal_8188 ), .Q ( new_AGEMA_signal_8189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3706 ( .C ( clk ), .D ( new_AGEMA_signal_8194 ), .Q ( new_AGEMA_signal_8195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3712 ( .C ( clk ), .D ( new_AGEMA_signal_8200 ), .Q ( new_AGEMA_signal_8201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3718 ( .C ( clk ), .D ( new_AGEMA_signal_8206 ), .Q ( new_AGEMA_signal_8207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3724 ( .C ( clk ), .D ( new_AGEMA_signal_8212 ), .Q ( new_AGEMA_signal_8213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3814 ( .C ( clk ), .D ( new_AGEMA_signal_8302 ), .Q ( new_AGEMA_signal_8303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3822 ( .C ( clk ), .D ( new_AGEMA_signal_8310 ), .Q ( new_AGEMA_signal_8311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3830 ( .C ( clk ), .D ( new_AGEMA_signal_8318 ), .Q ( new_AGEMA_signal_8319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3838 ( .C ( clk ), .D ( new_AGEMA_signal_8326 ), .Q ( new_AGEMA_signal_8327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3846 ( .C ( clk ), .D ( new_AGEMA_signal_8334 ), .Q ( new_AGEMA_signal_8335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3854 ( .C ( clk ), .D ( new_AGEMA_signal_8342 ), .Q ( new_AGEMA_signal_8343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3862 ( .C ( clk ), .D ( new_AGEMA_signal_8350 ), .Q ( new_AGEMA_signal_8351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3870 ( .C ( clk ), .D ( new_AGEMA_signal_8358 ), .Q ( new_AGEMA_signal_8359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3878 ( .C ( clk ), .D ( new_AGEMA_signal_8366 ), .Q ( new_AGEMA_signal_8367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3886 ( .C ( clk ), .D ( new_AGEMA_signal_8374 ), .Q ( new_AGEMA_signal_8375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3894 ( .C ( clk ), .D ( new_AGEMA_signal_8382 ), .Q ( new_AGEMA_signal_8383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3902 ( .C ( clk ), .D ( new_AGEMA_signal_8390 ), .Q ( new_AGEMA_signal_8391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3930 ( .C ( clk ), .D ( new_AGEMA_signal_8418 ), .Q ( new_AGEMA_signal_8419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3940 ( .C ( clk ), .D ( new_AGEMA_signal_8428 ), .Q ( new_AGEMA_signal_8429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3950 ( .C ( clk ), .D ( new_AGEMA_signal_8438 ), .Q ( new_AGEMA_signal_8439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3958 ( .C ( clk ), .D ( new_AGEMA_signal_8446 ), .Q ( new_AGEMA_signal_8447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3966 ( .C ( clk ), .D ( new_AGEMA_signal_8454 ), .Q ( new_AGEMA_signal_8455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3974 ( .C ( clk ), .D ( new_AGEMA_signal_8462 ), .Q ( new_AGEMA_signal_8463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3982 ( .C ( clk ), .D ( new_AGEMA_signal_8470 ), .Q ( new_AGEMA_signal_8471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3990 ( .C ( clk ), .D ( new_AGEMA_signal_8478 ), .Q ( new_AGEMA_signal_8479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3998 ( .C ( clk ), .D ( new_AGEMA_signal_8486 ), .Q ( new_AGEMA_signal_8487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4006 ( .C ( clk ), .D ( new_AGEMA_signal_8494 ), .Q ( new_AGEMA_signal_8495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4014 ( .C ( clk ), .D ( new_AGEMA_signal_8502 ), .Q ( new_AGEMA_signal_8503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4022 ( .C ( clk ), .D ( new_AGEMA_signal_8510 ), .Q ( new_AGEMA_signal_8511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4080 ( .C ( clk ), .D ( new_AGEMA_signal_8568 ), .Q ( new_AGEMA_signal_8569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4090 ( .C ( clk ), .D ( new_AGEMA_signal_8578 ), .Q ( new_AGEMA_signal_8579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4100 ( .C ( clk ), .D ( new_AGEMA_signal_8588 ), .Q ( new_AGEMA_signal_8589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4108 ( .C ( clk ), .D ( new_AGEMA_signal_8596 ), .Q ( new_AGEMA_signal_8597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4116 ( .C ( clk ), .D ( new_AGEMA_signal_8604 ), .Q ( new_AGEMA_signal_8605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4124 ( .C ( clk ), .D ( new_AGEMA_signal_8612 ), .Q ( new_AGEMA_signal_8613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4150 ( .C ( clk ), .D ( new_AGEMA_signal_8638 ), .Q ( new_AGEMA_signal_8639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4158 ( .C ( clk ), .D ( new_AGEMA_signal_8646 ), .Q ( new_AGEMA_signal_8647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4166 ( .C ( clk ), .D ( new_AGEMA_signal_8654 ), .Q ( new_AGEMA_signal_8655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4174 ( .C ( clk ), .D ( new_AGEMA_signal_8662 ), .Q ( new_AGEMA_signal_8663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4182 ( .C ( clk ), .D ( new_AGEMA_signal_8670 ), .Q ( new_AGEMA_signal_8671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4190 ( .C ( clk ), .D ( new_AGEMA_signal_8678 ), .Q ( new_AGEMA_signal_8679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4228 ( .C ( clk ), .D ( new_AGEMA_signal_8716 ), .Q ( new_AGEMA_signal_8717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4236 ( .C ( clk ), .D ( new_AGEMA_signal_8724 ), .Q ( new_AGEMA_signal_8725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4244 ( .C ( clk ), .D ( new_AGEMA_signal_8732 ), .Q ( new_AGEMA_signal_8733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4426 ( .C ( clk ), .D ( new_AGEMA_signal_8914 ), .Q ( new_AGEMA_signal_8915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4436 ( .C ( clk ), .D ( new_AGEMA_signal_8924 ), .Q ( new_AGEMA_signal_8925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4446 ( .C ( clk ), .D ( new_AGEMA_signal_8934 ), .Q ( new_AGEMA_signal_8935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5014 ( .C ( clk ), .D ( new_AGEMA_signal_9502 ), .Q ( new_AGEMA_signal_9503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5028 ( .C ( clk ), .D ( new_AGEMA_signal_9516 ), .Q ( new_AGEMA_signal_9517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5042 ( .C ( clk ), .D ( new_AGEMA_signal_9530 ), .Q ( new_AGEMA_signal_9531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5080 ( .C ( clk ), .D ( new_AGEMA_signal_9568 ), .Q ( new_AGEMA_signal_9569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5094 ( .C ( clk ), .D ( new_AGEMA_signal_9582 ), .Q ( new_AGEMA_signal_9583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5108 ( .C ( clk ), .D ( new_AGEMA_signal_9596 ), .Q ( new_AGEMA_signal_9597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5188 ( .C ( clk ), .D ( new_AGEMA_signal_9676 ), .Q ( new_AGEMA_signal_9677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5204 ( .C ( clk ), .D ( new_AGEMA_signal_9692 ), .Q ( new_AGEMA_signal_9693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5220 ( .C ( clk ), .D ( new_AGEMA_signal_9708 ), .Q ( new_AGEMA_signal_9709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5254 ( .C ( clk ), .D ( new_AGEMA_signal_9742 ), .Q ( new_AGEMA_signal_9743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5270 ( .C ( clk ), .D ( new_AGEMA_signal_9758 ), .Q ( new_AGEMA_signal_9759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5286 ( .C ( clk ), .D ( new_AGEMA_signal_9774 ), .Q ( new_AGEMA_signal_9775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5482 ( .C ( clk ), .D ( new_AGEMA_signal_9970 ), .Q ( new_AGEMA_signal_9971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5500 ( .C ( clk ), .D ( new_AGEMA_signal_9988 ), .Q ( new_AGEMA_signal_9989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5518 ( .C ( clk ), .D ( new_AGEMA_signal_10006 ), .Q ( new_AGEMA_signal_10007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5632 ( .C ( clk ), .D ( new_AGEMA_signal_10120 ), .Q ( new_AGEMA_signal_10121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5652 ( .C ( clk ), .D ( new_AGEMA_signal_10140 ), .Q ( new_AGEMA_signal_10141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5672 ( .C ( clk ), .D ( new_AGEMA_signal_10160 ), .Q ( new_AGEMA_signal_10161 ) ) ;

    /* cells in depth 9 */
    buf_clk new_AGEMA_reg_buffer_2555 ( .C ( clk ), .D ( new_AGEMA_signal_7043 ), .Q ( new_AGEMA_signal_7044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2559 ( .C ( clk ), .D ( new_AGEMA_signal_7047 ), .Q ( new_AGEMA_signal_7048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2563 ( .C ( clk ), .D ( new_AGEMA_signal_7051 ), .Q ( new_AGEMA_signal_7052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2567 ( .C ( clk ), .D ( new_AGEMA_signal_7055 ), .Q ( new_AGEMA_signal_7056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2571 ( .C ( clk ), .D ( new_AGEMA_signal_7059 ), .Q ( new_AGEMA_signal_7060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2575 ( .C ( clk ), .D ( new_AGEMA_signal_7063 ), .Q ( new_AGEMA_signal_7064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2583 ( .C ( clk ), .D ( new_AGEMA_signal_7071 ), .Q ( new_AGEMA_signal_7072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2591 ( .C ( clk ), .D ( new_AGEMA_signal_7079 ), .Q ( new_AGEMA_signal_7080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2599 ( .C ( clk ), .D ( new_AGEMA_signal_7087 ), .Q ( new_AGEMA_signal_7088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2601 ( .C ( clk ), .D ( n1978 ), .Q ( new_AGEMA_signal_7090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2603 ( .C ( clk ), .D ( new_AGEMA_signal_2022 ), .Q ( new_AGEMA_signal_7092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2605 ( .C ( clk ), .D ( new_AGEMA_signal_2023 ), .Q ( new_AGEMA_signal_7094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2613 ( .C ( clk ), .D ( new_AGEMA_signal_7101 ), .Q ( new_AGEMA_signal_7102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2621 ( .C ( clk ), .D ( new_AGEMA_signal_7109 ), .Q ( new_AGEMA_signal_7110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2629 ( .C ( clk ), .D ( new_AGEMA_signal_7117 ), .Q ( new_AGEMA_signal_7118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2635 ( .C ( clk ), .D ( new_AGEMA_signal_7123 ), .Q ( new_AGEMA_signal_7124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2641 ( .C ( clk ), .D ( new_AGEMA_signal_7129 ), .Q ( new_AGEMA_signal_7130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2647 ( .C ( clk ), .D ( new_AGEMA_signal_7135 ), .Q ( new_AGEMA_signal_7136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2651 ( .C ( clk ), .D ( new_AGEMA_signal_7139 ), .Q ( new_AGEMA_signal_7140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2655 ( .C ( clk ), .D ( new_AGEMA_signal_7143 ), .Q ( new_AGEMA_signal_7144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2659 ( .C ( clk ), .D ( new_AGEMA_signal_7147 ), .Q ( new_AGEMA_signal_7148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2665 ( .C ( clk ), .D ( new_AGEMA_signal_7153 ), .Q ( new_AGEMA_signal_7154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2671 ( .C ( clk ), .D ( new_AGEMA_signal_7159 ), .Q ( new_AGEMA_signal_7160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2677 ( .C ( clk ), .D ( new_AGEMA_signal_7165 ), .Q ( new_AGEMA_signal_7166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2679 ( .C ( clk ), .D ( new_AGEMA_signal_6877 ), .Q ( new_AGEMA_signal_7168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2681 ( .C ( clk ), .D ( new_AGEMA_signal_6881 ), .Q ( new_AGEMA_signal_7170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2683 ( .C ( clk ), .D ( new_AGEMA_signal_6885 ), .Q ( new_AGEMA_signal_7172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2689 ( .C ( clk ), .D ( new_AGEMA_signal_7177 ), .Q ( new_AGEMA_signal_7178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2695 ( .C ( clk ), .D ( new_AGEMA_signal_7183 ), .Q ( new_AGEMA_signal_7184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2701 ( .C ( clk ), .D ( new_AGEMA_signal_7189 ), .Q ( new_AGEMA_signal_7190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2707 ( .C ( clk ), .D ( new_AGEMA_signal_7195 ), .Q ( new_AGEMA_signal_7196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2713 ( .C ( clk ), .D ( new_AGEMA_signal_7201 ), .Q ( new_AGEMA_signal_7202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2719 ( .C ( clk ), .D ( new_AGEMA_signal_7207 ), .Q ( new_AGEMA_signal_7208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2721 ( .C ( clk ), .D ( n2091 ), .Q ( new_AGEMA_signal_7210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2723 ( .C ( clk ), .D ( new_AGEMA_signal_2058 ), .Q ( new_AGEMA_signal_7212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2725 ( .C ( clk ), .D ( new_AGEMA_signal_2059 ), .Q ( new_AGEMA_signal_7214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2729 ( .C ( clk ), .D ( new_AGEMA_signal_7217 ), .Q ( new_AGEMA_signal_7218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2733 ( .C ( clk ), .D ( new_AGEMA_signal_7221 ), .Q ( new_AGEMA_signal_7222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2737 ( .C ( clk ), .D ( new_AGEMA_signal_7225 ), .Q ( new_AGEMA_signal_7226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2743 ( .C ( clk ), .D ( new_AGEMA_signal_7231 ), .Q ( new_AGEMA_signal_7232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2749 ( .C ( clk ), .D ( new_AGEMA_signal_7237 ), .Q ( new_AGEMA_signal_7238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2755 ( .C ( clk ), .D ( new_AGEMA_signal_7243 ), .Q ( new_AGEMA_signal_7244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2761 ( .C ( clk ), .D ( new_AGEMA_signal_7249 ), .Q ( new_AGEMA_signal_7250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2767 ( .C ( clk ), .D ( new_AGEMA_signal_7255 ), .Q ( new_AGEMA_signal_7256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2773 ( .C ( clk ), .D ( new_AGEMA_signal_7261 ), .Q ( new_AGEMA_signal_7262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2775 ( .C ( clk ), .D ( n2543 ), .Q ( new_AGEMA_signal_7264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2777 ( .C ( clk ), .D ( new_AGEMA_signal_2070 ), .Q ( new_AGEMA_signal_7266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2779 ( .C ( clk ), .D ( new_AGEMA_signal_2071 ), .Q ( new_AGEMA_signal_7268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2785 ( .C ( clk ), .D ( new_AGEMA_signal_7273 ), .Q ( new_AGEMA_signal_7274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2791 ( .C ( clk ), .D ( new_AGEMA_signal_7279 ), .Q ( new_AGEMA_signal_7280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2797 ( .C ( clk ), .D ( new_AGEMA_signal_7285 ), .Q ( new_AGEMA_signal_7286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2799 ( .C ( clk ), .D ( n2159 ), .Q ( new_AGEMA_signal_7288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2801 ( .C ( clk ), .D ( new_AGEMA_signal_2078 ), .Q ( new_AGEMA_signal_7290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2803 ( .C ( clk ), .D ( new_AGEMA_signal_2079 ), .Q ( new_AGEMA_signal_7292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2807 ( .C ( clk ), .D ( new_AGEMA_signal_7295 ), .Q ( new_AGEMA_signal_7296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2811 ( .C ( clk ), .D ( new_AGEMA_signal_7299 ), .Q ( new_AGEMA_signal_7300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2815 ( .C ( clk ), .D ( new_AGEMA_signal_7303 ), .Q ( new_AGEMA_signal_7304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2819 ( .C ( clk ), .D ( new_AGEMA_signal_7307 ), .Q ( new_AGEMA_signal_7308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2823 ( .C ( clk ), .D ( new_AGEMA_signal_7311 ), .Q ( new_AGEMA_signal_7312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2827 ( .C ( clk ), .D ( new_AGEMA_signal_7315 ), .Q ( new_AGEMA_signal_7316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2829 ( .C ( clk ), .D ( new_AGEMA_signal_6857 ), .Q ( new_AGEMA_signal_7318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2831 ( .C ( clk ), .D ( new_AGEMA_signal_6859 ), .Q ( new_AGEMA_signal_7320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2833 ( .C ( clk ), .D ( new_AGEMA_signal_6861 ), .Q ( new_AGEMA_signal_7322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2841 ( .C ( clk ), .D ( new_AGEMA_signal_7329 ), .Q ( new_AGEMA_signal_7330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2849 ( .C ( clk ), .D ( new_AGEMA_signal_7337 ), .Q ( new_AGEMA_signal_7338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2857 ( .C ( clk ), .D ( new_AGEMA_signal_7345 ), .Q ( new_AGEMA_signal_7346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2863 ( .C ( clk ), .D ( new_AGEMA_signal_7351 ), .Q ( new_AGEMA_signal_7352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2869 ( .C ( clk ), .D ( new_AGEMA_signal_7357 ), .Q ( new_AGEMA_signal_7358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2875 ( .C ( clk ), .D ( new_AGEMA_signal_7363 ), .Q ( new_AGEMA_signal_7364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2879 ( .C ( clk ), .D ( new_AGEMA_signal_7367 ), .Q ( new_AGEMA_signal_7368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2883 ( .C ( clk ), .D ( new_AGEMA_signal_7371 ), .Q ( new_AGEMA_signal_7372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2887 ( .C ( clk ), .D ( new_AGEMA_signal_7375 ), .Q ( new_AGEMA_signal_7376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2891 ( .C ( clk ), .D ( new_AGEMA_signal_7379 ), .Q ( new_AGEMA_signal_7380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2895 ( .C ( clk ), .D ( new_AGEMA_signal_7383 ), .Q ( new_AGEMA_signal_7384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2899 ( .C ( clk ), .D ( new_AGEMA_signal_7387 ), .Q ( new_AGEMA_signal_7388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2901 ( .C ( clk ), .D ( n2270 ), .Q ( new_AGEMA_signal_7390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2903 ( .C ( clk ), .D ( new_AGEMA_signal_1830 ), .Q ( new_AGEMA_signal_7392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2905 ( .C ( clk ), .D ( new_AGEMA_signal_1831 ), .Q ( new_AGEMA_signal_7394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2907 ( .C ( clk ), .D ( n2285 ), .Q ( new_AGEMA_signal_7396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2909 ( .C ( clk ), .D ( new_AGEMA_signal_2114 ), .Q ( new_AGEMA_signal_7398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2911 ( .C ( clk ), .D ( new_AGEMA_signal_2115 ), .Q ( new_AGEMA_signal_7400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2915 ( .C ( clk ), .D ( new_AGEMA_signal_7403 ), .Q ( new_AGEMA_signal_7404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2919 ( .C ( clk ), .D ( new_AGEMA_signal_7407 ), .Q ( new_AGEMA_signal_7408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2923 ( .C ( clk ), .D ( new_AGEMA_signal_7411 ), .Q ( new_AGEMA_signal_7412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2927 ( .C ( clk ), .D ( new_AGEMA_signal_7415 ), .Q ( new_AGEMA_signal_7416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2931 ( .C ( clk ), .D ( new_AGEMA_signal_7419 ), .Q ( new_AGEMA_signal_7420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2935 ( .C ( clk ), .D ( new_AGEMA_signal_7423 ), .Q ( new_AGEMA_signal_7424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2937 ( .C ( clk ), .D ( n2334 ), .Q ( new_AGEMA_signal_7426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2939 ( .C ( clk ), .D ( new_AGEMA_signal_1852 ), .Q ( new_AGEMA_signal_7428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2941 ( .C ( clk ), .D ( new_AGEMA_signal_1853 ), .Q ( new_AGEMA_signal_7430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2947 ( .C ( clk ), .D ( new_AGEMA_signal_7435 ), .Q ( new_AGEMA_signal_7436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2953 ( .C ( clk ), .D ( new_AGEMA_signal_7441 ), .Q ( new_AGEMA_signal_7442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2959 ( .C ( clk ), .D ( new_AGEMA_signal_7447 ), .Q ( new_AGEMA_signal_7448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2963 ( .C ( clk ), .D ( new_AGEMA_signal_7451 ), .Q ( new_AGEMA_signal_7452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2967 ( .C ( clk ), .D ( new_AGEMA_signal_7455 ), .Q ( new_AGEMA_signal_7456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2971 ( .C ( clk ), .D ( new_AGEMA_signal_7459 ), .Q ( new_AGEMA_signal_7460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2973 ( .C ( clk ), .D ( new_AGEMA_signal_6869 ), .Q ( new_AGEMA_signal_7462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2975 ( .C ( clk ), .D ( new_AGEMA_signal_6871 ), .Q ( new_AGEMA_signal_7464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2977 ( .C ( clk ), .D ( new_AGEMA_signal_6873 ), .Q ( new_AGEMA_signal_7466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2981 ( .C ( clk ), .D ( new_AGEMA_signal_7469 ), .Q ( new_AGEMA_signal_7470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2985 ( .C ( clk ), .D ( new_AGEMA_signal_7473 ), .Q ( new_AGEMA_signal_7474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2989 ( .C ( clk ), .D ( new_AGEMA_signal_7477 ), .Q ( new_AGEMA_signal_7478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2993 ( .C ( clk ), .D ( new_AGEMA_signal_7481 ), .Q ( new_AGEMA_signal_7482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2997 ( .C ( clk ), .D ( new_AGEMA_signal_7485 ), .Q ( new_AGEMA_signal_7486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3001 ( .C ( clk ), .D ( new_AGEMA_signal_7489 ), .Q ( new_AGEMA_signal_7490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3005 ( .C ( clk ), .D ( new_AGEMA_signal_7493 ), .Q ( new_AGEMA_signal_7494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3009 ( .C ( clk ), .D ( new_AGEMA_signal_7497 ), .Q ( new_AGEMA_signal_7498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3013 ( .C ( clk ), .D ( new_AGEMA_signal_7501 ), .Q ( new_AGEMA_signal_7502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3015 ( .C ( clk ), .D ( n2435 ), .Q ( new_AGEMA_signal_7504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3017 ( .C ( clk ), .D ( new_AGEMA_signal_1890 ), .Q ( new_AGEMA_signal_7506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3019 ( .C ( clk ), .D ( new_AGEMA_signal_1891 ), .Q ( new_AGEMA_signal_7508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3023 ( .C ( clk ), .D ( new_AGEMA_signal_7511 ), .Q ( new_AGEMA_signal_7512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3027 ( .C ( clk ), .D ( new_AGEMA_signal_7515 ), .Q ( new_AGEMA_signal_7516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3031 ( .C ( clk ), .D ( new_AGEMA_signal_7519 ), .Q ( new_AGEMA_signal_7520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3033 ( .C ( clk ), .D ( new_AGEMA_signal_6755 ), .Q ( new_AGEMA_signal_7522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3035 ( .C ( clk ), .D ( new_AGEMA_signal_6757 ), .Q ( new_AGEMA_signal_7524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3037 ( .C ( clk ), .D ( new_AGEMA_signal_6759 ), .Q ( new_AGEMA_signal_7526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3043 ( .C ( clk ), .D ( new_AGEMA_signal_7531 ), .Q ( new_AGEMA_signal_7532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3049 ( .C ( clk ), .D ( new_AGEMA_signal_7537 ), .Q ( new_AGEMA_signal_7538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3055 ( .C ( clk ), .D ( new_AGEMA_signal_7543 ), .Q ( new_AGEMA_signal_7544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3061 ( .C ( clk ), .D ( new_AGEMA_signal_7549 ), .Q ( new_AGEMA_signal_7550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3067 ( .C ( clk ), .D ( new_AGEMA_signal_7555 ), .Q ( new_AGEMA_signal_7556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3073 ( .C ( clk ), .D ( new_AGEMA_signal_7561 ), .Q ( new_AGEMA_signal_7562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3077 ( .C ( clk ), .D ( new_AGEMA_signal_7565 ), .Q ( new_AGEMA_signal_7566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3081 ( .C ( clk ), .D ( new_AGEMA_signal_7569 ), .Q ( new_AGEMA_signal_7570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3085 ( .C ( clk ), .D ( new_AGEMA_signal_7573 ), .Q ( new_AGEMA_signal_7574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3087 ( .C ( clk ), .D ( new_AGEMA_signal_6723 ), .Q ( new_AGEMA_signal_7576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3089 ( .C ( clk ), .D ( new_AGEMA_signal_6729 ), .Q ( new_AGEMA_signal_7578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3091 ( .C ( clk ), .D ( new_AGEMA_signal_6735 ), .Q ( new_AGEMA_signal_7580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3099 ( .C ( clk ), .D ( new_AGEMA_signal_7587 ), .Q ( new_AGEMA_signal_7588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3107 ( .C ( clk ), .D ( new_AGEMA_signal_7595 ), .Q ( new_AGEMA_signal_7596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3115 ( .C ( clk ), .D ( new_AGEMA_signal_7603 ), .Q ( new_AGEMA_signal_7604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3117 ( .C ( clk ), .D ( n2547 ), .Q ( new_AGEMA_signal_7606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3119 ( .C ( clk ), .D ( new_AGEMA_signal_1926 ), .Q ( new_AGEMA_signal_7608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3121 ( .C ( clk ), .D ( new_AGEMA_signal_1927 ), .Q ( new_AGEMA_signal_7610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3125 ( .C ( clk ), .D ( new_AGEMA_signal_7613 ), .Q ( new_AGEMA_signal_7614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3129 ( .C ( clk ), .D ( new_AGEMA_signal_7617 ), .Q ( new_AGEMA_signal_7618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3133 ( .C ( clk ), .D ( new_AGEMA_signal_7621 ), .Q ( new_AGEMA_signal_7622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3137 ( .C ( clk ), .D ( new_AGEMA_signal_7625 ), .Q ( new_AGEMA_signal_7626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3141 ( .C ( clk ), .D ( new_AGEMA_signal_7629 ), .Q ( new_AGEMA_signal_7630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3145 ( .C ( clk ), .D ( new_AGEMA_signal_7633 ), .Q ( new_AGEMA_signal_7634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3149 ( .C ( clk ), .D ( new_AGEMA_signal_7637 ), .Q ( new_AGEMA_signal_7638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3153 ( .C ( clk ), .D ( new_AGEMA_signal_7641 ), .Q ( new_AGEMA_signal_7642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3157 ( .C ( clk ), .D ( new_AGEMA_signal_7645 ), .Q ( new_AGEMA_signal_7646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3161 ( .C ( clk ), .D ( new_AGEMA_signal_7649 ), .Q ( new_AGEMA_signal_7650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3165 ( .C ( clk ), .D ( new_AGEMA_signal_7653 ), .Q ( new_AGEMA_signal_7654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3169 ( .C ( clk ), .D ( new_AGEMA_signal_7657 ), .Q ( new_AGEMA_signal_7658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3173 ( .C ( clk ), .D ( new_AGEMA_signal_7661 ), .Q ( new_AGEMA_signal_7662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3177 ( .C ( clk ), .D ( new_AGEMA_signal_7665 ), .Q ( new_AGEMA_signal_7666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3181 ( .C ( clk ), .D ( new_AGEMA_signal_7669 ), .Q ( new_AGEMA_signal_7670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3189 ( .C ( clk ), .D ( new_AGEMA_signal_7677 ), .Q ( new_AGEMA_signal_7678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3197 ( .C ( clk ), .D ( new_AGEMA_signal_7685 ), .Q ( new_AGEMA_signal_7686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3205 ( .C ( clk ), .D ( new_AGEMA_signal_7693 ), .Q ( new_AGEMA_signal_7694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3207 ( .C ( clk ), .D ( n2758 ), .Q ( new_AGEMA_signal_7696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3209 ( .C ( clk ), .D ( new_AGEMA_signal_2216 ), .Q ( new_AGEMA_signal_7698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3211 ( .C ( clk ), .D ( new_AGEMA_signal_2217 ), .Q ( new_AGEMA_signal_7700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3215 ( .C ( clk ), .D ( new_AGEMA_signal_7703 ), .Q ( new_AGEMA_signal_7704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3219 ( .C ( clk ), .D ( new_AGEMA_signal_7707 ), .Q ( new_AGEMA_signal_7708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3223 ( .C ( clk ), .D ( new_AGEMA_signal_7711 ), .Q ( new_AGEMA_signal_7712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3225 ( .C ( clk ), .D ( n2797 ), .Q ( new_AGEMA_signal_7714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3227 ( .C ( clk ), .D ( new_AGEMA_signal_2224 ), .Q ( new_AGEMA_signal_7716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3229 ( .C ( clk ), .D ( new_AGEMA_signal_2225 ), .Q ( new_AGEMA_signal_7718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3235 ( .C ( clk ), .D ( new_AGEMA_signal_7723 ), .Q ( new_AGEMA_signal_7724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3241 ( .C ( clk ), .D ( new_AGEMA_signal_7729 ), .Q ( new_AGEMA_signal_7730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3247 ( .C ( clk ), .D ( new_AGEMA_signal_7735 ), .Q ( new_AGEMA_signal_7736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3259 ( .C ( clk ), .D ( new_AGEMA_signal_7747 ), .Q ( new_AGEMA_signal_7748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3267 ( .C ( clk ), .D ( new_AGEMA_signal_7755 ), .Q ( new_AGEMA_signal_7756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3275 ( .C ( clk ), .D ( new_AGEMA_signal_7763 ), .Q ( new_AGEMA_signal_7764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3285 ( .C ( clk ), .D ( n2012 ), .Q ( new_AGEMA_signal_7774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3289 ( .C ( clk ), .D ( new_AGEMA_signal_2032 ), .Q ( new_AGEMA_signal_7778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3293 ( .C ( clk ), .D ( new_AGEMA_signal_2033 ), .Q ( new_AGEMA_signal_7782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3301 ( .C ( clk ), .D ( new_AGEMA_signal_7789 ), .Q ( new_AGEMA_signal_7790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3309 ( .C ( clk ), .D ( new_AGEMA_signal_7797 ), .Q ( new_AGEMA_signal_7798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3317 ( .C ( clk ), .D ( new_AGEMA_signal_7805 ), .Q ( new_AGEMA_signal_7806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3329 ( .C ( clk ), .D ( new_AGEMA_signal_7817 ), .Q ( new_AGEMA_signal_7818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3335 ( .C ( clk ), .D ( new_AGEMA_signal_7823 ), .Q ( new_AGEMA_signal_7824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3341 ( .C ( clk ), .D ( new_AGEMA_signal_7829 ), .Q ( new_AGEMA_signal_7830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3345 ( .C ( clk ), .D ( n2652 ), .Q ( new_AGEMA_signal_7834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3349 ( .C ( clk ), .D ( new_AGEMA_signal_2050 ), .Q ( new_AGEMA_signal_7838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3353 ( .C ( clk ), .D ( new_AGEMA_signal_2051 ), .Q ( new_AGEMA_signal_7842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3361 ( .C ( clk ), .D ( new_AGEMA_signal_7849 ), .Q ( new_AGEMA_signal_7850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3369 ( .C ( clk ), .D ( new_AGEMA_signal_7857 ), .Q ( new_AGEMA_signal_7858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3377 ( .C ( clk ), .D ( new_AGEMA_signal_7865 ), .Q ( new_AGEMA_signal_7866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3381 ( .C ( clk ), .D ( n2143 ), .Q ( new_AGEMA_signal_7870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3385 ( .C ( clk ), .D ( new_AGEMA_signal_2074 ), .Q ( new_AGEMA_signal_7874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3389 ( .C ( clk ), .D ( new_AGEMA_signal_2075 ), .Q ( new_AGEMA_signal_7878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3395 ( .C ( clk ), .D ( new_AGEMA_signal_7883 ), .Q ( new_AGEMA_signal_7884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3401 ( .C ( clk ), .D ( new_AGEMA_signal_7889 ), .Q ( new_AGEMA_signal_7890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3407 ( .C ( clk ), .D ( new_AGEMA_signal_7895 ), .Q ( new_AGEMA_signal_7896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3413 ( .C ( clk ), .D ( new_AGEMA_signal_7901 ), .Q ( new_AGEMA_signal_7902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3419 ( .C ( clk ), .D ( new_AGEMA_signal_7907 ), .Q ( new_AGEMA_signal_7908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3425 ( .C ( clk ), .D ( new_AGEMA_signal_7913 ), .Q ( new_AGEMA_signal_7914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3431 ( .C ( clk ), .D ( new_AGEMA_signal_7919 ), .Q ( new_AGEMA_signal_7920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3437 ( .C ( clk ), .D ( new_AGEMA_signal_7925 ), .Q ( new_AGEMA_signal_7926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3443 ( .C ( clk ), .D ( new_AGEMA_signal_7931 ), .Q ( new_AGEMA_signal_7932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3449 ( .C ( clk ), .D ( new_AGEMA_signal_7937 ), .Q ( new_AGEMA_signal_7938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3455 ( .C ( clk ), .D ( new_AGEMA_signal_7943 ), .Q ( new_AGEMA_signal_7944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3461 ( .C ( clk ), .D ( new_AGEMA_signal_7949 ), .Q ( new_AGEMA_signal_7950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3467 ( .C ( clk ), .D ( new_AGEMA_signal_7955 ), .Q ( new_AGEMA_signal_7956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3473 ( .C ( clk ), .D ( new_AGEMA_signal_7961 ), .Q ( new_AGEMA_signal_7962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3479 ( .C ( clk ), .D ( new_AGEMA_signal_7967 ), .Q ( new_AGEMA_signal_7968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3483 ( .C ( clk ), .D ( n2297 ), .Q ( new_AGEMA_signal_7972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3487 ( .C ( clk ), .D ( new_AGEMA_signal_2120 ), .Q ( new_AGEMA_signal_7976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3491 ( .C ( clk ), .D ( new_AGEMA_signal_2121 ), .Q ( new_AGEMA_signal_7980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3499 ( .C ( clk ), .D ( new_AGEMA_signal_7987 ), .Q ( new_AGEMA_signal_7988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3507 ( .C ( clk ), .D ( new_AGEMA_signal_7995 ), .Q ( new_AGEMA_signal_7996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3515 ( .C ( clk ), .D ( new_AGEMA_signal_8003 ), .Q ( new_AGEMA_signal_8004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3519 ( .C ( clk ), .D ( n2336 ), .Q ( new_AGEMA_signal_8008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3523 ( .C ( clk ), .D ( new_AGEMA_signal_2310 ), .Q ( new_AGEMA_signal_8012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3527 ( .C ( clk ), .D ( new_AGEMA_signal_2311 ), .Q ( new_AGEMA_signal_8016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3533 ( .C ( clk ), .D ( new_AGEMA_signal_8021 ), .Q ( new_AGEMA_signal_8022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3539 ( .C ( clk ), .D ( new_AGEMA_signal_8027 ), .Q ( new_AGEMA_signal_8028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3545 ( .C ( clk ), .D ( new_AGEMA_signal_8033 ), .Q ( new_AGEMA_signal_8034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3553 ( .C ( clk ), .D ( new_AGEMA_signal_8041 ), .Q ( new_AGEMA_signal_8042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3561 ( .C ( clk ), .D ( new_AGEMA_signal_8049 ), .Q ( new_AGEMA_signal_8050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3569 ( .C ( clk ), .D ( new_AGEMA_signal_8057 ), .Q ( new_AGEMA_signal_8058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3581 ( .C ( clk ), .D ( new_AGEMA_signal_8069 ), .Q ( new_AGEMA_signal_8070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3587 ( .C ( clk ), .D ( new_AGEMA_signal_8075 ), .Q ( new_AGEMA_signal_8076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3593 ( .C ( clk ), .D ( new_AGEMA_signal_8081 ), .Q ( new_AGEMA_signal_8082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3611 ( .C ( clk ), .D ( new_AGEMA_signal_8099 ), .Q ( new_AGEMA_signal_8100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3617 ( .C ( clk ), .D ( new_AGEMA_signal_8105 ), .Q ( new_AGEMA_signal_8106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3623 ( .C ( clk ), .D ( new_AGEMA_signal_8111 ), .Q ( new_AGEMA_signal_8112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3629 ( .C ( clk ), .D ( new_AGEMA_signal_8117 ), .Q ( new_AGEMA_signal_8118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3635 ( .C ( clk ), .D ( new_AGEMA_signal_8123 ), .Q ( new_AGEMA_signal_8124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3641 ( .C ( clk ), .D ( new_AGEMA_signal_8129 ), .Q ( new_AGEMA_signal_8130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3649 ( .C ( clk ), .D ( new_AGEMA_signal_8137 ), .Q ( new_AGEMA_signal_8138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3657 ( .C ( clk ), .D ( new_AGEMA_signal_8145 ), .Q ( new_AGEMA_signal_8146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3665 ( .C ( clk ), .D ( new_AGEMA_signal_8153 ), .Q ( new_AGEMA_signal_8154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3673 ( .C ( clk ), .D ( new_AGEMA_signal_8161 ), .Q ( new_AGEMA_signal_8162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3681 ( .C ( clk ), .D ( new_AGEMA_signal_8169 ), .Q ( new_AGEMA_signal_8170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3689 ( .C ( clk ), .D ( new_AGEMA_signal_8177 ), .Q ( new_AGEMA_signal_8178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3695 ( .C ( clk ), .D ( new_AGEMA_signal_8183 ), .Q ( new_AGEMA_signal_8184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3701 ( .C ( clk ), .D ( new_AGEMA_signal_8189 ), .Q ( new_AGEMA_signal_8190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3707 ( .C ( clk ), .D ( new_AGEMA_signal_8195 ), .Q ( new_AGEMA_signal_8196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3713 ( .C ( clk ), .D ( new_AGEMA_signal_8201 ), .Q ( new_AGEMA_signal_8202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3719 ( .C ( clk ), .D ( new_AGEMA_signal_8207 ), .Q ( new_AGEMA_signal_8208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3725 ( .C ( clk ), .D ( new_AGEMA_signal_8213 ), .Q ( new_AGEMA_signal_8214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3735 ( .C ( clk ), .D ( n2658 ), .Q ( new_AGEMA_signal_8224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3739 ( .C ( clk ), .D ( new_AGEMA_signal_2014 ), .Q ( new_AGEMA_signal_8228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3743 ( .C ( clk ), .D ( new_AGEMA_signal_2015 ), .Q ( new_AGEMA_signal_8232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3747 ( .C ( clk ), .D ( n2698 ), .Q ( new_AGEMA_signal_8236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3751 ( .C ( clk ), .D ( new_AGEMA_signal_2204 ), .Q ( new_AGEMA_signal_8240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3755 ( .C ( clk ), .D ( new_AGEMA_signal_2205 ), .Q ( new_AGEMA_signal_8244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3759 ( .C ( clk ), .D ( n2800 ), .Q ( new_AGEMA_signal_8248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3763 ( .C ( clk ), .D ( new_AGEMA_signal_2220 ), .Q ( new_AGEMA_signal_8252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3767 ( .C ( clk ), .D ( new_AGEMA_signal_2221 ), .Q ( new_AGEMA_signal_8256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3777 ( .C ( clk ), .D ( n1936 ), .Q ( new_AGEMA_signal_8266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3783 ( .C ( clk ), .D ( new_AGEMA_signal_1998 ), .Q ( new_AGEMA_signal_8272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3789 ( .C ( clk ), .D ( new_AGEMA_signal_1999 ), .Q ( new_AGEMA_signal_8278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3815 ( .C ( clk ), .D ( new_AGEMA_signal_8303 ), .Q ( new_AGEMA_signal_8304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3823 ( .C ( clk ), .D ( new_AGEMA_signal_8311 ), .Q ( new_AGEMA_signal_8312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3831 ( .C ( clk ), .D ( new_AGEMA_signal_8319 ), .Q ( new_AGEMA_signal_8320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3839 ( .C ( clk ), .D ( new_AGEMA_signal_8327 ), .Q ( new_AGEMA_signal_8328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3847 ( .C ( clk ), .D ( new_AGEMA_signal_8335 ), .Q ( new_AGEMA_signal_8336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3855 ( .C ( clk ), .D ( new_AGEMA_signal_8343 ), .Q ( new_AGEMA_signal_8344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3863 ( .C ( clk ), .D ( new_AGEMA_signal_8351 ), .Q ( new_AGEMA_signal_8352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3871 ( .C ( clk ), .D ( new_AGEMA_signal_8359 ), .Q ( new_AGEMA_signal_8360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3879 ( .C ( clk ), .D ( new_AGEMA_signal_8367 ), .Q ( new_AGEMA_signal_8368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3887 ( .C ( clk ), .D ( new_AGEMA_signal_8375 ), .Q ( new_AGEMA_signal_8376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3895 ( .C ( clk ), .D ( new_AGEMA_signal_8383 ), .Q ( new_AGEMA_signal_8384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3903 ( .C ( clk ), .D ( new_AGEMA_signal_8391 ), .Q ( new_AGEMA_signal_8392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3909 ( .C ( clk ), .D ( n2099 ), .Q ( new_AGEMA_signal_8398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3915 ( .C ( clk ), .D ( new_AGEMA_signal_2056 ), .Q ( new_AGEMA_signal_8404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3921 ( .C ( clk ), .D ( new_AGEMA_signal_2057 ), .Q ( new_AGEMA_signal_8410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3931 ( .C ( clk ), .D ( new_AGEMA_signal_8419 ), .Q ( new_AGEMA_signal_8420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3941 ( .C ( clk ), .D ( new_AGEMA_signal_8429 ), .Q ( new_AGEMA_signal_8430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3951 ( .C ( clk ), .D ( new_AGEMA_signal_8439 ), .Q ( new_AGEMA_signal_8440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3959 ( .C ( clk ), .D ( new_AGEMA_signal_8447 ), .Q ( new_AGEMA_signal_8448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3967 ( .C ( clk ), .D ( new_AGEMA_signal_8455 ), .Q ( new_AGEMA_signal_8456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3975 ( .C ( clk ), .D ( new_AGEMA_signal_8463 ), .Q ( new_AGEMA_signal_8464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3983 ( .C ( clk ), .D ( new_AGEMA_signal_8471 ), .Q ( new_AGEMA_signal_8472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3991 ( .C ( clk ), .D ( new_AGEMA_signal_8479 ), .Q ( new_AGEMA_signal_8480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3999 ( .C ( clk ), .D ( new_AGEMA_signal_8487 ), .Q ( new_AGEMA_signal_8488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4007 ( .C ( clk ), .D ( new_AGEMA_signal_8495 ), .Q ( new_AGEMA_signal_8496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4015 ( .C ( clk ), .D ( new_AGEMA_signal_8503 ), .Q ( new_AGEMA_signal_8504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4023 ( .C ( clk ), .D ( new_AGEMA_signal_8511 ), .Q ( new_AGEMA_signal_8512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4047 ( .C ( clk ), .D ( n2301 ), .Q ( new_AGEMA_signal_8536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4053 ( .C ( clk ), .D ( new_AGEMA_signal_2124 ), .Q ( new_AGEMA_signal_8542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4059 ( .C ( clk ), .D ( new_AGEMA_signal_2125 ), .Q ( new_AGEMA_signal_8548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4081 ( .C ( clk ), .D ( new_AGEMA_signal_8569 ), .Q ( new_AGEMA_signal_8570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4091 ( .C ( clk ), .D ( new_AGEMA_signal_8579 ), .Q ( new_AGEMA_signal_8580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4101 ( .C ( clk ), .D ( new_AGEMA_signal_8589 ), .Q ( new_AGEMA_signal_8590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4109 ( .C ( clk ), .D ( new_AGEMA_signal_8597 ), .Q ( new_AGEMA_signal_8598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4117 ( .C ( clk ), .D ( new_AGEMA_signal_8605 ), .Q ( new_AGEMA_signal_8606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4125 ( .C ( clk ), .D ( new_AGEMA_signal_8613 ), .Q ( new_AGEMA_signal_8614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4151 ( .C ( clk ), .D ( new_AGEMA_signal_8639 ), .Q ( new_AGEMA_signal_8640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4159 ( .C ( clk ), .D ( new_AGEMA_signal_8647 ), .Q ( new_AGEMA_signal_8648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4167 ( .C ( clk ), .D ( new_AGEMA_signal_8655 ), .Q ( new_AGEMA_signal_8656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4175 ( .C ( clk ), .D ( new_AGEMA_signal_8663 ), .Q ( new_AGEMA_signal_8664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4183 ( .C ( clk ), .D ( new_AGEMA_signal_8671 ), .Q ( new_AGEMA_signal_8672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4191 ( .C ( clk ), .D ( new_AGEMA_signal_8679 ), .Q ( new_AGEMA_signal_8680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4197 ( .C ( clk ), .D ( new_AGEMA_signal_6673 ), .Q ( new_AGEMA_signal_8686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4203 ( .C ( clk ), .D ( new_AGEMA_signal_6677 ), .Q ( new_AGEMA_signal_8692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4209 ( .C ( clk ), .D ( new_AGEMA_signal_6681 ), .Q ( new_AGEMA_signal_8698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4229 ( .C ( clk ), .D ( new_AGEMA_signal_8717 ), .Q ( new_AGEMA_signal_8718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4237 ( .C ( clk ), .D ( new_AGEMA_signal_8725 ), .Q ( new_AGEMA_signal_8726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4245 ( .C ( clk ), .D ( new_AGEMA_signal_8733 ), .Q ( new_AGEMA_signal_8734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4323 ( .C ( clk ), .D ( new_AGEMA_signal_7009 ), .Q ( new_AGEMA_signal_8812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4331 ( .C ( clk ), .D ( new_AGEMA_signal_7013 ), .Q ( new_AGEMA_signal_8820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4339 ( .C ( clk ), .D ( new_AGEMA_signal_7017 ), .Q ( new_AGEMA_signal_8828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4377 ( .C ( clk ), .D ( n2102 ), .Q ( new_AGEMA_signal_8866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4385 ( .C ( clk ), .D ( new_AGEMA_signal_2064 ), .Q ( new_AGEMA_signal_8874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4393 ( .C ( clk ), .D ( new_AGEMA_signal_2065 ), .Q ( new_AGEMA_signal_8882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4401 ( .C ( clk ), .D ( new_AGEMA_signal_6551 ), .Q ( new_AGEMA_signal_8890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4409 ( .C ( clk ), .D ( new_AGEMA_signal_6553 ), .Q ( new_AGEMA_signal_8898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4417 ( .C ( clk ), .D ( new_AGEMA_signal_6555 ), .Q ( new_AGEMA_signal_8906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4427 ( .C ( clk ), .D ( new_AGEMA_signal_8915 ), .Q ( new_AGEMA_signal_8916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4437 ( .C ( clk ), .D ( new_AGEMA_signal_8925 ), .Q ( new_AGEMA_signal_8926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4447 ( .C ( clk ), .D ( new_AGEMA_signal_8935 ), .Q ( new_AGEMA_signal_8936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4455 ( .C ( clk ), .D ( new_AGEMA_signal_6829 ), .Q ( new_AGEMA_signal_8944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4463 ( .C ( clk ), .D ( new_AGEMA_signal_6833 ), .Q ( new_AGEMA_signal_8952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4471 ( .C ( clk ), .D ( new_AGEMA_signal_6837 ), .Q ( new_AGEMA_signal_8960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4527 ( .C ( clk ), .D ( n2367 ), .Q ( new_AGEMA_signal_9016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4535 ( .C ( clk ), .D ( new_AGEMA_signal_1858 ), .Q ( new_AGEMA_signal_9024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4543 ( .C ( clk ), .D ( new_AGEMA_signal_1859 ), .Q ( new_AGEMA_signal_9032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4575 ( .C ( clk ), .D ( n2591 ), .Q ( new_AGEMA_signal_9064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4583 ( .C ( clk ), .D ( new_AGEMA_signal_2186 ), .Q ( new_AGEMA_signal_9072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4591 ( .C ( clk ), .D ( new_AGEMA_signal_2187 ), .Q ( new_AGEMA_signal_9080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4707 ( .C ( clk ), .D ( n2105 ), .Q ( new_AGEMA_signal_9196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4717 ( .C ( clk ), .D ( new_AGEMA_signal_2054 ), .Q ( new_AGEMA_signal_9206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4727 ( .C ( clk ), .D ( new_AGEMA_signal_2055 ), .Q ( new_AGEMA_signal_9216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4977 ( .C ( clk ), .D ( n2106 ), .Q ( new_AGEMA_signal_9466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4989 ( .C ( clk ), .D ( new_AGEMA_signal_1772 ), .Q ( new_AGEMA_signal_9478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5001 ( .C ( clk ), .D ( new_AGEMA_signal_1773 ), .Q ( new_AGEMA_signal_9490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5015 ( .C ( clk ), .D ( new_AGEMA_signal_9503 ), .Q ( new_AGEMA_signal_9504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5029 ( .C ( clk ), .D ( new_AGEMA_signal_9517 ), .Q ( new_AGEMA_signal_9518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5043 ( .C ( clk ), .D ( new_AGEMA_signal_9531 ), .Q ( new_AGEMA_signal_9532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5081 ( .C ( clk ), .D ( new_AGEMA_signal_9569 ), .Q ( new_AGEMA_signal_9570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5095 ( .C ( clk ), .D ( new_AGEMA_signal_9583 ), .Q ( new_AGEMA_signal_9584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5109 ( .C ( clk ), .D ( new_AGEMA_signal_9597 ), .Q ( new_AGEMA_signal_9598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5189 ( .C ( clk ), .D ( new_AGEMA_signal_9677 ), .Q ( new_AGEMA_signal_9678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5205 ( .C ( clk ), .D ( new_AGEMA_signal_9693 ), .Q ( new_AGEMA_signal_9694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5221 ( .C ( clk ), .D ( new_AGEMA_signal_9709 ), .Q ( new_AGEMA_signal_9710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5255 ( .C ( clk ), .D ( new_AGEMA_signal_9743 ), .Q ( new_AGEMA_signal_9744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5271 ( .C ( clk ), .D ( new_AGEMA_signal_9759 ), .Q ( new_AGEMA_signal_9760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5287 ( .C ( clk ), .D ( new_AGEMA_signal_9775 ), .Q ( new_AGEMA_signal_9776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5403 ( .C ( clk ), .D ( n2155 ), .Q ( new_AGEMA_signal_9892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5419 ( .C ( clk ), .D ( new_AGEMA_signal_1776 ), .Q ( new_AGEMA_signal_9908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5435 ( .C ( clk ), .D ( new_AGEMA_signal_1777 ), .Q ( new_AGEMA_signal_9924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5483 ( .C ( clk ), .D ( new_AGEMA_signal_9971 ), .Q ( new_AGEMA_signal_9972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5501 ( .C ( clk ), .D ( new_AGEMA_signal_9989 ), .Q ( new_AGEMA_signal_9990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5519 ( .C ( clk ), .D ( new_AGEMA_signal_10007 ), .Q ( new_AGEMA_signal_10008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5633 ( .C ( clk ), .D ( new_AGEMA_signal_10121 ), .Q ( new_AGEMA_signal_10122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5653 ( .C ( clk ), .D ( new_AGEMA_signal_10141 ), .Q ( new_AGEMA_signal_10142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5673 ( .C ( clk ), .D ( new_AGEMA_signal_10161 ), .Q ( new_AGEMA_signal_10162 ) ) ;

    /* cells in depth 10 */
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1983 ( .a ({new_AGEMA_signal_6447, new_AGEMA_signal_6443, new_AGEMA_signal_6439}), .b ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, n1928}), .clk ( clk ), .r ({Fresh[1727], Fresh[1726], Fresh[1725]}), .c ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, n1934}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U1998 ( .a ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, n1931}), .b ({new_AGEMA_signal_6459, new_AGEMA_signal_6455, new_AGEMA_signal_6451}), .clk ( clk ), .r ({Fresh[1730], Fresh[1729], Fresh[1728]}), .c ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, n1932}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2015 ( .a ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, n1939}), .b ({new_AGEMA_signal_6465, new_AGEMA_signal_6463, new_AGEMA_signal_6461}), .clk ( clk ), .r ({Fresh[1733], Fresh[1732], Fresh[1731]}), .c ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, n1940}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2033 ( .a ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, n1948}), .b ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, n1947}), .clk ( clk ), .r ({Fresh[1736], Fresh[1735], Fresh[1734]}), .c ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, n1961}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2050 ( .a ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, n1954}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, n1953}), .clk ( clk ), .r ({Fresh[1739], Fresh[1738], Fresh[1737]}), .c ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, n1955}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2066 ( .a ({new_AGEMA_signal_6471, new_AGEMA_signal_6469, new_AGEMA_signal_6467}), .b ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, n1965}), .clk ( clk ), .r ({Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, n1967}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2085 ( .a ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, n1970}), .b ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, n1969}), .clk ( clk ), .r ({Fresh[1745], Fresh[1744], Fresh[1743]}), .c ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, n1984}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2103 ( .a ({new_AGEMA_signal_6483, new_AGEMA_signal_6479, new_AGEMA_signal_6475}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, n1975}), .clk ( clk ), .r ({Fresh[1748], Fresh[1747], Fresh[1746]}), .c ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, n1977}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2108 ( .a ({new_AGEMA_signal_6489, new_AGEMA_signal_6487, new_AGEMA_signal_6485}), .b ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, n1980}), .clk ( clk ), .r ({Fresh[1751], Fresh[1750], Fresh[1749]}), .c ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, n1981}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2115 ( .a ({new_AGEMA_signal_6501, new_AGEMA_signal_6497, new_AGEMA_signal_6493}), .b ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, n1986}), .clk ( clk ), .r ({Fresh[1754], Fresh[1753], Fresh[1752]}), .c ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, n1987}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2127 ( .a ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, n1997}), .b ({new_AGEMA_signal_6507, new_AGEMA_signal_6505, new_AGEMA_signal_6503}), .clk ( clk ), .r ({Fresh[1757], Fresh[1756], Fresh[1755]}), .c ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, n1998}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2146 ( .a ({new_AGEMA_signal_6519, new_AGEMA_signal_6515, new_AGEMA_signal_6511}), .b ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, n2007}), .clk ( clk ), .r ({Fresh[1760], Fresh[1759], Fresh[1758]}), .c ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, n2010}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2162 ( .a ({new_AGEMA_signal_6531, new_AGEMA_signal_6527, new_AGEMA_signal_6523}), .b ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, n2021}), .clk ( clk ), .r ({Fresh[1763], Fresh[1762], Fresh[1761]}), .c ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, n2024}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2177 ( .a ({new_AGEMA_signal_6537, new_AGEMA_signal_6535, new_AGEMA_signal_6533}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, n2032}), .clk ( clk ), .r ({Fresh[1766], Fresh[1765], Fresh[1764]}), .c ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, n2035}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2186 ( .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, n2041}), .b ({new_AGEMA_signal_6543, new_AGEMA_signal_6541, new_AGEMA_signal_6539}), .clk ( clk ), .r ({Fresh[1769], Fresh[1768], Fresh[1767]}), .c ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, n2054}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2190 ( .a ({new_AGEMA_signal_6549, new_AGEMA_signal_6547, new_AGEMA_signal_6545}), .b ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, n2043}), .clk ( clk ), .r ({Fresh[1772], Fresh[1771], Fresh[1770]}), .c ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, n2048}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2195 ( .a ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, n2046}), .b ({new_AGEMA_signal_6555, new_AGEMA_signal_6553, new_AGEMA_signal_6551}), .clk ( clk ), .r ({Fresh[1775], Fresh[1774], Fresh[1773]}), .c ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, n2047}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2206 ( .a ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, n2058}), .b ({new_AGEMA_signal_6567, new_AGEMA_signal_6563, new_AGEMA_signal_6559}), .clk ( clk ), .r ({Fresh[1778], Fresh[1777], Fresh[1776]}), .c ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, n2059}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2213 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, n2063}), .b ({new_AGEMA_signal_6579, new_AGEMA_signal_6575, new_AGEMA_signal_6571}), .clk ( clk ), .r ({Fresh[1781], Fresh[1780], Fresh[1779]}), .c ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, n2064}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2229 ( .a ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, n2076}), .b ({new_AGEMA_signal_6591, new_AGEMA_signal_6587, new_AGEMA_signal_6583}), .clk ( clk ), .r ({Fresh[1784], Fresh[1783], Fresh[1782]}), .c ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, n2077}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2249 ( .a ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, n2090}), .b ({new_AGEMA_signal_6597, new_AGEMA_signal_6595, new_AGEMA_signal_6593}), .clk ( clk ), .r ({Fresh[1787], Fresh[1786], Fresh[1785]}), .c ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, n2158}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2255 ( .a ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, n2093}), .b ({new_AGEMA_signal_6603, new_AGEMA_signal_6601, new_AGEMA_signal_6599}), .clk ( clk ), .r ({Fresh[1790], Fresh[1789], Fresh[1788]}), .c ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, n2095}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2274 ( .a ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, n2116}), .b ({new_AGEMA_signal_6609, new_AGEMA_signal_6607, new_AGEMA_signal_6605}), .clk ( clk ), .r ({Fresh[1793], Fresh[1792], Fresh[1791]}), .c ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, n2117}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2283 ( .a ({new_AGEMA_signal_6621, new_AGEMA_signal_6617, new_AGEMA_signal_6613}), .b ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, n2120}), .clk ( clk ), .r ({Fresh[1796], Fresh[1795], Fresh[1794]}), .c ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, n2123}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2300 ( .a ({new_AGEMA_signal_6627, new_AGEMA_signal_6625, new_AGEMA_signal_6623}), .b ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, n2134}), .clk ( clk ), .r ({Fresh[1799], Fresh[1798], Fresh[1797]}), .c ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, n2135}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2309 ( .a ({new_AGEMA_signal_6639, new_AGEMA_signal_6635, new_AGEMA_signal_6631}), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, n2140}), .clk ( clk ), .r ({Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, n2141}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2327 ( .a ({new_AGEMA_signal_6657, new_AGEMA_signal_6651, new_AGEMA_signal_6645}), .b ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, n2161}), .clk ( clk ), .r ({Fresh[1805], Fresh[1804], Fresh[1803]}), .c ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, n2166}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2331 ( .a ({new_AGEMA_signal_6669, new_AGEMA_signal_6665, new_AGEMA_signal_6661}), .b ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, n2164}), .clk ( clk ), .r ({Fresh[1808], Fresh[1807], Fresh[1806]}), .c ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, n2165}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2346 ( .a ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, n2179}), .b ({new_AGEMA_signal_6681, new_AGEMA_signal_6677, new_AGEMA_signal_6673}), .clk ( clk ), .r ({Fresh[1811], Fresh[1810], Fresh[1809]}), .c ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, n2180}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2360 ( .a ({new_AGEMA_signal_6687, new_AGEMA_signal_6685, new_AGEMA_signal_6683}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, n2192}), .clk ( clk ), .r ({Fresh[1814], Fresh[1813], Fresh[1812]}), .c ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, n2194}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2372 ( .a ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, n2203}), .b ({new_AGEMA_signal_6693, new_AGEMA_signal_6691, new_AGEMA_signal_6689}), .clk ( clk ), .r ({Fresh[1817], Fresh[1816], Fresh[1815]}), .c ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, n2204}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2389 ( .a ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, n2224}), .b ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, n2223}), .clk ( clk ), .r ({Fresh[1820], Fresh[1819], Fresh[1818]}), .c ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, n2225}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2394 ( .a ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, n2229}), .b ({new_AGEMA_signal_6699, new_AGEMA_signal_6697, new_AGEMA_signal_6695}), .clk ( clk ), .r ({Fresh[1823], Fresh[1822], Fresh[1821]}), .c ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, n2230}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2400 ( .a ({new_AGEMA_signal_6705, new_AGEMA_signal_6703, new_AGEMA_signal_6701}), .b ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, n2234}), .clk ( clk ), .r ({Fresh[1826], Fresh[1825], Fresh[1824]}), .c ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, n2236}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2412 ( .a ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, n2246}), .b ({new_AGEMA_signal_6717, new_AGEMA_signal_6713, new_AGEMA_signal_6709}), .clk ( clk ), .r ({Fresh[1829], Fresh[1828], Fresh[1827]}), .c ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, n2247}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2419 ( .a ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, n2254}), .b ({new_AGEMA_signal_6735, new_AGEMA_signal_6729, new_AGEMA_signal_6723}), .clk ( clk ), .r ({Fresh[1832], Fresh[1831], Fresh[1830]}), .c ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, n2255}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2427 ( .a ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, n2263}), .b ({new_AGEMA_signal_6747, new_AGEMA_signal_6743, new_AGEMA_signal_6739}), .clk ( clk ), .r ({Fresh[1835], Fresh[1834], Fresh[1833]}), .c ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, n2264}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2435 ( .a ({new_AGEMA_signal_6753, new_AGEMA_signal_6751, new_AGEMA_signal_6749}), .b ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, n2267}), .clk ( clk ), .r ({Fresh[1838], Fresh[1837], Fresh[1836]}), .c ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, n2271}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2446 ( .a ({new_AGEMA_signal_6501, new_AGEMA_signal_6497, new_AGEMA_signal_6493}), .b ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, n2279}), .clk ( clk ), .r ({Fresh[1841], Fresh[1840], Fresh[1839]}), .c ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, n2280}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2451 ( .a ({new_AGEMA_signal_6759, new_AGEMA_signal_6757, new_AGEMA_signal_6755}), .b ({new_AGEMA_signal_1835, new_AGEMA_signal_1834, n2283}), .clk ( clk ), .r ({Fresh[1844], Fresh[1843], Fresh[1842]}), .c ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, n2286}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2461 ( .a ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, n2686}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, n2289}), .clk ( clk ), .r ({Fresh[1847], Fresh[1846], Fresh[1845]}), .c ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, n2304}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2466 ( .a ({new_AGEMA_signal_6765, new_AGEMA_signal_6763, new_AGEMA_signal_6761}), .b ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, n2292}), .clk ( clk ), .r ({Fresh[1850], Fresh[1849], Fresh[1848]}), .c ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, n2295}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2488 ( .a ({new_AGEMA_signal_2127, new_AGEMA_signal_2126, n2321}), .b ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, n2320}), .clk ( clk ), .r ({Fresh[1853], Fresh[1852], Fresh[1851]}), .c ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, n2322}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2499 ( .a ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, n2332}), .b ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, n2331}), .clk ( clk ), .r ({Fresh[1856], Fresh[1855], Fresh[1854]}), .c ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, n2333}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2509 ( .a ({new_AGEMA_signal_6777, new_AGEMA_signal_6773, new_AGEMA_signal_6769}), .b ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, n2342}), .clk ( clk ), .r ({Fresh[1859], Fresh[1858], Fresh[1857]}), .c ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, n2345}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2526 ( .a ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, n2358}), .b ({new_AGEMA_signal_6783, new_AGEMA_signal_6781, new_AGEMA_signal_6779}), .clk ( clk ), .r ({Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, n2361}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2549 ( .a ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, n2387}), .b ({new_AGEMA_signal_6789, new_AGEMA_signal_6787, new_AGEMA_signal_6785}), .clk ( clk ), .r ({Fresh[1865], Fresh[1864], Fresh[1863]}), .c ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, n2388}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2556 ( .a ({new_AGEMA_signal_6801, new_AGEMA_signal_6797, new_AGEMA_signal_6793}), .b ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, n2392}), .clk ( clk ), .r ({Fresh[1868], Fresh[1867], Fresh[1866]}), .c ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, n2393}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2567 ( .a ({new_AGEMA_signal_6813, new_AGEMA_signal_6809, new_AGEMA_signal_6805}), .b ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, n2404}), .clk ( clk ), .r ({Fresh[1871], Fresh[1870], Fresh[1869]}), .c ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, n2405}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2571 ( .a ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, n2409}), .b ({new_AGEMA_signal_6825, new_AGEMA_signal_6821, new_AGEMA_signal_6817}), .clk ( clk ), .r ({Fresh[1874], Fresh[1873], Fresh[1872]}), .c ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, n2410}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2576 ( .a ({new_AGEMA_signal_6837, new_AGEMA_signal_6833, new_AGEMA_signal_6829}), .b ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, n2414}), .clk ( clk ), .r ({Fresh[1877], Fresh[1876], Fresh[1875]}), .c ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, n2421}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2579 ( .a ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, n2418}), .b ({new_AGEMA_signal_6849, new_AGEMA_signal_6845, new_AGEMA_signal_6841}), .clk ( clk ), .r ({Fresh[1880], Fresh[1879], Fresh[1878]}), .c ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, n2419}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2590 ( .a ({new_AGEMA_signal_6855, new_AGEMA_signal_6853, new_AGEMA_signal_6851}), .b ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, n2432}), .clk ( clk ), .r ({Fresh[1883], Fresh[1882], Fresh[1881]}), .c ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, n2436}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2604 ( .a ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, n2449}), .b ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, n2448}), .clk ( clk ), .r ({Fresh[1886], Fresh[1885], Fresh[1884]}), .c ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, n2450}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2610 ( .a ({new_AGEMA_signal_6861, new_AGEMA_signal_6859, new_AGEMA_signal_6857}), .b ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, n2455}), .clk ( clk ), .r ({Fresh[1889], Fresh[1888], Fresh[1887]}), .c ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, n2456}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2613 ( .a ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, n2460}), .b ({new_AGEMA_signal_6867, new_AGEMA_signal_6865, new_AGEMA_signal_6863}), .clk ( clk ), .r ({Fresh[1892], Fresh[1891], Fresh[1890]}), .c ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, n2461}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2619 ( .a ({new_AGEMA_signal_6873, new_AGEMA_signal_6871, new_AGEMA_signal_6869}), .b ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, n2466}), .clk ( clk ), .r ({Fresh[1895], Fresh[1894], Fresh[1893]}), .c ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, n2469}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2630 ( .a ({new_AGEMA_signal_6885, new_AGEMA_signal_6881, new_AGEMA_signal_6877}), .b ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, n2477}), .clk ( clk ), .r ({Fresh[1898], Fresh[1897], Fresh[1896]}), .c ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, n2478}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2635 ( .a ({new_AGEMA_signal_6897, new_AGEMA_signal_6893, new_AGEMA_signal_6889}), .b ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, n2482}), .clk ( clk ), .r ({Fresh[1901], Fresh[1900], Fresh[1899]}), .c ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, n2484}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2643 ( .a ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, n2490}), .b ({new_AGEMA_signal_6903, new_AGEMA_signal_6901, new_AGEMA_signal_6899}), .clk ( clk ), .r ({Fresh[1904], Fresh[1903], Fresh[1902]}), .c ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, n2491}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2649 ( .a ({new_AGEMA_signal_6909, new_AGEMA_signal_6907, new_AGEMA_signal_6905}), .b ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, n2496}), .clk ( clk ), .r ({Fresh[1907], Fresh[1906], Fresh[1905]}), .c ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, n2500}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2656 ( .a ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, n2507}), .b ({new_AGEMA_signal_6915, new_AGEMA_signal_6913, new_AGEMA_signal_6911}), .clk ( clk ), .r ({Fresh[1910], Fresh[1909], Fresh[1908]}), .c ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, n2508}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2670 ( .a ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, n2525}), .b ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, n2524}), .clk ( clk ), .r ({Fresh[1913], Fresh[1912], Fresh[1911]}), .c ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, n2526}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2679 ( .a ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, n2537}), .b ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, n2536}), .clk ( clk ), .r ({Fresh[1916], Fresh[1915], Fresh[1914]}), .c ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, n2539}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2682 ( .a ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, n2543}), .b ({new_AGEMA_signal_6921, new_AGEMA_signal_6919, new_AGEMA_signal_6917}), .clk ( clk ), .r ({Fresh[1919], Fresh[1918], Fresh[1917]}), .c ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, n2548}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2694 ( .a ({new_AGEMA_signal_6927, new_AGEMA_signal_6925, new_AGEMA_signal_6923}), .b ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, n2557}), .clk ( clk ), .r ({Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, n2568}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2700 ( .a ({new_AGEMA_signal_6933, new_AGEMA_signal_6931, new_AGEMA_signal_6929}), .b ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, n2565}), .clk ( clk ), .r ({Fresh[1925], Fresh[1924], Fresh[1923]}), .c ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, n2567}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2710 ( .a ({new_AGEMA_signal_6939, new_AGEMA_signal_6937, new_AGEMA_signal_6935}), .b ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, n2580}), .clk ( clk ), .r ({Fresh[1928], Fresh[1927], Fresh[1926]}), .c ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, n2583}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2728 ( .a ({new_AGEMA_signal_6945, new_AGEMA_signal_6943, new_AGEMA_signal_6941}), .b ({new_AGEMA_signal_1623, new_AGEMA_signal_1622, n2602}), .clk ( clk ), .r ({Fresh[1931], Fresh[1930], Fresh[1929]}), .c ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, n2604}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2739 ( .a ({new_AGEMA_signal_6951, new_AGEMA_signal_6949, new_AGEMA_signal_6947}), .b ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, n2619}), .clk ( clk ), .r ({Fresh[1934], Fresh[1933], Fresh[1932]}), .c ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, n2621}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2745 ( .a ({new_AGEMA_signal_6963, new_AGEMA_signal_6959, new_AGEMA_signal_6955}), .b ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, n2628}), .clk ( clk ), .r ({Fresh[1937], Fresh[1936], Fresh[1935]}), .c ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, n2633}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2756 ( .a ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, n2649}), .b ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, n2648}), .clk ( clk ), .r ({Fresh[1940], Fresh[1939], Fresh[1938]}), .c ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, n2660}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2759 ( .a ({new_AGEMA_signal_6969, new_AGEMA_signal_6967, new_AGEMA_signal_6965}), .b ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, n2652}), .clk ( clk ), .r ({Fresh[1943], Fresh[1942], Fresh[1941]}), .c ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, n2656}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2766 ( .a ({new_AGEMA_signal_6975, new_AGEMA_signal_6973, new_AGEMA_signal_6971}), .b ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, n2664}), .clk ( clk ), .r ({Fresh[1946], Fresh[1945], Fresh[1944]}), .c ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, n2666}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2774 ( .a ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, n2681}), .b ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, n2680}), .clk ( clk ), .r ({Fresh[1949], Fresh[1948], Fresh[1947]}), .c ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, n2706}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2777 ( .a ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, n2686}), .b ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, n2685}), .clk ( clk ), .r ({Fresh[1952], Fresh[1951], Fresh[1950]}), .c ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, n2704}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2781 ( .a ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, n2692}), .b ({new_AGEMA_signal_6981, new_AGEMA_signal_6979, new_AGEMA_signal_6977}), .clk ( clk ), .r ({Fresh[1955], Fresh[1954], Fresh[1953]}), .c ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, n2696}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2794 ( .a ({new_AGEMA_signal_6987, new_AGEMA_signal_6985, new_AGEMA_signal_6983}), .b ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, n2716}), .clk ( clk ), .r ({Fresh[1958], Fresh[1957], Fresh[1956]}), .c ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, n2718}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2801 ( .a ({new_AGEMA_signal_6993, new_AGEMA_signal_6991, new_AGEMA_signal_6989}), .b ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, n2728}), .clk ( clk ), .r ({Fresh[1961], Fresh[1960], Fresh[1959]}), .c ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, n2730}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2805 ( .a ({new_AGEMA_signal_7005, new_AGEMA_signal_7001, new_AGEMA_signal_6997}), .b ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, n2735}), .clk ( clk ), .r ({Fresh[1964], Fresh[1963], Fresh[1962]}), .c ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, n2745}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2809 ( .a ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, n2743}), .b ({new_AGEMA_signal_7017, new_AGEMA_signal_7013, new_AGEMA_signal_7009}), .clk ( clk ), .r ({Fresh[1967], Fresh[1966], Fresh[1965]}), .c ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, n2744}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2814 ( .a ({new_AGEMA_signal_6753, new_AGEMA_signal_6751, new_AGEMA_signal_6749}), .b ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, n2751}), .clk ( clk ), .r ({Fresh[1970], Fresh[1969], Fresh[1968]}), .c ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, n2759}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2821 ( .a ({new_AGEMA_signal_7029, new_AGEMA_signal_7025, new_AGEMA_signal_7021}), .b ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, n2764}), .clk ( clk ), .r ({Fresh[1973], Fresh[1972], Fresh[1971]}), .c ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, n2771}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2833 ( .a ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, n2788}), .b ({new_AGEMA_signal_7041, new_AGEMA_signal_7037, new_AGEMA_signal_7033}), .clk ( clk ), .r ({Fresh[1976], Fresh[1975], Fresh[1974]}), .c ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, n2798}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2850 ( .a ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, n2822}), .b ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, n2821}), .clk ( clk ), .r ({Fresh[1979], Fresh[1978], Fresh[1977]}), .c ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, n2826}) ) ;
    buf_clk new_AGEMA_reg_buffer_2556 ( .C ( clk ), .D ( new_AGEMA_signal_7044 ), .Q ( new_AGEMA_signal_7045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2560 ( .C ( clk ), .D ( new_AGEMA_signal_7048 ), .Q ( new_AGEMA_signal_7049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2564 ( .C ( clk ), .D ( new_AGEMA_signal_7052 ), .Q ( new_AGEMA_signal_7053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2568 ( .C ( clk ), .D ( new_AGEMA_signal_7056 ), .Q ( new_AGEMA_signal_7057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2572 ( .C ( clk ), .D ( new_AGEMA_signal_7060 ), .Q ( new_AGEMA_signal_7061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2576 ( .C ( clk ), .D ( new_AGEMA_signal_7064 ), .Q ( new_AGEMA_signal_7065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2584 ( .C ( clk ), .D ( new_AGEMA_signal_7072 ), .Q ( new_AGEMA_signal_7073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2592 ( .C ( clk ), .D ( new_AGEMA_signal_7080 ), .Q ( new_AGEMA_signal_7081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2600 ( .C ( clk ), .D ( new_AGEMA_signal_7088 ), .Q ( new_AGEMA_signal_7089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2602 ( .C ( clk ), .D ( new_AGEMA_signal_7090 ), .Q ( new_AGEMA_signal_7091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2604 ( .C ( clk ), .D ( new_AGEMA_signal_7092 ), .Q ( new_AGEMA_signal_7093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2606 ( .C ( clk ), .D ( new_AGEMA_signal_7094 ), .Q ( new_AGEMA_signal_7095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2614 ( .C ( clk ), .D ( new_AGEMA_signal_7102 ), .Q ( new_AGEMA_signal_7103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2622 ( .C ( clk ), .D ( new_AGEMA_signal_7110 ), .Q ( new_AGEMA_signal_7111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2630 ( .C ( clk ), .D ( new_AGEMA_signal_7118 ), .Q ( new_AGEMA_signal_7119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2636 ( .C ( clk ), .D ( new_AGEMA_signal_7124 ), .Q ( new_AGEMA_signal_7125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2642 ( .C ( clk ), .D ( new_AGEMA_signal_7130 ), .Q ( new_AGEMA_signal_7131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2648 ( .C ( clk ), .D ( new_AGEMA_signal_7136 ), .Q ( new_AGEMA_signal_7137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2652 ( .C ( clk ), .D ( new_AGEMA_signal_7140 ), .Q ( new_AGEMA_signal_7141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2656 ( .C ( clk ), .D ( new_AGEMA_signal_7144 ), .Q ( new_AGEMA_signal_7145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2660 ( .C ( clk ), .D ( new_AGEMA_signal_7148 ), .Q ( new_AGEMA_signal_7149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2666 ( .C ( clk ), .D ( new_AGEMA_signal_7154 ), .Q ( new_AGEMA_signal_7155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2672 ( .C ( clk ), .D ( new_AGEMA_signal_7160 ), .Q ( new_AGEMA_signal_7161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2678 ( .C ( clk ), .D ( new_AGEMA_signal_7166 ), .Q ( new_AGEMA_signal_7167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2680 ( .C ( clk ), .D ( new_AGEMA_signal_7168 ), .Q ( new_AGEMA_signal_7169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2682 ( .C ( clk ), .D ( new_AGEMA_signal_7170 ), .Q ( new_AGEMA_signal_7171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2684 ( .C ( clk ), .D ( new_AGEMA_signal_7172 ), .Q ( new_AGEMA_signal_7173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2690 ( .C ( clk ), .D ( new_AGEMA_signal_7178 ), .Q ( new_AGEMA_signal_7179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2696 ( .C ( clk ), .D ( new_AGEMA_signal_7184 ), .Q ( new_AGEMA_signal_7185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2702 ( .C ( clk ), .D ( new_AGEMA_signal_7190 ), .Q ( new_AGEMA_signal_7191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2708 ( .C ( clk ), .D ( new_AGEMA_signal_7196 ), .Q ( new_AGEMA_signal_7197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2714 ( .C ( clk ), .D ( new_AGEMA_signal_7202 ), .Q ( new_AGEMA_signal_7203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2720 ( .C ( clk ), .D ( new_AGEMA_signal_7208 ), .Q ( new_AGEMA_signal_7209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2722 ( .C ( clk ), .D ( new_AGEMA_signal_7210 ), .Q ( new_AGEMA_signal_7211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2724 ( .C ( clk ), .D ( new_AGEMA_signal_7212 ), .Q ( new_AGEMA_signal_7213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2726 ( .C ( clk ), .D ( new_AGEMA_signal_7214 ), .Q ( new_AGEMA_signal_7215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2730 ( .C ( clk ), .D ( new_AGEMA_signal_7218 ), .Q ( new_AGEMA_signal_7219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2734 ( .C ( clk ), .D ( new_AGEMA_signal_7222 ), .Q ( new_AGEMA_signal_7223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2738 ( .C ( clk ), .D ( new_AGEMA_signal_7226 ), .Q ( new_AGEMA_signal_7227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2744 ( .C ( clk ), .D ( new_AGEMA_signal_7232 ), .Q ( new_AGEMA_signal_7233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2750 ( .C ( clk ), .D ( new_AGEMA_signal_7238 ), .Q ( new_AGEMA_signal_7239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2756 ( .C ( clk ), .D ( new_AGEMA_signal_7244 ), .Q ( new_AGEMA_signal_7245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2762 ( .C ( clk ), .D ( new_AGEMA_signal_7250 ), .Q ( new_AGEMA_signal_7251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2768 ( .C ( clk ), .D ( new_AGEMA_signal_7256 ), .Q ( new_AGEMA_signal_7257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2774 ( .C ( clk ), .D ( new_AGEMA_signal_7262 ), .Q ( new_AGEMA_signal_7263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2776 ( .C ( clk ), .D ( new_AGEMA_signal_7264 ), .Q ( new_AGEMA_signal_7265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2778 ( .C ( clk ), .D ( new_AGEMA_signal_7266 ), .Q ( new_AGEMA_signal_7267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2780 ( .C ( clk ), .D ( new_AGEMA_signal_7268 ), .Q ( new_AGEMA_signal_7269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2786 ( .C ( clk ), .D ( new_AGEMA_signal_7274 ), .Q ( new_AGEMA_signal_7275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2792 ( .C ( clk ), .D ( new_AGEMA_signal_7280 ), .Q ( new_AGEMA_signal_7281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2798 ( .C ( clk ), .D ( new_AGEMA_signal_7286 ), .Q ( new_AGEMA_signal_7287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2800 ( .C ( clk ), .D ( new_AGEMA_signal_7288 ), .Q ( new_AGEMA_signal_7289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2802 ( .C ( clk ), .D ( new_AGEMA_signal_7290 ), .Q ( new_AGEMA_signal_7291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2804 ( .C ( clk ), .D ( new_AGEMA_signal_7292 ), .Q ( new_AGEMA_signal_7293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2808 ( .C ( clk ), .D ( new_AGEMA_signal_7296 ), .Q ( new_AGEMA_signal_7297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2812 ( .C ( clk ), .D ( new_AGEMA_signal_7300 ), .Q ( new_AGEMA_signal_7301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2816 ( .C ( clk ), .D ( new_AGEMA_signal_7304 ), .Q ( new_AGEMA_signal_7305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2820 ( .C ( clk ), .D ( new_AGEMA_signal_7308 ), .Q ( new_AGEMA_signal_7309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2824 ( .C ( clk ), .D ( new_AGEMA_signal_7312 ), .Q ( new_AGEMA_signal_7313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2828 ( .C ( clk ), .D ( new_AGEMA_signal_7316 ), .Q ( new_AGEMA_signal_7317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2830 ( .C ( clk ), .D ( new_AGEMA_signal_7318 ), .Q ( new_AGEMA_signal_7319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2832 ( .C ( clk ), .D ( new_AGEMA_signal_7320 ), .Q ( new_AGEMA_signal_7321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2834 ( .C ( clk ), .D ( new_AGEMA_signal_7322 ), .Q ( new_AGEMA_signal_7323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2842 ( .C ( clk ), .D ( new_AGEMA_signal_7330 ), .Q ( new_AGEMA_signal_7331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2850 ( .C ( clk ), .D ( new_AGEMA_signal_7338 ), .Q ( new_AGEMA_signal_7339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2858 ( .C ( clk ), .D ( new_AGEMA_signal_7346 ), .Q ( new_AGEMA_signal_7347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2864 ( .C ( clk ), .D ( new_AGEMA_signal_7352 ), .Q ( new_AGEMA_signal_7353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2870 ( .C ( clk ), .D ( new_AGEMA_signal_7358 ), .Q ( new_AGEMA_signal_7359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2876 ( .C ( clk ), .D ( new_AGEMA_signal_7364 ), .Q ( new_AGEMA_signal_7365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2880 ( .C ( clk ), .D ( new_AGEMA_signal_7368 ), .Q ( new_AGEMA_signal_7369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2884 ( .C ( clk ), .D ( new_AGEMA_signal_7372 ), .Q ( new_AGEMA_signal_7373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2888 ( .C ( clk ), .D ( new_AGEMA_signal_7376 ), .Q ( new_AGEMA_signal_7377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2892 ( .C ( clk ), .D ( new_AGEMA_signal_7380 ), .Q ( new_AGEMA_signal_7381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2896 ( .C ( clk ), .D ( new_AGEMA_signal_7384 ), .Q ( new_AGEMA_signal_7385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2900 ( .C ( clk ), .D ( new_AGEMA_signal_7388 ), .Q ( new_AGEMA_signal_7389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2902 ( .C ( clk ), .D ( new_AGEMA_signal_7390 ), .Q ( new_AGEMA_signal_7391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2904 ( .C ( clk ), .D ( new_AGEMA_signal_7392 ), .Q ( new_AGEMA_signal_7393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2906 ( .C ( clk ), .D ( new_AGEMA_signal_7394 ), .Q ( new_AGEMA_signal_7395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2908 ( .C ( clk ), .D ( new_AGEMA_signal_7396 ), .Q ( new_AGEMA_signal_7397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2910 ( .C ( clk ), .D ( new_AGEMA_signal_7398 ), .Q ( new_AGEMA_signal_7399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2912 ( .C ( clk ), .D ( new_AGEMA_signal_7400 ), .Q ( new_AGEMA_signal_7401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2916 ( .C ( clk ), .D ( new_AGEMA_signal_7404 ), .Q ( new_AGEMA_signal_7405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2920 ( .C ( clk ), .D ( new_AGEMA_signal_7408 ), .Q ( new_AGEMA_signal_7409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2924 ( .C ( clk ), .D ( new_AGEMA_signal_7412 ), .Q ( new_AGEMA_signal_7413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2928 ( .C ( clk ), .D ( new_AGEMA_signal_7416 ), .Q ( new_AGEMA_signal_7417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2932 ( .C ( clk ), .D ( new_AGEMA_signal_7420 ), .Q ( new_AGEMA_signal_7421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2936 ( .C ( clk ), .D ( new_AGEMA_signal_7424 ), .Q ( new_AGEMA_signal_7425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2938 ( .C ( clk ), .D ( new_AGEMA_signal_7426 ), .Q ( new_AGEMA_signal_7427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2940 ( .C ( clk ), .D ( new_AGEMA_signal_7428 ), .Q ( new_AGEMA_signal_7429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2942 ( .C ( clk ), .D ( new_AGEMA_signal_7430 ), .Q ( new_AGEMA_signal_7431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2948 ( .C ( clk ), .D ( new_AGEMA_signal_7436 ), .Q ( new_AGEMA_signal_7437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2954 ( .C ( clk ), .D ( new_AGEMA_signal_7442 ), .Q ( new_AGEMA_signal_7443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2960 ( .C ( clk ), .D ( new_AGEMA_signal_7448 ), .Q ( new_AGEMA_signal_7449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2964 ( .C ( clk ), .D ( new_AGEMA_signal_7452 ), .Q ( new_AGEMA_signal_7453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2968 ( .C ( clk ), .D ( new_AGEMA_signal_7456 ), .Q ( new_AGEMA_signal_7457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2972 ( .C ( clk ), .D ( new_AGEMA_signal_7460 ), .Q ( new_AGEMA_signal_7461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2974 ( .C ( clk ), .D ( new_AGEMA_signal_7462 ), .Q ( new_AGEMA_signal_7463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2976 ( .C ( clk ), .D ( new_AGEMA_signal_7464 ), .Q ( new_AGEMA_signal_7465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2978 ( .C ( clk ), .D ( new_AGEMA_signal_7466 ), .Q ( new_AGEMA_signal_7467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2982 ( .C ( clk ), .D ( new_AGEMA_signal_7470 ), .Q ( new_AGEMA_signal_7471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2986 ( .C ( clk ), .D ( new_AGEMA_signal_7474 ), .Q ( new_AGEMA_signal_7475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2990 ( .C ( clk ), .D ( new_AGEMA_signal_7478 ), .Q ( new_AGEMA_signal_7479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2994 ( .C ( clk ), .D ( new_AGEMA_signal_7482 ), .Q ( new_AGEMA_signal_7483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2998 ( .C ( clk ), .D ( new_AGEMA_signal_7486 ), .Q ( new_AGEMA_signal_7487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3002 ( .C ( clk ), .D ( new_AGEMA_signal_7490 ), .Q ( new_AGEMA_signal_7491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3006 ( .C ( clk ), .D ( new_AGEMA_signal_7494 ), .Q ( new_AGEMA_signal_7495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3010 ( .C ( clk ), .D ( new_AGEMA_signal_7498 ), .Q ( new_AGEMA_signal_7499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3014 ( .C ( clk ), .D ( new_AGEMA_signal_7502 ), .Q ( new_AGEMA_signal_7503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3016 ( .C ( clk ), .D ( new_AGEMA_signal_7504 ), .Q ( new_AGEMA_signal_7505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3018 ( .C ( clk ), .D ( new_AGEMA_signal_7506 ), .Q ( new_AGEMA_signal_7507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3020 ( .C ( clk ), .D ( new_AGEMA_signal_7508 ), .Q ( new_AGEMA_signal_7509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3024 ( .C ( clk ), .D ( new_AGEMA_signal_7512 ), .Q ( new_AGEMA_signal_7513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3028 ( .C ( clk ), .D ( new_AGEMA_signal_7516 ), .Q ( new_AGEMA_signal_7517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3032 ( .C ( clk ), .D ( new_AGEMA_signal_7520 ), .Q ( new_AGEMA_signal_7521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3034 ( .C ( clk ), .D ( new_AGEMA_signal_7522 ), .Q ( new_AGEMA_signal_7523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3036 ( .C ( clk ), .D ( new_AGEMA_signal_7524 ), .Q ( new_AGEMA_signal_7525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3038 ( .C ( clk ), .D ( new_AGEMA_signal_7526 ), .Q ( new_AGEMA_signal_7527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3044 ( .C ( clk ), .D ( new_AGEMA_signal_7532 ), .Q ( new_AGEMA_signal_7533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3050 ( .C ( clk ), .D ( new_AGEMA_signal_7538 ), .Q ( new_AGEMA_signal_7539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3056 ( .C ( clk ), .D ( new_AGEMA_signal_7544 ), .Q ( new_AGEMA_signal_7545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3062 ( .C ( clk ), .D ( new_AGEMA_signal_7550 ), .Q ( new_AGEMA_signal_7551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3068 ( .C ( clk ), .D ( new_AGEMA_signal_7556 ), .Q ( new_AGEMA_signal_7557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3074 ( .C ( clk ), .D ( new_AGEMA_signal_7562 ), .Q ( new_AGEMA_signal_7563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3078 ( .C ( clk ), .D ( new_AGEMA_signal_7566 ), .Q ( new_AGEMA_signal_7567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3082 ( .C ( clk ), .D ( new_AGEMA_signal_7570 ), .Q ( new_AGEMA_signal_7571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3086 ( .C ( clk ), .D ( new_AGEMA_signal_7574 ), .Q ( new_AGEMA_signal_7575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3088 ( .C ( clk ), .D ( new_AGEMA_signal_7576 ), .Q ( new_AGEMA_signal_7577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3090 ( .C ( clk ), .D ( new_AGEMA_signal_7578 ), .Q ( new_AGEMA_signal_7579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3092 ( .C ( clk ), .D ( new_AGEMA_signal_7580 ), .Q ( new_AGEMA_signal_7581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3100 ( .C ( clk ), .D ( new_AGEMA_signal_7588 ), .Q ( new_AGEMA_signal_7589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3108 ( .C ( clk ), .D ( new_AGEMA_signal_7596 ), .Q ( new_AGEMA_signal_7597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3116 ( .C ( clk ), .D ( new_AGEMA_signal_7604 ), .Q ( new_AGEMA_signal_7605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3118 ( .C ( clk ), .D ( new_AGEMA_signal_7606 ), .Q ( new_AGEMA_signal_7607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3120 ( .C ( clk ), .D ( new_AGEMA_signal_7608 ), .Q ( new_AGEMA_signal_7609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3122 ( .C ( clk ), .D ( new_AGEMA_signal_7610 ), .Q ( new_AGEMA_signal_7611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3126 ( .C ( clk ), .D ( new_AGEMA_signal_7614 ), .Q ( new_AGEMA_signal_7615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3130 ( .C ( clk ), .D ( new_AGEMA_signal_7618 ), .Q ( new_AGEMA_signal_7619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3134 ( .C ( clk ), .D ( new_AGEMA_signal_7622 ), .Q ( new_AGEMA_signal_7623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3138 ( .C ( clk ), .D ( new_AGEMA_signal_7626 ), .Q ( new_AGEMA_signal_7627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3142 ( .C ( clk ), .D ( new_AGEMA_signal_7630 ), .Q ( new_AGEMA_signal_7631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3146 ( .C ( clk ), .D ( new_AGEMA_signal_7634 ), .Q ( new_AGEMA_signal_7635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3150 ( .C ( clk ), .D ( new_AGEMA_signal_7638 ), .Q ( new_AGEMA_signal_7639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3154 ( .C ( clk ), .D ( new_AGEMA_signal_7642 ), .Q ( new_AGEMA_signal_7643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3158 ( .C ( clk ), .D ( new_AGEMA_signal_7646 ), .Q ( new_AGEMA_signal_7647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3162 ( .C ( clk ), .D ( new_AGEMA_signal_7650 ), .Q ( new_AGEMA_signal_7651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3166 ( .C ( clk ), .D ( new_AGEMA_signal_7654 ), .Q ( new_AGEMA_signal_7655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3170 ( .C ( clk ), .D ( new_AGEMA_signal_7658 ), .Q ( new_AGEMA_signal_7659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3174 ( .C ( clk ), .D ( new_AGEMA_signal_7662 ), .Q ( new_AGEMA_signal_7663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3178 ( .C ( clk ), .D ( new_AGEMA_signal_7666 ), .Q ( new_AGEMA_signal_7667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3182 ( .C ( clk ), .D ( new_AGEMA_signal_7670 ), .Q ( new_AGEMA_signal_7671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3190 ( .C ( clk ), .D ( new_AGEMA_signal_7678 ), .Q ( new_AGEMA_signal_7679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3198 ( .C ( clk ), .D ( new_AGEMA_signal_7686 ), .Q ( new_AGEMA_signal_7687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3206 ( .C ( clk ), .D ( new_AGEMA_signal_7694 ), .Q ( new_AGEMA_signal_7695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3208 ( .C ( clk ), .D ( new_AGEMA_signal_7696 ), .Q ( new_AGEMA_signal_7697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3210 ( .C ( clk ), .D ( new_AGEMA_signal_7698 ), .Q ( new_AGEMA_signal_7699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3212 ( .C ( clk ), .D ( new_AGEMA_signal_7700 ), .Q ( new_AGEMA_signal_7701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3216 ( .C ( clk ), .D ( new_AGEMA_signal_7704 ), .Q ( new_AGEMA_signal_7705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3220 ( .C ( clk ), .D ( new_AGEMA_signal_7708 ), .Q ( new_AGEMA_signal_7709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3224 ( .C ( clk ), .D ( new_AGEMA_signal_7712 ), .Q ( new_AGEMA_signal_7713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3226 ( .C ( clk ), .D ( new_AGEMA_signal_7714 ), .Q ( new_AGEMA_signal_7715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3228 ( .C ( clk ), .D ( new_AGEMA_signal_7716 ), .Q ( new_AGEMA_signal_7717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3230 ( .C ( clk ), .D ( new_AGEMA_signal_7718 ), .Q ( new_AGEMA_signal_7719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3236 ( .C ( clk ), .D ( new_AGEMA_signal_7724 ), .Q ( new_AGEMA_signal_7725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3242 ( .C ( clk ), .D ( new_AGEMA_signal_7730 ), .Q ( new_AGEMA_signal_7731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3248 ( .C ( clk ), .D ( new_AGEMA_signal_7736 ), .Q ( new_AGEMA_signal_7737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3260 ( .C ( clk ), .D ( new_AGEMA_signal_7748 ), .Q ( new_AGEMA_signal_7749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3268 ( .C ( clk ), .D ( new_AGEMA_signal_7756 ), .Q ( new_AGEMA_signal_7757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3276 ( .C ( clk ), .D ( new_AGEMA_signal_7764 ), .Q ( new_AGEMA_signal_7765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3286 ( .C ( clk ), .D ( new_AGEMA_signal_7774 ), .Q ( new_AGEMA_signal_7775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3290 ( .C ( clk ), .D ( new_AGEMA_signal_7778 ), .Q ( new_AGEMA_signal_7779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3294 ( .C ( clk ), .D ( new_AGEMA_signal_7782 ), .Q ( new_AGEMA_signal_7783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3302 ( .C ( clk ), .D ( new_AGEMA_signal_7790 ), .Q ( new_AGEMA_signal_7791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3310 ( .C ( clk ), .D ( new_AGEMA_signal_7798 ), .Q ( new_AGEMA_signal_7799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3318 ( .C ( clk ), .D ( new_AGEMA_signal_7806 ), .Q ( new_AGEMA_signal_7807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3330 ( .C ( clk ), .D ( new_AGEMA_signal_7818 ), .Q ( new_AGEMA_signal_7819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3336 ( .C ( clk ), .D ( new_AGEMA_signal_7824 ), .Q ( new_AGEMA_signal_7825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3342 ( .C ( clk ), .D ( new_AGEMA_signal_7830 ), .Q ( new_AGEMA_signal_7831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3346 ( .C ( clk ), .D ( new_AGEMA_signal_7834 ), .Q ( new_AGEMA_signal_7835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3350 ( .C ( clk ), .D ( new_AGEMA_signal_7838 ), .Q ( new_AGEMA_signal_7839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3354 ( .C ( clk ), .D ( new_AGEMA_signal_7842 ), .Q ( new_AGEMA_signal_7843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3362 ( .C ( clk ), .D ( new_AGEMA_signal_7850 ), .Q ( new_AGEMA_signal_7851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3370 ( .C ( clk ), .D ( new_AGEMA_signal_7858 ), .Q ( new_AGEMA_signal_7859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3378 ( .C ( clk ), .D ( new_AGEMA_signal_7866 ), .Q ( new_AGEMA_signal_7867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3382 ( .C ( clk ), .D ( new_AGEMA_signal_7870 ), .Q ( new_AGEMA_signal_7871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3386 ( .C ( clk ), .D ( new_AGEMA_signal_7874 ), .Q ( new_AGEMA_signal_7875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3390 ( .C ( clk ), .D ( new_AGEMA_signal_7878 ), .Q ( new_AGEMA_signal_7879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3396 ( .C ( clk ), .D ( new_AGEMA_signal_7884 ), .Q ( new_AGEMA_signal_7885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3402 ( .C ( clk ), .D ( new_AGEMA_signal_7890 ), .Q ( new_AGEMA_signal_7891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3408 ( .C ( clk ), .D ( new_AGEMA_signal_7896 ), .Q ( new_AGEMA_signal_7897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3414 ( .C ( clk ), .D ( new_AGEMA_signal_7902 ), .Q ( new_AGEMA_signal_7903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3420 ( .C ( clk ), .D ( new_AGEMA_signal_7908 ), .Q ( new_AGEMA_signal_7909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3426 ( .C ( clk ), .D ( new_AGEMA_signal_7914 ), .Q ( new_AGEMA_signal_7915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3432 ( .C ( clk ), .D ( new_AGEMA_signal_7920 ), .Q ( new_AGEMA_signal_7921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3438 ( .C ( clk ), .D ( new_AGEMA_signal_7926 ), .Q ( new_AGEMA_signal_7927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3444 ( .C ( clk ), .D ( new_AGEMA_signal_7932 ), .Q ( new_AGEMA_signal_7933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3450 ( .C ( clk ), .D ( new_AGEMA_signal_7938 ), .Q ( new_AGEMA_signal_7939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3456 ( .C ( clk ), .D ( new_AGEMA_signal_7944 ), .Q ( new_AGEMA_signal_7945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3462 ( .C ( clk ), .D ( new_AGEMA_signal_7950 ), .Q ( new_AGEMA_signal_7951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3468 ( .C ( clk ), .D ( new_AGEMA_signal_7956 ), .Q ( new_AGEMA_signal_7957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3474 ( .C ( clk ), .D ( new_AGEMA_signal_7962 ), .Q ( new_AGEMA_signal_7963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3480 ( .C ( clk ), .D ( new_AGEMA_signal_7968 ), .Q ( new_AGEMA_signal_7969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3484 ( .C ( clk ), .D ( new_AGEMA_signal_7972 ), .Q ( new_AGEMA_signal_7973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3488 ( .C ( clk ), .D ( new_AGEMA_signal_7976 ), .Q ( new_AGEMA_signal_7977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3492 ( .C ( clk ), .D ( new_AGEMA_signal_7980 ), .Q ( new_AGEMA_signal_7981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3500 ( .C ( clk ), .D ( new_AGEMA_signal_7988 ), .Q ( new_AGEMA_signal_7989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3508 ( .C ( clk ), .D ( new_AGEMA_signal_7996 ), .Q ( new_AGEMA_signal_7997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3516 ( .C ( clk ), .D ( new_AGEMA_signal_8004 ), .Q ( new_AGEMA_signal_8005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3520 ( .C ( clk ), .D ( new_AGEMA_signal_8008 ), .Q ( new_AGEMA_signal_8009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3524 ( .C ( clk ), .D ( new_AGEMA_signal_8012 ), .Q ( new_AGEMA_signal_8013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3528 ( .C ( clk ), .D ( new_AGEMA_signal_8016 ), .Q ( new_AGEMA_signal_8017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3534 ( .C ( clk ), .D ( new_AGEMA_signal_8022 ), .Q ( new_AGEMA_signal_8023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3540 ( .C ( clk ), .D ( new_AGEMA_signal_8028 ), .Q ( new_AGEMA_signal_8029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3546 ( .C ( clk ), .D ( new_AGEMA_signal_8034 ), .Q ( new_AGEMA_signal_8035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3554 ( .C ( clk ), .D ( new_AGEMA_signal_8042 ), .Q ( new_AGEMA_signal_8043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3562 ( .C ( clk ), .D ( new_AGEMA_signal_8050 ), .Q ( new_AGEMA_signal_8051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3570 ( .C ( clk ), .D ( new_AGEMA_signal_8058 ), .Q ( new_AGEMA_signal_8059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3582 ( .C ( clk ), .D ( new_AGEMA_signal_8070 ), .Q ( new_AGEMA_signal_8071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3588 ( .C ( clk ), .D ( new_AGEMA_signal_8076 ), .Q ( new_AGEMA_signal_8077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3594 ( .C ( clk ), .D ( new_AGEMA_signal_8082 ), .Q ( new_AGEMA_signal_8083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3612 ( .C ( clk ), .D ( new_AGEMA_signal_8100 ), .Q ( new_AGEMA_signal_8101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3618 ( .C ( clk ), .D ( new_AGEMA_signal_8106 ), .Q ( new_AGEMA_signal_8107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3624 ( .C ( clk ), .D ( new_AGEMA_signal_8112 ), .Q ( new_AGEMA_signal_8113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3630 ( .C ( clk ), .D ( new_AGEMA_signal_8118 ), .Q ( new_AGEMA_signal_8119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3636 ( .C ( clk ), .D ( new_AGEMA_signal_8124 ), .Q ( new_AGEMA_signal_8125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3642 ( .C ( clk ), .D ( new_AGEMA_signal_8130 ), .Q ( new_AGEMA_signal_8131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3650 ( .C ( clk ), .D ( new_AGEMA_signal_8138 ), .Q ( new_AGEMA_signal_8139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3658 ( .C ( clk ), .D ( new_AGEMA_signal_8146 ), .Q ( new_AGEMA_signal_8147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3666 ( .C ( clk ), .D ( new_AGEMA_signal_8154 ), .Q ( new_AGEMA_signal_8155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3674 ( .C ( clk ), .D ( new_AGEMA_signal_8162 ), .Q ( new_AGEMA_signal_8163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3682 ( .C ( clk ), .D ( new_AGEMA_signal_8170 ), .Q ( new_AGEMA_signal_8171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3690 ( .C ( clk ), .D ( new_AGEMA_signal_8178 ), .Q ( new_AGEMA_signal_8179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3696 ( .C ( clk ), .D ( new_AGEMA_signal_8184 ), .Q ( new_AGEMA_signal_8185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3702 ( .C ( clk ), .D ( new_AGEMA_signal_8190 ), .Q ( new_AGEMA_signal_8191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3708 ( .C ( clk ), .D ( new_AGEMA_signal_8196 ), .Q ( new_AGEMA_signal_8197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3714 ( .C ( clk ), .D ( new_AGEMA_signal_8202 ), .Q ( new_AGEMA_signal_8203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3720 ( .C ( clk ), .D ( new_AGEMA_signal_8208 ), .Q ( new_AGEMA_signal_8209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3726 ( .C ( clk ), .D ( new_AGEMA_signal_8214 ), .Q ( new_AGEMA_signal_8215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3736 ( .C ( clk ), .D ( new_AGEMA_signal_8224 ), .Q ( new_AGEMA_signal_8225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3740 ( .C ( clk ), .D ( new_AGEMA_signal_8228 ), .Q ( new_AGEMA_signal_8229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3744 ( .C ( clk ), .D ( new_AGEMA_signal_8232 ), .Q ( new_AGEMA_signal_8233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3748 ( .C ( clk ), .D ( new_AGEMA_signal_8236 ), .Q ( new_AGEMA_signal_8237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3752 ( .C ( clk ), .D ( new_AGEMA_signal_8240 ), .Q ( new_AGEMA_signal_8241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3756 ( .C ( clk ), .D ( new_AGEMA_signal_8244 ), .Q ( new_AGEMA_signal_8245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3760 ( .C ( clk ), .D ( new_AGEMA_signal_8248 ), .Q ( new_AGEMA_signal_8249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3764 ( .C ( clk ), .D ( new_AGEMA_signal_8252 ), .Q ( new_AGEMA_signal_8253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3768 ( .C ( clk ), .D ( new_AGEMA_signal_8256 ), .Q ( new_AGEMA_signal_8257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3778 ( .C ( clk ), .D ( new_AGEMA_signal_8266 ), .Q ( new_AGEMA_signal_8267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3784 ( .C ( clk ), .D ( new_AGEMA_signal_8272 ), .Q ( new_AGEMA_signal_8273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3790 ( .C ( clk ), .D ( new_AGEMA_signal_8278 ), .Q ( new_AGEMA_signal_8279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3816 ( .C ( clk ), .D ( new_AGEMA_signal_8304 ), .Q ( new_AGEMA_signal_8305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3824 ( .C ( clk ), .D ( new_AGEMA_signal_8312 ), .Q ( new_AGEMA_signal_8313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3832 ( .C ( clk ), .D ( new_AGEMA_signal_8320 ), .Q ( new_AGEMA_signal_8321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3840 ( .C ( clk ), .D ( new_AGEMA_signal_8328 ), .Q ( new_AGEMA_signal_8329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3848 ( .C ( clk ), .D ( new_AGEMA_signal_8336 ), .Q ( new_AGEMA_signal_8337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3856 ( .C ( clk ), .D ( new_AGEMA_signal_8344 ), .Q ( new_AGEMA_signal_8345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3864 ( .C ( clk ), .D ( new_AGEMA_signal_8352 ), .Q ( new_AGEMA_signal_8353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3872 ( .C ( clk ), .D ( new_AGEMA_signal_8360 ), .Q ( new_AGEMA_signal_8361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3880 ( .C ( clk ), .D ( new_AGEMA_signal_8368 ), .Q ( new_AGEMA_signal_8369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3888 ( .C ( clk ), .D ( new_AGEMA_signal_8376 ), .Q ( new_AGEMA_signal_8377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3896 ( .C ( clk ), .D ( new_AGEMA_signal_8384 ), .Q ( new_AGEMA_signal_8385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3904 ( .C ( clk ), .D ( new_AGEMA_signal_8392 ), .Q ( new_AGEMA_signal_8393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3910 ( .C ( clk ), .D ( new_AGEMA_signal_8398 ), .Q ( new_AGEMA_signal_8399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3916 ( .C ( clk ), .D ( new_AGEMA_signal_8404 ), .Q ( new_AGEMA_signal_8405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3922 ( .C ( clk ), .D ( new_AGEMA_signal_8410 ), .Q ( new_AGEMA_signal_8411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3932 ( .C ( clk ), .D ( new_AGEMA_signal_8420 ), .Q ( new_AGEMA_signal_8421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3942 ( .C ( clk ), .D ( new_AGEMA_signal_8430 ), .Q ( new_AGEMA_signal_8431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3952 ( .C ( clk ), .D ( new_AGEMA_signal_8440 ), .Q ( new_AGEMA_signal_8441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3960 ( .C ( clk ), .D ( new_AGEMA_signal_8448 ), .Q ( new_AGEMA_signal_8449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3968 ( .C ( clk ), .D ( new_AGEMA_signal_8456 ), .Q ( new_AGEMA_signal_8457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3976 ( .C ( clk ), .D ( new_AGEMA_signal_8464 ), .Q ( new_AGEMA_signal_8465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3984 ( .C ( clk ), .D ( new_AGEMA_signal_8472 ), .Q ( new_AGEMA_signal_8473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3992 ( .C ( clk ), .D ( new_AGEMA_signal_8480 ), .Q ( new_AGEMA_signal_8481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4000 ( .C ( clk ), .D ( new_AGEMA_signal_8488 ), .Q ( new_AGEMA_signal_8489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4008 ( .C ( clk ), .D ( new_AGEMA_signal_8496 ), .Q ( new_AGEMA_signal_8497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4016 ( .C ( clk ), .D ( new_AGEMA_signal_8504 ), .Q ( new_AGEMA_signal_8505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4024 ( .C ( clk ), .D ( new_AGEMA_signal_8512 ), .Q ( new_AGEMA_signal_8513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4048 ( .C ( clk ), .D ( new_AGEMA_signal_8536 ), .Q ( new_AGEMA_signal_8537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4054 ( .C ( clk ), .D ( new_AGEMA_signal_8542 ), .Q ( new_AGEMA_signal_8543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4060 ( .C ( clk ), .D ( new_AGEMA_signal_8548 ), .Q ( new_AGEMA_signal_8549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4082 ( .C ( clk ), .D ( new_AGEMA_signal_8570 ), .Q ( new_AGEMA_signal_8571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4092 ( .C ( clk ), .D ( new_AGEMA_signal_8580 ), .Q ( new_AGEMA_signal_8581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4102 ( .C ( clk ), .D ( new_AGEMA_signal_8590 ), .Q ( new_AGEMA_signal_8591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4110 ( .C ( clk ), .D ( new_AGEMA_signal_8598 ), .Q ( new_AGEMA_signal_8599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4118 ( .C ( clk ), .D ( new_AGEMA_signal_8606 ), .Q ( new_AGEMA_signal_8607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4126 ( .C ( clk ), .D ( new_AGEMA_signal_8614 ), .Q ( new_AGEMA_signal_8615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4152 ( .C ( clk ), .D ( new_AGEMA_signal_8640 ), .Q ( new_AGEMA_signal_8641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4160 ( .C ( clk ), .D ( new_AGEMA_signal_8648 ), .Q ( new_AGEMA_signal_8649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4168 ( .C ( clk ), .D ( new_AGEMA_signal_8656 ), .Q ( new_AGEMA_signal_8657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4176 ( .C ( clk ), .D ( new_AGEMA_signal_8664 ), .Q ( new_AGEMA_signal_8665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4184 ( .C ( clk ), .D ( new_AGEMA_signal_8672 ), .Q ( new_AGEMA_signal_8673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4192 ( .C ( clk ), .D ( new_AGEMA_signal_8680 ), .Q ( new_AGEMA_signal_8681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4198 ( .C ( clk ), .D ( new_AGEMA_signal_8686 ), .Q ( new_AGEMA_signal_8687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4204 ( .C ( clk ), .D ( new_AGEMA_signal_8692 ), .Q ( new_AGEMA_signal_8693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4210 ( .C ( clk ), .D ( new_AGEMA_signal_8698 ), .Q ( new_AGEMA_signal_8699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4230 ( .C ( clk ), .D ( new_AGEMA_signal_8718 ), .Q ( new_AGEMA_signal_8719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4238 ( .C ( clk ), .D ( new_AGEMA_signal_8726 ), .Q ( new_AGEMA_signal_8727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4246 ( .C ( clk ), .D ( new_AGEMA_signal_8734 ), .Q ( new_AGEMA_signal_8735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4324 ( .C ( clk ), .D ( new_AGEMA_signal_8812 ), .Q ( new_AGEMA_signal_8813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4332 ( .C ( clk ), .D ( new_AGEMA_signal_8820 ), .Q ( new_AGEMA_signal_8821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4340 ( .C ( clk ), .D ( new_AGEMA_signal_8828 ), .Q ( new_AGEMA_signal_8829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4378 ( .C ( clk ), .D ( new_AGEMA_signal_8866 ), .Q ( new_AGEMA_signal_8867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4386 ( .C ( clk ), .D ( new_AGEMA_signal_8874 ), .Q ( new_AGEMA_signal_8875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4394 ( .C ( clk ), .D ( new_AGEMA_signal_8882 ), .Q ( new_AGEMA_signal_8883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4402 ( .C ( clk ), .D ( new_AGEMA_signal_8890 ), .Q ( new_AGEMA_signal_8891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4410 ( .C ( clk ), .D ( new_AGEMA_signal_8898 ), .Q ( new_AGEMA_signal_8899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4418 ( .C ( clk ), .D ( new_AGEMA_signal_8906 ), .Q ( new_AGEMA_signal_8907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4428 ( .C ( clk ), .D ( new_AGEMA_signal_8916 ), .Q ( new_AGEMA_signal_8917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4438 ( .C ( clk ), .D ( new_AGEMA_signal_8926 ), .Q ( new_AGEMA_signal_8927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4448 ( .C ( clk ), .D ( new_AGEMA_signal_8936 ), .Q ( new_AGEMA_signal_8937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4456 ( .C ( clk ), .D ( new_AGEMA_signal_8944 ), .Q ( new_AGEMA_signal_8945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4464 ( .C ( clk ), .D ( new_AGEMA_signal_8952 ), .Q ( new_AGEMA_signal_8953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4472 ( .C ( clk ), .D ( new_AGEMA_signal_8960 ), .Q ( new_AGEMA_signal_8961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4528 ( .C ( clk ), .D ( new_AGEMA_signal_9016 ), .Q ( new_AGEMA_signal_9017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4536 ( .C ( clk ), .D ( new_AGEMA_signal_9024 ), .Q ( new_AGEMA_signal_9025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4544 ( .C ( clk ), .D ( new_AGEMA_signal_9032 ), .Q ( new_AGEMA_signal_9033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4576 ( .C ( clk ), .D ( new_AGEMA_signal_9064 ), .Q ( new_AGEMA_signal_9065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4584 ( .C ( clk ), .D ( new_AGEMA_signal_9072 ), .Q ( new_AGEMA_signal_9073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4592 ( .C ( clk ), .D ( new_AGEMA_signal_9080 ), .Q ( new_AGEMA_signal_9081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4708 ( .C ( clk ), .D ( new_AGEMA_signal_9196 ), .Q ( new_AGEMA_signal_9197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4718 ( .C ( clk ), .D ( new_AGEMA_signal_9206 ), .Q ( new_AGEMA_signal_9207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4728 ( .C ( clk ), .D ( new_AGEMA_signal_9216 ), .Q ( new_AGEMA_signal_9217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4978 ( .C ( clk ), .D ( new_AGEMA_signal_9466 ), .Q ( new_AGEMA_signal_9467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4990 ( .C ( clk ), .D ( new_AGEMA_signal_9478 ), .Q ( new_AGEMA_signal_9479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5002 ( .C ( clk ), .D ( new_AGEMA_signal_9490 ), .Q ( new_AGEMA_signal_9491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5016 ( .C ( clk ), .D ( new_AGEMA_signal_9504 ), .Q ( new_AGEMA_signal_9505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5030 ( .C ( clk ), .D ( new_AGEMA_signal_9518 ), .Q ( new_AGEMA_signal_9519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5044 ( .C ( clk ), .D ( new_AGEMA_signal_9532 ), .Q ( new_AGEMA_signal_9533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5082 ( .C ( clk ), .D ( new_AGEMA_signal_9570 ), .Q ( new_AGEMA_signal_9571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5096 ( .C ( clk ), .D ( new_AGEMA_signal_9584 ), .Q ( new_AGEMA_signal_9585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5110 ( .C ( clk ), .D ( new_AGEMA_signal_9598 ), .Q ( new_AGEMA_signal_9599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5190 ( .C ( clk ), .D ( new_AGEMA_signal_9678 ), .Q ( new_AGEMA_signal_9679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5206 ( .C ( clk ), .D ( new_AGEMA_signal_9694 ), .Q ( new_AGEMA_signal_9695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5222 ( .C ( clk ), .D ( new_AGEMA_signal_9710 ), .Q ( new_AGEMA_signal_9711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5256 ( .C ( clk ), .D ( new_AGEMA_signal_9744 ), .Q ( new_AGEMA_signal_9745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5272 ( .C ( clk ), .D ( new_AGEMA_signal_9760 ), .Q ( new_AGEMA_signal_9761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5288 ( .C ( clk ), .D ( new_AGEMA_signal_9776 ), .Q ( new_AGEMA_signal_9777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5404 ( .C ( clk ), .D ( new_AGEMA_signal_9892 ), .Q ( new_AGEMA_signal_9893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5420 ( .C ( clk ), .D ( new_AGEMA_signal_9908 ), .Q ( new_AGEMA_signal_9909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5436 ( .C ( clk ), .D ( new_AGEMA_signal_9924 ), .Q ( new_AGEMA_signal_9925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5484 ( .C ( clk ), .D ( new_AGEMA_signal_9972 ), .Q ( new_AGEMA_signal_9973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5502 ( .C ( clk ), .D ( new_AGEMA_signal_9990 ), .Q ( new_AGEMA_signal_9991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5520 ( .C ( clk ), .D ( new_AGEMA_signal_10008 ), .Q ( new_AGEMA_signal_10009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5634 ( .C ( clk ), .D ( new_AGEMA_signal_10122 ), .Q ( new_AGEMA_signal_10123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5654 ( .C ( clk ), .D ( new_AGEMA_signal_10142 ), .Q ( new_AGEMA_signal_10143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5674 ( .C ( clk ), .D ( new_AGEMA_signal_10162 ), .Q ( new_AGEMA_signal_10163 ) ) ;

    /* cells in depth 11 */
    buf_clk new_AGEMA_reg_buffer_3249 ( .C ( clk ), .D ( n1934 ), .Q ( new_AGEMA_signal_7738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3251 ( .C ( clk ), .D ( new_AGEMA_signal_2228 ), .Q ( new_AGEMA_signal_7740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3253 ( .C ( clk ), .D ( new_AGEMA_signal_2229 ), .Q ( new_AGEMA_signal_7742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3261 ( .C ( clk ), .D ( new_AGEMA_signal_7749 ), .Q ( new_AGEMA_signal_7750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3269 ( .C ( clk ), .D ( new_AGEMA_signal_7757 ), .Q ( new_AGEMA_signal_7758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3277 ( .C ( clk ), .D ( new_AGEMA_signal_7765 ), .Q ( new_AGEMA_signal_7766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3279 ( .C ( clk ), .D ( n1981 ), .Q ( new_AGEMA_signal_7768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3281 ( .C ( clk ), .D ( new_AGEMA_signal_2244 ), .Q ( new_AGEMA_signal_7770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3283 ( .C ( clk ), .D ( new_AGEMA_signal_2245 ), .Q ( new_AGEMA_signal_7772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3287 ( .C ( clk ), .D ( new_AGEMA_signal_7775 ), .Q ( new_AGEMA_signal_7776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3291 ( .C ( clk ), .D ( new_AGEMA_signal_7779 ), .Q ( new_AGEMA_signal_7780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3295 ( .C ( clk ), .D ( new_AGEMA_signal_7783 ), .Q ( new_AGEMA_signal_7784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3303 ( .C ( clk ), .D ( new_AGEMA_signal_7791 ), .Q ( new_AGEMA_signal_7792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3311 ( .C ( clk ), .D ( new_AGEMA_signal_7799 ), .Q ( new_AGEMA_signal_7800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3319 ( .C ( clk ), .D ( new_AGEMA_signal_7807 ), .Q ( new_AGEMA_signal_7808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3321 ( .C ( clk ), .D ( new_AGEMA_signal_7103 ), .Q ( new_AGEMA_signal_7810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3323 ( .C ( clk ), .D ( new_AGEMA_signal_7111 ), .Q ( new_AGEMA_signal_7812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3325 ( .C ( clk ), .D ( new_AGEMA_signal_7119 ), .Q ( new_AGEMA_signal_7814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3331 ( .C ( clk ), .D ( new_AGEMA_signal_7819 ), .Q ( new_AGEMA_signal_7820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3337 ( .C ( clk ), .D ( new_AGEMA_signal_7825 ), .Q ( new_AGEMA_signal_7826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3343 ( .C ( clk ), .D ( new_AGEMA_signal_7831 ), .Q ( new_AGEMA_signal_7832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3347 ( .C ( clk ), .D ( new_AGEMA_signal_7835 ), .Q ( new_AGEMA_signal_7836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3351 ( .C ( clk ), .D ( new_AGEMA_signal_7839 ), .Q ( new_AGEMA_signal_7840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3355 ( .C ( clk ), .D ( new_AGEMA_signal_7843 ), .Q ( new_AGEMA_signal_7844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3363 ( .C ( clk ), .D ( new_AGEMA_signal_7851 ), .Q ( new_AGEMA_signal_7852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3371 ( .C ( clk ), .D ( new_AGEMA_signal_7859 ), .Q ( new_AGEMA_signal_7860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3379 ( .C ( clk ), .D ( new_AGEMA_signal_7867 ), .Q ( new_AGEMA_signal_7868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3383 ( .C ( clk ), .D ( new_AGEMA_signal_7871 ), .Q ( new_AGEMA_signal_7872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3387 ( .C ( clk ), .D ( new_AGEMA_signal_7875 ), .Q ( new_AGEMA_signal_7876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3391 ( .C ( clk ), .D ( new_AGEMA_signal_7879 ), .Q ( new_AGEMA_signal_7880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3397 ( .C ( clk ), .D ( new_AGEMA_signal_7885 ), .Q ( new_AGEMA_signal_7886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3403 ( .C ( clk ), .D ( new_AGEMA_signal_7891 ), .Q ( new_AGEMA_signal_7892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3409 ( .C ( clk ), .D ( new_AGEMA_signal_7897 ), .Q ( new_AGEMA_signal_7898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3415 ( .C ( clk ), .D ( new_AGEMA_signal_7903 ), .Q ( new_AGEMA_signal_7904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3421 ( .C ( clk ), .D ( new_AGEMA_signal_7909 ), .Q ( new_AGEMA_signal_7910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3427 ( .C ( clk ), .D ( new_AGEMA_signal_7915 ), .Q ( new_AGEMA_signal_7916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3433 ( .C ( clk ), .D ( new_AGEMA_signal_7921 ), .Q ( new_AGEMA_signal_7922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3439 ( .C ( clk ), .D ( new_AGEMA_signal_7927 ), .Q ( new_AGEMA_signal_7928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3445 ( .C ( clk ), .D ( new_AGEMA_signal_7933 ), .Q ( new_AGEMA_signal_7934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3451 ( .C ( clk ), .D ( new_AGEMA_signal_7939 ), .Q ( new_AGEMA_signal_7940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3457 ( .C ( clk ), .D ( new_AGEMA_signal_7945 ), .Q ( new_AGEMA_signal_7946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3463 ( .C ( clk ), .D ( new_AGEMA_signal_7951 ), .Q ( new_AGEMA_signal_7952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3469 ( .C ( clk ), .D ( new_AGEMA_signal_7957 ), .Q ( new_AGEMA_signal_7958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3475 ( .C ( clk ), .D ( new_AGEMA_signal_7963 ), .Q ( new_AGEMA_signal_7964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3481 ( .C ( clk ), .D ( new_AGEMA_signal_7969 ), .Q ( new_AGEMA_signal_7970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3485 ( .C ( clk ), .D ( new_AGEMA_signal_7973 ), .Q ( new_AGEMA_signal_7974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3489 ( .C ( clk ), .D ( new_AGEMA_signal_7977 ), .Q ( new_AGEMA_signal_7978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3493 ( .C ( clk ), .D ( new_AGEMA_signal_7981 ), .Q ( new_AGEMA_signal_7982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3501 ( .C ( clk ), .D ( new_AGEMA_signal_7989 ), .Q ( new_AGEMA_signal_7990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3509 ( .C ( clk ), .D ( new_AGEMA_signal_7997 ), .Q ( new_AGEMA_signal_7998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3517 ( .C ( clk ), .D ( new_AGEMA_signal_8005 ), .Q ( new_AGEMA_signal_8006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3521 ( .C ( clk ), .D ( new_AGEMA_signal_8009 ), .Q ( new_AGEMA_signal_8010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3525 ( .C ( clk ), .D ( new_AGEMA_signal_8013 ), .Q ( new_AGEMA_signal_8014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3529 ( .C ( clk ), .D ( new_AGEMA_signal_8017 ), .Q ( new_AGEMA_signal_8018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3535 ( .C ( clk ), .D ( new_AGEMA_signal_8023 ), .Q ( new_AGEMA_signal_8024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3541 ( .C ( clk ), .D ( new_AGEMA_signal_8029 ), .Q ( new_AGEMA_signal_8030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3547 ( .C ( clk ), .D ( new_AGEMA_signal_8035 ), .Q ( new_AGEMA_signal_8036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3555 ( .C ( clk ), .D ( new_AGEMA_signal_8043 ), .Q ( new_AGEMA_signal_8044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3563 ( .C ( clk ), .D ( new_AGEMA_signal_8051 ), .Q ( new_AGEMA_signal_8052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3571 ( .C ( clk ), .D ( new_AGEMA_signal_8059 ), .Q ( new_AGEMA_signal_8060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3573 ( .C ( clk ), .D ( new_AGEMA_signal_7523 ), .Q ( new_AGEMA_signal_8062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3575 ( .C ( clk ), .D ( new_AGEMA_signal_7525 ), .Q ( new_AGEMA_signal_8064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3577 ( .C ( clk ), .D ( new_AGEMA_signal_7527 ), .Q ( new_AGEMA_signal_8066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3583 ( .C ( clk ), .D ( new_AGEMA_signal_8071 ), .Q ( new_AGEMA_signal_8072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3589 ( .C ( clk ), .D ( new_AGEMA_signal_8077 ), .Q ( new_AGEMA_signal_8078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3595 ( .C ( clk ), .D ( new_AGEMA_signal_8083 ), .Q ( new_AGEMA_signal_8084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3597 ( .C ( clk ), .D ( n2410 ), .Q ( new_AGEMA_signal_8086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3599 ( .C ( clk ), .D ( new_AGEMA_signal_2322 ), .Q ( new_AGEMA_signal_8088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3601 ( .C ( clk ), .D ( new_AGEMA_signal_2323 ), .Q ( new_AGEMA_signal_8090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3603 ( .C ( clk ), .D ( n2421 ), .Q ( new_AGEMA_signal_8092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3605 ( .C ( clk ), .D ( new_AGEMA_signal_2324 ), .Q ( new_AGEMA_signal_8094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3607 ( .C ( clk ), .D ( new_AGEMA_signal_2325 ), .Q ( new_AGEMA_signal_8096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3613 ( .C ( clk ), .D ( new_AGEMA_signal_8101 ), .Q ( new_AGEMA_signal_8102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3619 ( .C ( clk ), .D ( new_AGEMA_signal_8107 ), .Q ( new_AGEMA_signal_8108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3625 ( .C ( clk ), .D ( new_AGEMA_signal_8113 ), .Q ( new_AGEMA_signal_8114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3631 ( .C ( clk ), .D ( new_AGEMA_signal_8119 ), .Q ( new_AGEMA_signal_8120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3637 ( .C ( clk ), .D ( new_AGEMA_signal_8125 ), .Q ( new_AGEMA_signal_8126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3643 ( .C ( clk ), .D ( new_AGEMA_signal_8131 ), .Q ( new_AGEMA_signal_8132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3651 ( .C ( clk ), .D ( new_AGEMA_signal_8139 ), .Q ( new_AGEMA_signal_8140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3659 ( .C ( clk ), .D ( new_AGEMA_signal_8147 ), .Q ( new_AGEMA_signal_8148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3667 ( .C ( clk ), .D ( new_AGEMA_signal_8155 ), .Q ( new_AGEMA_signal_8156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3675 ( .C ( clk ), .D ( new_AGEMA_signal_8163 ), .Q ( new_AGEMA_signal_8164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3683 ( .C ( clk ), .D ( new_AGEMA_signal_8171 ), .Q ( new_AGEMA_signal_8172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3691 ( .C ( clk ), .D ( new_AGEMA_signal_8179 ), .Q ( new_AGEMA_signal_8180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3697 ( .C ( clk ), .D ( new_AGEMA_signal_8185 ), .Q ( new_AGEMA_signal_8186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3703 ( .C ( clk ), .D ( new_AGEMA_signal_8191 ), .Q ( new_AGEMA_signal_8192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3709 ( .C ( clk ), .D ( new_AGEMA_signal_8197 ), .Q ( new_AGEMA_signal_8198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3715 ( .C ( clk ), .D ( new_AGEMA_signal_8203 ), .Q ( new_AGEMA_signal_8204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3721 ( .C ( clk ), .D ( new_AGEMA_signal_8209 ), .Q ( new_AGEMA_signal_8210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3727 ( .C ( clk ), .D ( new_AGEMA_signal_8215 ), .Q ( new_AGEMA_signal_8216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3729 ( .C ( clk ), .D ( new_AGEMA_signal_7495 ), .Q ( new_AGEMA_signal_8218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3731 ( .C ( clk ), .D ( new_AGEMA_signal_7499 ), .Q ( new_AGEMA_signal_8220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3733 ( .C ( clk ), .D ( new_AGEMA_signal_7503 ), .Q ( new_AGEMA_signal_8222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3737 ( .C ( clk ), .D ( new_AGEMA_signal_8225 ), .Q ( new_AGEMA_signal_8226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3741 ( .C ( clk ), .D ( new_AGEMA_signal_8229 ), .Q ( new_AGEMA_signal_8230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3745 ( .C ( clk ), .D ( new_AGEMA_signal_8233 ), .Q ( new_AGEMA_signal_8234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3749 ( .C ( clk ), .D ( new_AGEMA_signal_8237 ), .Q ( new_AGEMA_signal_8238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3753 ( .C ( clk ), .D ( new_AGEMA_signal_8241 ), .Q ( new_AGEMA_signal_8242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3757 ( .C ( clk ), .D ( new_AGEMA_signal_8245 ), .Q ( new_AGEMA_signal_8246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3761 ( .C ( clk ), .D ( new_AGEMA_signal_8249 ), .Q ( new_AGEMA_signal_8250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3765 ( .C ( clk ), .D ( new_AGEMA_signal_8253 ), .Q ( new_AGEMA_signal_8254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3769 ( .C ( clk ), .D ( new_AGEMA_signal_8257 ), .Q ( new_AGEMA_signal_8258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3771 ( .C ( clk ), .D ( new_AGEMA_signal_7331 ), .Q ( new_AGEMA_signal_8260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3773 ( .C ( clk ), .D ( new_AGEMA_signal_7339 ), .Q ( new_AGEMA_signal_8262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3775 ( .C ( clk ), .D ( new_AGEMA_signal_7347 ), .Q ( new_AGEMA_signal_8264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3779 ( .C ( clk ), .D ( new_AGEMA_signal_8267 ), .Q ( new_AGEMA_signal_8268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3785 ( .C ( clk ), .D ( new_AGEMA_signal_8273 ), .Q ( new_AGEMA_signal_8274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3791 ( .C ( clk ), .D ( new_AGEMA_signal_8279 ), .Q ( new_AGEMA_signal_8280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3801 ( .C ( clk ), .D ( n1984 ), .Q ( new_AGEMA_signal_8290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3805 ( .C ( clk ), .D ( new_AGEMA_signal_2396 ), .Q ( new_AGEMA_signal_8294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3809 ( .C ( clk ), .D ( new_AGEMA_signal_2397 ), .Q ( new_AGEMA_signal_8298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3817 ( .C ( clk ), .D ( new_AGEMA_signal_8305 ), .Q ( new_AGEMA_signal_8306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3825 ( .C ( clk ), .D ( new_AGEMA_signal_8313 ), .Q ( new_AGEMA_signal_8314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3833 ( .C ( clk ), .D ( new_AGEMA_signal_8321 ), .Q ( new_AGEMA_signal_8322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3841 ( .C ( clk ), .D ( new_AGEMA_signal_8329 ), .Q ( new_AGEMA_signal_8330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3849 ( .C ( clk ), .D ( new_AGEMA_signal_8337 ), .Q ( new_AGEMA_signal_8338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3857 ( .C ( clk ), .D ( new_AGEMA_signal_8345 ), .Q ( new_AGEMA_signal_8346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3865 ( .C ( clk ), .D ( new_AGEMA_signal_8353 ), .Q ( new_AGEMA_signal_8354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3873 ( .C ( clk ), .D ( new_AGEMA_signal_8361 ), .Q ( new_AGEMA_signal_8362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3881 ( .C ( clk ), .D ( new_AGEMA_signal_8369 ), .Q ( new_AGEMA_signal_8370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3889 ( .C ( clk ), .D ( new_AGEMA_signal_8377 ), .Q ( new_AGEMA_signal_8378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3897 ( .C ( clk ), .D ( new_AGEMA_signal_8385 ), .Q ( new_AGEMA_signal_8386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3905 ( .C ( clk ), .D ( new_AGEMA_signal_8393 ), .Q ( new_AGEMA_signal_8394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3911 ( .C ( clk ), .D ( new_AGEMA_signal_8399 ), .Q ( new_AGEMA_signal_8400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3917 ( .C ( clk ), .D ( new_AGEMA_signal_8405 ), .Q ( new_AGEMA_signal_8406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3923 ( .C ( clk ), .D ( new_AGEMA_signal_8411 ), .Q ( new_AGEMA_signal_8412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3933 ( .C ( clk ), .D ( new_AGEMA_signal_8421 ), .Q ( new_AGEMA_signal_8422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3943 ( .C ( clk ), .D ( new_AGEMA_signal_8431 ), .Q ( new_AGEMA_signal_8432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3953 ( .C ( clk ), .D ( new_AGEMA_signal_8441 ), .Q ( new_AGEMA_signal_8442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3961 ( .C ( clk ), .D ( new_AGEMA_signal_8449 ), .Q ( new_AGEMA_signal_8450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3969 ( .C ( clk ), .D ( new_AGEMA_signal_8457 ), .Q ( new_AGEMA_signal_8458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3977 ( .C ( clk ), .D ( new_AGEMA_signal_8465 ), .Q ( new_AGEMA_signal_8466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3985 ( .C ( clk ), .D ( new_AGEMA_signal_8473 ), .Q ( new_AGEMA_signal_8474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3993 ( .C ( clk ), .D ( new_AGEMA_signal_8481 ), .Q ( new_AGEMA_signal_8482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4001 ( .C ( clk ), .D ( new_AGEMA_signal_8489 ), .Q ( new_AGEMA_signal_8490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4009 ( .C ( clk ), .D ( new_AGEMA_signal_8497 ), .Q ( new_AGEMA_signal_8498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4017 ( .C ( clk ), .D ( new_AGEMA_signal_8505 ), .Q ( new_AGEMA_signal_8506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4025 ( .C ( clk ), .D ( new_AGEMA_signal_8513 ), .Q ( new_AGEMA_signal_8514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4035 ( .C ( clk ), .D ( new_AGEMA_signal_7513 ), .Q ( new_AGEMA_signal_8524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4039 ( .C ( clk ), .D ( new_AGEMA_signal_7517 ), .Q ( new_AGEMA_signal_8528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4043 ( .C ( clk ), .D ( new_AGEMA_signal_7521 ), .Q ( new_AGEMA_signal_8532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4049 ( .C ( clk ), .D ( new_AGEMA_signal_8537 ), .Q ( new_AGEMA_signal_8538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4055 ( .C ( clk ), .D ( new_AGEMA_signal_8543 ), .Q ( new_AGEMA_signal_8544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4061 ( .C ( clk ), .D ( new_AGEMA_signal_8549 ), .Q ( new_AGEMA_signal_8550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4065 ( .C ( clk ), .D ( new_AGEMA_signal_7179 ), .Q ( new_AGEMA_signal_8554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4069 ( .C ( clk ), .D ( new_AGEMA_signal_7185 ), .Q ( new_AGEMA_signal_8558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4073 ( .C ( clk ), .D ( new_AGEMA_signal_7191 ), .Q ( new_AGEMA_signal_8562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4083 ( .C ( clk ), .D ( new_AGEMA_signal_8571 ), .Q ( new_AGEMA_signal_8572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4093 ( .C ( clk ), .D ( new_AGEMA_signal_8581 ), .Q ( new_AGEMA_signal_8582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4103 ( .C ( clk ), .D ( new_AGEMA_signal_8591 ), .Q ( new_AGEMA_signal_8592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4111 ( .C ( clk ), .D ( new_AGEMA_signal_8599 ), .Q ( new_AGEMA_signal_8600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4119 ( .C ( clk ), .D ( new_AGEMA_signal_8607 ), .Q ( new_AGEMA_signal_8608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4127 ( .C ( clk ), .D ( new_AGEMA_signal_8615 ), .Q ( new_AGEMA_signal_8616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4131 ( .C ( clk ), .D ( n2478 ), .Q ( new_AGEMA_signal_8620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4135 ( .C ( clk ), .D ( new_AGEMA_signal_2164 ), .Q ( new_AGEMA_signal_8624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4139 ( .C ( clk ), .D ( new_AGEMA_signal_2165 ), .Q ( new_AGEMA_signal_8628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4153 ( .C ( clk ), .D ( new_AGEMA_signal_8641 ), .Q ( new_AGEMA_signal_8642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4161 ( .C ( clk ), .D ( new_AGEMA_signal_8649 ), .Q ( new_AGEMA_signal_8650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4169 ( .C ( clk ), .D ( new_AGEMA_signal_8657 ), .Q ( new_AGEMA_signal_8658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4177 ( .C ( clk ), .D ( new_AGEMA_signal_8665 ), .Q ( new_AGEMA_signal_8666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4185 ( .C ( clk ), .D ( new_AGEMA_signal_8673 ), .Q ( new_AGEMA_signal_8674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4193 ( .C ( clk ), .D ( new_AGEMA_signal_8681 ), .Q ( new_AGEMA_signal_8682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4199 ( .C ( clk ), .D ( new_AGEMA_signal_8687 ), .Q ( new_AGEMA_signal_8688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4205 ( .C ( clk ), .D ( new_AGEMA_signal_8693 ), .Q ( new_AGEMA_signal_8694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4211 ( .C ( clk ), .D ( new_AGEMA_signal_8699 ), .Q ( new_AGEMA_signal_8700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4215 ( .C ( clk ), .D ( n2660 ), .Q ( new_AGEMA_signal_8704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4219 ( .C ( clk ), .D ( new_AGEMA_signal_2364 ), .Q ( new_AGEMA_signal_8708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4223 ( .C ( clk ), .D ( new_AGEMA_signal_2365 ), .Q ( new_AGEMA_signal_8712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4231 ( .C ( clk ), .D ( new_AGEMA_signal_8719 ), .Q ( new_AGEMA_signal_8720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4239 ( .C ( clk ), .D ( new_AGEMA_signal_8727 ), .Q ( new_AGEMA_signal_8728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4247 ( .C ( clk ), .D ( new_AGEMA_signal_8735 ), .Q ( new_AGEMA_signal_8736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4257 ( .C ( clk ), .D ( n1940 ), .Q ( new_AGEMA_signal_8746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4263 ( .C ( clk ), .D ( new_AGEMA_signal_2232 ), .Q ( new_AGEMA_signal_8752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4269 ( .C ( clk ), .D ( new_AGEMA_signal_2233 ), .Q ( new_AGEMA_signal_8758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4275 ( .C ( clk ), .D ( n1961 ), .Q ( new_AGEMA_signal_8764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4281 ( .C ( clk ), .D ( new_AGEMA_signal_2234 ), .Q ( new_AGEMA_signal_8770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4287 ( .C ( clk ), .D ( new_AGEMA_signal_2235 ), .Q ( new_AGEMA_signal_8776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4293 ( .C ( clk ), .D ( n1987 ), .Q ( new_AGEMA_signal_8782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4299 ( .C ( clk ), .D ( new_AGEMA_signal_2028 ), .Q ( new_AGEMA_signal_8788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4305 ( .C ( clk ), .D ( new_AGEMA_signal_2029 ), .Q ( new_AGEMA_signal_8794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4325 ( .C ( clk ), .D ( new_AGEMA_signal_8813 ), .Q ( new_AGEMA_signal_8814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4333 ( .C ( clk ), .D ( new_AGEMA_signal_8821 ), .Q ( new_AGEMA_signal_8822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4341 ( .C ( clk ), .D ( new_AGEMA_signal_8829 ), .Q ( new_AGEMA_signal_8830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4347 ( .C ( clk ), .D ( n2054 ), .Q ( new_AGEMA_signal_8836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4353 ( .C ( clk ), .D ( new_AGEMA_signal_2254 ), .Q ( new_AGEMA_signal_8842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4359 ( .C ( clk ), .D ( new_AGEMA_signal_2255 ), .Q ( new_AGEMA_signal_8848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4379 ( .C ( clk ), .D ( new_AGEMA_signal_8867 ), .Q ( new_AGEMA_signal_8868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4387 ( .C ( clk ), .D ( new_AGEMA_signal_8875 ), .Q ( new_AGEMA_signal_8876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4395 ( .C ( clk ), .D ( new_AGEMA_signal_8883 ), .Q ( new_AGEMA_signal_8884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4403 ( .C ( clk ), .D ( new_AGEMA_signal_8891 ), .Q ( new_AGEMA_signal_8892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4411 ( .C ( clk ), .D ( new_AGEMA_signal_8899 ), .Q ( new_AGEMA_signal_8900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4419 ( .C ( clk ), .D ( new_AGEMA_signal_8907 ), .Q ( new_AGEMA_signal_8908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4429 ( .C ( clk ), .D ( new_AGEMA_signal_8917 ), .Q ( new_AGEMA_signal_8918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4439 ( .C ( clk ), .D ( new_AGEMA_signal_8927 ), .Q ( new_AGEMA_signal_8928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4449 ( .C ( clk ), .D ( new_AGEMA_signal_8937 ), .Q ( new_AGEMA_signal_8938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4457 ( .C ( clk ), .D ( new_AGEMA_signal_8945 ), .Q ( new_AGEMA_signal_8946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4465 ( .C ( clk ), .D ( new_AGEMA_signal_8953 ), .Q ( new_AGEMA_signal_8954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4473 ( .C ( clk ), .D ( new_AGEMA_signal_8961 ), .Q ( new_AGEMA_signal_8962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4479 ( .C ( clk ), .D ( n2255 ), .Q ( new_AGEMA_signal_8968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4485 ( .C ( clk ), .D ( new_AGEMA_signal_2294 ), .Q ( new_AGEMA_signal_8974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4491 ( .C ( clk ), .D ( new_AGEMA_signal_2295 ), .Q ( new_AGEMA_signal_8980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4509 ( .C ( clk ), .D ( n2304 ), .Q ( new_AGEMA_signal_8998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4515 ( .C ( clk ), .D ( new_AGEMA_signal_2302 ), .Q ( new_AGEMA_signal_9004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4521 ( .C ( clk ), .D ( new_AGEMA_signal_2303 ), .Q ( new_AGEMA_signal_9010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4529 ( .C ( clk ), .D ( new_AGEMA_signal_9017 ), .Q ( new_AGEMA_signal_9018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4537 ( .C ( clk ), .D ( new_AGEMA_signal_9025 ), .Q ( new_AGEMA_signal_9026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4545 ( .C ( clk ), .D ( new_AGEMA_signal_9033 ), .Q ( new_AGEMA_signal_9034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4551 ( .C ( clk ), .D ( n2450 ), .Q ( new_AGEMA_signal_9040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4557 ( .C ( clk ), .D ( new_AGEMA_signal_2330 ), .Q ( new_AGEMA_signal_9046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4563 ( .C ( clk ), .D ( new_AGEMA_signal_2331 ), .Q ( new_AGEMA_signal_9052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4577 ( .C ( clk ), .D ( new_AGEMA_signal_9065 ), .Q ( new_AGEMA_signal_9066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4585 ( .C ( clk ), .D ( new_AGEMA_signal_9073 ), .Q ( new_AGEMA_signal_9074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4593 ( .C ( clk ), .D ( new_AGEMA_signal_9081 ), .Q ( new_AGEMA_signal_9082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4611 ( .C ( clk ), .D ( n2666 ), .Q ( new_AGEMA_signal_9100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4617 ( .C ( clk ), .D ( new_AGEMA_signal_2368 ), .Q ( new_AGEMA_signal_9106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4623 ( .C ( clk ), .D ( new_AGEMA_signal_2369 ), .Q ( new_AGEMA_signal_9112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4629 ( .C ( clk ), .D ( n2704 ), .Q ( new_AGEMA_signal_9118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4635 ( .C ( clk ), .D ( new_AGEMA_signal_2372 ), .Q ( new_AGEMA_signal_9124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4641 ( .C ( clk ), .D ( new_AGEMA_signal_2373 ), .Q ( new_AGEMA_signal_9130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4709 ( .C ( clk ), .D ( new_AGEMA_signal_9197 ), .Q ( new_AGEMA_signal_9198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4719 ( .C ( clk ), .D ( new_AGEMA_signal_9207 ), .Q ( new_AGEMA_signal_9208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4729 ( .C ( clk ), .D ( new_AGEMA_signal_9217 ), .Q ( new_AGEMA_signal_9218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4797 ( .C ( clk ), .D ( n2280 ), .Q ( new_AGEMA_signal_9286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4805 ( .C ( clk ), .D ( new_AGEMA_signal_2110 ), .Q ( new_AGEMA_signal_9294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4813 ( .C ( clk ), .D ( new_AGEMA_signal_2111 ), .Q ( new_AGEMA_signal_9302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4839 ( .C ( clk ), .D ( new_AGEMA_signal_7169 ), .Q ( new_AGEMA_signal_9328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4847 ( .C ( clk ), .D ( new_AGEMA_signal_7171 ), .Q ( new_AGEMA_signal_9336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4855 ( .C ( clk ), .D ( new_AGEMA_signal_7173 ), .Q ( new_AGEMA_signal_9344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4863 ( .C ( clk ), .D ( n2456 ), .Q ( new_AGEMA_signal_9352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4871 ( .C ( clk ), .D ( new_AGEMA_signal_2332 ), .Q ( new_AGEMA_signal_9360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4879 ( .C ( clk ), .D ( new_AGEMA_signal_2333 ), .Q ( new_AGEMA_signal_9368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4917 ( .C ( clk ), .D ( n2706 ), .Q ( new_AGEMA_signal_9406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4925 ( .C ( clk ), .D ( new_AGEMA_signal_2370 ), .Q ( new_AGEMA_signal_9414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4933 ( .C ( clk ), .D ( new_AGEMA_signal_2371 ), .Q ( new_AGEMA_signal_9422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4979 ( .C ( clk ), .D ( new_AGEMA_signal_9467 ), .Q ( new_AGEMA_signal_9468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4991 ( .C ( clk ), .D ( new_AGEMA_signal_9479 ), .Q ( new_AGEMA_signal_9480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5003 ( .C ( clk ), .D ( new_AGEMA_signal_9491 ), .Q ( new_AGEMA_signal_9492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5017 ( .C ( clk ), .D ( new_AGEMA_signal_9505 ), .Q ( new_AGEMA_signal_9506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5031 ( .C ( clk ), .D ( new_AGEMA_signal_9519 ), .Q ( new_AGEMA_signal_9520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5045 ( .C ( clk ), .D ( new_AGEMA_signal_9533 ), .Q ( new_AGEMA_signal_9534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5083 ( .C ( clk ), .D ( new_AGEMA_signal_9571 ), .Q ( new_AGEMA_signal_9572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5097 ( .C ( clk ), .D ( new_AGEMA_signal_9585 ), .Q ( new_AGEMA_signal_9586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5111 ( .C ( clk ), .D ( new_AGEMA_signal_9599 ), .Q ( new_AGEMA_signal_9600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5191 ( .C ( clk ), .D ( new_AGEMA_signal_9679 ), .Q ( new_AGEMA_signal_9680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5207 ( .C ( clk ), .D ( new_AGEMA_signal_9695 ), .Q ( new_AGEMA_signal_9696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5223 ( .C ( clk ), .D ( new_AGEMA_signal_9711 ), .Q ( new_AGEMA_signal_9712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5257 ( .C ( clk ), .D ( new_AGEMA_signal_9745 ), .Q ( new_AGEMA_signal_9746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5273 ( .C ( clk ), .D ( new_AGEMA_signal_9761 ), .Q ( new_AGEMA_signal_9762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5289 ( .C ( clk ), .D ( new_AGEMA_signal_9777 ), .Q ( new_AGEMA_signal_9778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5405 ( .C ( clk ), .D ( new_AGEMA_signal_9893 ), .Q ( new_AGEMA_signal_9894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5421 ( .C ( clk ), .D ( new_AGEMA_signal_9909 ), .Q ( new_AGEMA_signal_9910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5437 ( .C ( clk ), .D ( new_AGEMA_signal_9925 ), .Q ( new_AGEMA_signal_9926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5485 ( .C ( clk ), .D ( new_AGEMA_signal_9973 ), .Q ( new_AGEMA_signal_9974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5503 ( .C ( clk ), .D ( new_AGEMA_signal_9991 ), .Q ( new_AGEMA_signal_9992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5521 ( .C ( clk ), .D ( new_AGEMA_signal_10009 ), .Q ( new_AGEMA_signal_10010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5635 ( .C ( clk ), .D ( new_AGEMA_signal_10123 ), .Q ( new_AGEMA_signal_10124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5655 ( .C ( clk ), .D ( new_AGEMA_signal_10143 ), .Q ( new_AGEMA_signal_10144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5675 ( .C ( clk ), .D ( new_AGEMA_signal_10163 ), .Q ( new_AGEMA_signal_10164 ) ) ;

    /* cells in depth 12 */
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2001 ( .a ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, n1932}), .b ({new_AGEMA_signal_7053, new_AGEMA_signal_7049, new_AGEMA_signal_7045}), .clk ( clk ), .r ({Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, n1933}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2051 ( .a ({new_AGEMA_signal_7065, new_AGEMA_signal_7061, new_AGEMA_signal_7057}), .b ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, n1955}), .clk ( clk ), .r ({Fresh[1985], Fresh[1984], Fresh[1983]}), .c ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, n1958}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2067 ( .a ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, n1967}), .b ({new_AGEMA_signal_7089, new_AGEMA_signal_7081, new_AGEMA_signal_7073}), .clk ( clk ), .r ({Fresh[1988], Fresh[1987], Fresh[1986]}), .c ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, n1990}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2104 ( .a ({new_AGEMA_signal_7095, new_AGEMA_signal_7093, new_AGEMA_signal_7091}), .b ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, n1977}), .clk ( clk ), .r ({Fresh[1991], Fresh[1990], Fresh[1989]}), .c ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, n1982}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2128 ( .a ({new_AGEMA_signal_7119, new_AGEMA_signal_7111, new_AGEMA_signal_7103}), .b ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, n1998}), .clk ( clk ), .r ({Fresh[1994], Fresh[1993], Fresh[1992]}), .c ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, n1999}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2148 ( .a ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, n2010}), .b ({new_AGEMA_signal_7137, new_AGEMA_signal_7131, new_AGEMA_signal_7125}), .clk ( clk ), .r ({Fresh[1997], Fresh[1996], Fresh[1995]}), .c ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, n2011}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2165 ( .a ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, n2024}), .b ({new_AGEMA_signal_7149, new_AGEMA_signal_7145, new_AGEMA_signal_7141}), .clk ( clk ), .r ({Fresh[2000], Fresh[1999], Fresh[1998]}), .c ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, n2025}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2179 ( .a ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, n2035}), .b ({new_AGEMA_signal_7167, new_AGEMA_signal_7161, new_AGEMA_signal_7155}), .clk ( clk ), .r ({Fresh[2003], Fresh[2002], Fresh[2001]}), .c ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, n2036}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2196 ( .a ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, n2048}), .b ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, n2047}), .clk ( clk ), .r ({Fresh[2006], Fresh[2005], Fresh[2004]}), .c ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, n2049}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2207 ( .a ({new_AGEMA_signal_7173, new_AGEMA_signal_7171, new_AGEMA_signal_7169}), .b ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, n2059}), .clk ( clk ), .r ({Fresh[2009], Fresh[2008], Fresh[2007]}), .c ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, n2072}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2214 ( .a ({new_AGEMA_signal_7191, new_AGEMA_signal_7185, new_AGEMA_signal_7179}), .b ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, n2064}), .clk ( clk ), .r ({Fresh[2012], Fresh[2011], Fresh[2010]}), .c ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, n2067}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2230 ( .a ({new_AGEMA_signal_7209, new_AGEMA_signal_7203, new_AGEMA_signal_7197}), .b ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, n2077}), .clk ( clk ), .r ({Fresh[2015], Fresh[2014], Fresh[2013]}), .c ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, n2078}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2250 ( .a ({new_AGEMA_signal_7215, new_AGEMA_signal_7213, new_AGEMA_signal_7211}), .b ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, n2158}), .clk ( clk ), .r ({Fresh[2018], Fresh[2017], Fresh[2016]}), .c ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, n2097}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2257 ( .a ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, n2095}), .b ({new_AGEMA_signal_7227, new_AGEMA_signal_7223, new_AGEMA_signal_7219}), .clk ( clk ), .r ({Fresh[2021], Fresh[2020], Fresh[2019]}), .c ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, n2096}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2275 ( .a ({new_AGEMA_signal_7245, new_AGEMA_signal_7239, new_AGEMA_signal_7233}), .b ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, n2117}), .clk ( clk ), .r ({Fresh[2024], Fresh[2023], Fresh[2022]}), .c ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, n2128}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2285 ( .a ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, n2123}), .b ({new_AGEMA_signal_7263, new_AGEMA_signal_7257, new_AGEMA_signal_7251}), .clk ( clk ), .r ({Fresh[2027], Fresh[2026], Fresh[2025]}), .c ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, n2124}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2301 ( .a ({new_AGEMA_signal_7269, new_AGEMA_signal_7267, new_AGEMA_signal_7265}), .b ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, n2135}), .clk ( clk ), .r ({Fresh[2030], Fresh[2029], Fresh[2028]}), .c ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, n2148}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2310 ( .a ({new_AGEMA_signal_7287, new_AGEMA_signal_7281, new_AGEMA_signal_7275}), .b ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, n2141}), .clk ( clk ), .r ({Fresh[2033], Fresh[2032], Fresh[2031]}), .c ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, n2142}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2325 ( .a ({new_AGEMA_signal_7293, new_AGEMA_signal_7291, new_AGEMA_signal_7289}), .b ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, n2158}), .clk ( clk ), .r ({Fresh[2036], Fresh[2035], Fresh[2034]}), .c ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, n2168}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2332 ( .a ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, n2166}), .b ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, n2165}), .clk ( clk ), .r ({Fresh[2039], Fresh[2038], Fresh[2037]}), .c ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, n2167}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2347 ( .a ({new_AGEMA_signal_7305, new_AGEMA_signal_7301, new_AGEMA_signal_7297}), .b ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, n2180}), .clk ( clk ), .r ({Fresh[2042], Fresh[2041], Fresh[2040]}), .c ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, n2184}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2361 ( .a ({new_AGEMA_signal_7317, new_AGEMA_signal_7313, new_AGEMA_signal_7309}), .b ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, n2194}), .clk ( clk ), .r ({Fresh[2045], Fresh[2044], Fresh[2043]}), .c ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, n2197}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2373 ( .a ({new_AGEMA_signal_7323, new_AGEMA_signal_7321, new_AGEMA_signal_7319}), .b ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, n2204}), .clk ( clk ), .r ({Fresh[2048], Fresh[2047], Fresh[2046]}), .c ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, n2205}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2390 ( .a ({new_AGEMA_signal_7347, new_AGEMA_signal_7339, new_AGEMA_signal_7331}), .b ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, n2225}), .clk ( clk ), .r ({Fresh[2051], Fresh[2050], Fresh[2049]}), .c ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, n2232}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2395 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, n2230}), .b ({new_AGEMA_signal_7365, new_AGEMA_signal_7359, new_AGEMA_signal_7353}), .clk ( clk ), .r ({Fresh[2054], Fresh[2053], Fresh[2052]}), .c ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, n2231}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2401 ( .a ({new_AGEMA_signal_7377, new_AGEMA_signal_7373, new_AGEMA_signal_7369}), .b ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, n2236}), .clk ( clk ), .r ({Fresh[2057], Fresh[2056], Fresh[2055]}), .c ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, n2239}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2413 ( .a ({new_AGEMA_signal_7389, new_AGEMA_signal_7385, new_AGEMA_signal_7381}), .b ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, n2247}), .clk ( clk ), .r ({Fresh[2060], Fresh[2059], Fresh[2058]}), .c ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, n2250}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2428 ( .a ({new_AGEMA_signal_7173, new_AGEMA_signal_7171, new_AGEMA_signal_7169}), .b ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, n2264}), .clk ( clk ), .r ({Fresh[2063], Fresh[2062], Fresh[2061]}), .c ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, n2276}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2439 ( .a ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, n2271}), .b ({new_AGEMA_signal_7395, new_AGEMA_signal_7393, new_AGEMA_signal_7391}), .clk ( clk ), .r ({Fresh[2066], Fresh[2065], Fresh[2064]}), .c ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, n2272}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2454 ( .a ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, n2286}), .b ({new_AGEMA_signal_7401, new_AGEMA_signal_7399, new_AGEMA_signal_7397}), .clk ( clk ), .r ({Fresh[2069], Fresh[2068], Fresh[2067]}), .c ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, n2306}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2468 ( .a ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, n2295}), .b ({new_AGEMA_signal_7413, new_AGEMA_signal_7409, new_AGEMA_signal_7405}), .clk ( clk ), .r ({Fresh[2072], Fresh[2071], Fresh[2070]}), .c ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, n2296}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2489 ( .a ({new_AGEMA_signal_7425, new_AGEMA_signal_7421, new_AGEMA_signal_7417}), .b ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, n2322}), .clk ( clk ), .r ({Fresh[2075], Fresh[2074], Fresh[2073]}), .c ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, n2324}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2500 ( .a ({new_AGEMA_signal_7431, new_AGEMA_signal_7429, new_AGEMA_signal_7427}), .b ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, n2333}), .clk ( clk ), .r ({Fresh[2078], Fresh[2077], Fresh[2076]}), .c ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, n2337}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2511 ( .a ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, n2345}), .b ({new_AGEMA_signal_7449, new_AGEMA_signal_7443, new_AGEMA_signal_7437}), .clk ( clk ), .r ({Fresh[2081], Fresh[2080], Fresh[2079]}), .c ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, n2350}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2528 ( .a ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, n2361}), .b ({new_AGEMA_signal_7461, new_AGEMA_signal_7457, new_AGEMA_signal_7453}), .clk ( clk ), .r ({Fresh[2084], Fresh[2083], Fresh[2082]}), .c ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, n2362}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2550 ( .a ({new_AGEMA_signal_7467, new_AGEMA_signal_7465, new_AGEMA_signal_7463}), .b ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, n2388}), .clk ( clk ), .r ({Fresh[2087], Fresh[2086], Fresh[2085]}), .c ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, n2389}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2557 ( .a ({new_AGEMA_signal_7479, new_AGEMA_signal_7475, new_AGEMA_signal_7471}), .b ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, n2393}), .clk ( clk ), .r ({Fresh[2090], Fresh[2089], Fresh[2088]}), .c ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, n2397}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2568 ( .a ({new_AGEMA_signal_7491, new_AGEMA_signal_7487, new_AGEMA_signal_7483}), .b ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, n2405}), .clk ( clk ), .r ({Fresh[2093], Fresh[2092], Fresh[2091]}), .c ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, n2411}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2580 ( .a ({new_AGEMA_signal_7503, new_AGEMA_signal_7499, new_AGEMA_signal_7495}), .b ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, n2419}), .clk ( clk ), .r ({Fresh[2096], Fresh[2095], Fresh[2094]}), .c ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, n2420}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2593 ( .a ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, n2436}), .b ({new_AGEMA_signal_7509, new_AGEMA_signal_7507, new_AGEMA_signal_7505}), .clk ( clk ), .r ({Fresh[2099], Fresh[2098], Fresh[2097]}), .c ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, n2440}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2614 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7517, new_AGEMA_signal_7513}), .b ({new_AGEMA_signal_2335, new_AGEMA_signal_2334, n2461}), .clk ( clk ), .r ({Fresh[2102], Fresh[2101], Fresh[2100]}), .c ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, n2516}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) U2621 ( .s ({new_AGEMA_signal_7527, new_AGEMA_signal_7525, new_AGEMA_signal_7523}), .b ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, n2469}), .a ({new_AGEMA_signal_7545, new_AGEMA_signal_7539, new_AGEMA_signal_7533}), .clk ( clk ), .r ({Fresh[2105], Fresh[2104], Fresh[2103]}), .c ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, n2471}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2636 ( .a ({new_AGEMA_signal_7563, new_AGEMA_signal_7557, new_AGEMA_signal_7551}), .b ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, n2484}), .clk ( clk ), .r ({Fresh[2108], Fresh[2107], Fresh[2106]}), .c ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, n2485}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2644 ( .a ({new_AGEMA_signal_7191, new_AGEMA_signal_7185, new_AGEMA_signal_7179}), .b ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, n2491}), .clk ( clk ), .r ({Fresh[2111], Fresh[2110], Fresh[2109]}), .c ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, n2502}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2651 ( .a ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, n2500}), .b ({new_AGEMA_signal_7575, new_AGEMA_signal_7571, new_AGEMA_signal_7567}), .clk ( clk ), .r ({Fresh[2114], Fresh[2113], Fresh[2112]}), .c ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, n2501}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2657 ( .a ({new_AGEMA_signal_7503, new_AGEMA_signal_7499, new_AGEMA_signal_7495}), .b ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, n2508}), .clk ( clk ), .r ({Fresh[2117], Fresh[2116], Fresh[2115]}), .c ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, n2509}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2671 ( .a ({new_AGEMA_signal_7581, new_AGEMA_signal_7579, new_AGEMA_signal_7577}), .b ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, n2526}), .clk ( clk ), .r ({Fresh[2120], Fresh[2119], Fresh[2118]}), .c ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, n2527}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2680 ( .a ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, n2539}), .b ({new_AGEMA_signal_7605, new_AGEMA_signal_7597, new_AGEMA_signal_7589}), .clk ( clk ), .r ({Fresh[2123], Fresh[2122], Fresh[2121]}), .c ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, n2550}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2685 ( .a ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, n2548}), .b ({new_AGEMA_signal_7611, new_AGEMA_signal_7609, new_AGEMA_signal_7607}), .clk ( clk ), .r ({Fresh[2126], Fresh[2125], Fresh[2124]}), .c ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, n2549}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2701 ( .a ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, n2568}), .b ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, n2567}), .clk ( clk ), .r ({Fresh[2129], Fresh[2128], Fresh[2127]}), .c ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, n2569}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2712 ( .a ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, n2583}), .b ({new_AGEMA_signal_7623, new_AGEMA_signal_7619, new_AGEMA_signal_7615}), .clk ( clk ), .r ({Fresh[2132], Fresh[2131], Fresh[2130]}), .c ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, n2584}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2729 ( .a ({new_AGEMA_signal_7635, new_AGEMA_signal_7631, new_AGEMA_signal_7627}), .b ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, n2604}), .clk ( clk ), .r ({Fresh[2135], Fresh[2134], Fresh[2133]}), .c ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, n2606}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2740 ( .a ({new_AGEMA_signal_7191, new_AGEMA_signal_7185, new_AGEMA_signal_7179}), .b ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, n2621}), .clk ( clk ), .r ({Fresh[2138], Fresh[2137], Fresh[2136]}), .c ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, n2622}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2747 ( .a ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, n2633}), .b ({new_AGEMA_signal_7647, new_AGEMA_signal_7643, new_AGEMA_signal_7639}), .clk ( clk ), .r ({Fresh[2141], Fresh[2140], Fresh[2139]}), .c ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, n2634}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2761 ( .a ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, n2656}), .b ({new_AGEMA_signal_7659, new_AGEMA_signal_7655, new_AGEMA_signal_7651}), .clk ( clk ), .r ({Fresh[2144], Fresh[2143], Fresh[2142]}), .c ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, n2657}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2783 ( .a ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, n2696}), .b ({new_AGEMA_signal_7671, new_AGEMA_signal_7667, new_AGEMA_signal_7663}), .clk ( clk ), .r ({Fresh[2147], Fresh[2146], Fresh[2145]}), .c ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, n2697}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2795 ( .a ({new_AGEMA_signal_7173, new_AGEMA_signal_7171, new_AGEMA_signal_7169}), .b ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, n2718}), .clk ( clk ), .r ({Fresh[2150], Fresh[2149], Fresh[2148]}), .c ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, n2808}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2802 ( .a ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, n2730}), .b ({new_AGEMA_signal_7695, new_AGEMA_signal_7687, new_AGEMA_signal_7679}), .clk ( clk ), .r ({Fresh[2153], Fresh[2152], Fresh[2151]}), .c ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, n2747}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2810 ( .a ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, n2745}), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, n2744}), .clk ( clk ), .r ({Fresh[2156], Fresh[2155], Fresh[2154]}), .c ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, n2746}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2818 ( .a ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, n2759}), .b ({new_AGEMA_signal_7701, new_AGEMA_signal_7699, new_AGEMA_signal_7697}), .clk ( clk ), .r ({Fresh[2159], Fresh[2158], Fresh[2157]}), .c ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, n2804}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2824 ( .a ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, n2771}), .b ({new_AGEMA_signal_7713, new_AGEMA_signal_7709, new_AGEMA_signal_7705}), .clk ( clk ), .r ({Fresh[2162], Fresh[2161], Fresh[2160]}), .c ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, n2802}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2838 ( .a ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, n2798}), .b ({new_AGEMA_signal_7719, new_AGEMA_signal_7717, new_AGEMA_signal_7715}), .clk ( clk ), .r ({Fresh[2165], Fresh[2164], Fresh[2163]}), .c ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, n2799}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2852 ( .a ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, n2826}), .b ({new_AGEMA_signal_7737, new_AGEMA_signal_7731, new_AGEMA_signal_7725}), .clk ( clk ), .r ({Fresh[2168], Fresh[2167], Fresh[2166]}), .c ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, n2827}) ) ;
    buf_clk new_AGEMA_reg_buffer_3250 ( .C ( clk ), .D ( new_AGEMA_signal_7738 ), .Q ( new_AGEMA_signal_7739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3252 ( .C ( clk ), .D ( new_AGEMA_signal_7740 ), .Q ( new_AGEMA_signal_7741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3254 ( .C ( clk ), .D ( new_AGEMA_signal_7742 ), .Q ( new_AGEMA_signal_7743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3262 ( .C ( clk ), .D ( new_AGEMA_signal_7750 ), .Q ( new_AGEMA_signal_7751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3270 ( .C ( clk ), .D ( new_AGEMA_signal_7758 ), .Q ( new_AGEMA_signal_7759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3278 ( .C ( clk ), .D ( new_AGEMA_signal_7766 ), .Q ( new_AGEMA_signal_7767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3280 ( .C ( clk ), .D ( new_AGEMA_signal_7768 ), .Q ( new_AGEMA_signal_7769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3282 ( .C ( clk ), .D ( new_AGEMA_signal_7770 ), .Q ( new_AGEMA_signal_7771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3284 ( .C ( clk ), .D ( new_AGEMA_signal_7772 ), .Q ( new_AGEMA_signal_7773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3288 ( .C ( clk ), .D ( new_AGEMA_signal_7776 ), .Q ( new_AGEMA_signal_7777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3292 ( .C ( clk ), .D ( new_AGEMA_signal_7780 ), .Q ( new_AGEMA_signal_7781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3296 ( .C ( clk ), .D ( new_AGEMA_signal_7784 ), .Q ( new_AGEMA_signal_7785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3304 ( .C ( clk ), .D ( new_AGEMA_signal_7792 ), .Q ( new_AGEMA_signal_7793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3312 ( .C ( clk ), .D ( new_AGEMA_signal_7800 ), .Q ( new_AGEMA_signal_7801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3320 ( .C ( clk ), .D ( new_AGEMA_signal_7808 ), .Q ( new_AGEMA_signal_7809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3322 ( .C ( clk ), .D ( new_AGEMA_signal_7810 ), .Q ( new_AGEMA_signal_7811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3324 ( .C ( clk ), .D ( new_AGEMA_signal_7812 ), .Q ( new_AGEMA_signal_7813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3326 ( .C ( clk ), .D ( new_AGEMA_signal_7814 ), .Q ( new_AGEMA_signal_7815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3332 ( .C ( clk ), .D ( new_AGEMA_signal_7820 ), .Q ( new_AGEMA_signal_7821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3338 ( .C ( clk ), .D ( new_AGEMA_signal_7826 ), .Q ( new_AGEMA_signal_7827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3344 ( .C ( clk ), .D ( new_AGEMA_signal_7832 ), .Q ( new_AGEMA_signal_7833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3348 ( .C ( clk ), .D ( new_AGEMA_signal_7836 ), .Q ( new_AGEMA_signal_7837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3352 ( .C ( clk ), .D ( new_AGEMA_signal_7840 ), .Q ( new_AGEMA_signal_7841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3356 ( .C ( clk ), .D ( new_AGEMA_signal_7844 ), .Q ( new_AGEMA_signal_7845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3364 ( .C ( clk ), .D ( new_AGEMA_signal_7852 ), .Q ( new_AGEMA_signal_7853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3372 ( .C ( clk ), .D ( new_AGEMA_signal_7860 ), .Q ( new_AGEMA_signal_7861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3380 ( .C ( clk ), .D ( new_AGEMA_signal_7868 ), .Q ( new_AGEMA_signal_7869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3384 ( .C ( clk ), .D ( new_AGEMA_signal_7872 ), .Q ( new_AGEMA_signal_7873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3388 ( .C ( clk ), .D ( new_AGEMA_signal_7876 ), .Q ( new_AGEMA_signal_7877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3392 ( .C ( clk ), .D ( new_AGEMA_signal_7880 ), .Q ( new_AGEMA_signal_7881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3398 ( .C ( clk ), .D ( new_AGEMA_signal_7886 ), .Q ( new_AGEMA_signal_7887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3404 ( .C ( clk ), .D ( new_AGEMA_signal_7892 ), .Q ( new_AGEMA_signal_7893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3410 ( .C ( clk ), .D ( new_AGEMA_signal_7898 ), .Q ( new_AGEMA_signal_7899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3416 ( .C ( clk ), .D ( new_AGEMA_signal_7904 ), .Q ( new_AGEMA_signal_7905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3422 ( .C ( clk ), .D ( new_AGEMA_signal_7910 ), .Q ( new_AGEMA_signal_7911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3428 ( .C ( clk ), .D ( new_AGEMA_signal_7916 ), .Q ( new_AGEMA_signal_7917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3434 ( .C ( clk ), .D ( new_AGEMA_signal_7922 ), .Q ( new_AGEMA_signal_7923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3440 ( .C ( clk ), .D ( new_AGEMA_signal_7928 ), .Q ( new_AGEMA_signal_7929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3446 ( .C ( clk ), .D ( new_AGEMA_signal_7934 ), .Q ( new_AGEMA_signal_7935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3452 ( .C ( clk ), .D ( new_AGEMA_signal_7940 ), .Q ( new_AGEMA_signal_7941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3458 ( .C ( clk ), .D ( new_AGEMA_signal_7946 ), .Q ( new_AGEMA_signal_7947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3464 ( .C ( clk ), .D ( new_AGEMA_signal_7952 ), .Q ( new_AGEMA_signal_7953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3470 ( .C ( clk ), .D ( new_AGEMA_signal_7958 ), .Q ( new_AGEMA_signal_7959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3476 ( .C ( clk ), .D ( new_AGEMA_signal_7964 ), .Q ( new_AGEMA_signal_7965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3482 ( .C ( clk ), .D ( new_AGEMA_signal_7970 ), .Q ( new_AGEMA_signal_7971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3486 ( .C ( clk ), .D ( new_AGEMA_signal_7974 ), .Q ( new_AGEMA_signal_7975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3490 ( .C ( clk ), .D ( new_AGEMA_signal_7978 ), .Q ( new_AGEMA_signal_7979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3494 ( .C ( clk ), .D ( new_AGEMA_signal_7982 ), .Q ( new_AGEMA_signal_7983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3502 ( .C ( clk ), .D ( new_AGEMA_signal_7990 ), .Q ( new_AGEMA_signal_7991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3510 ( .C ( clk ), .D ( new_AGEMA_signal_7998 ), .Q ( new_AGEMA_signal_7999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3518 ( .C ( clk ), .D ( new_AGEMA_signal_8006 ), .Q ( new_AGEMA_signal_8007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3522 ( .C ( clk ), .D ( new_AGEMA_signal_8010 ), .Q ( new_AGEMA_signal_8011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3526 ( .C ( clk ), .D ( new_AGEMA_signal_8014 ), .Q ( new_AGEMA_signal_8015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3530 ( .C ( clk ), .D ( new_AGEMA_signal_8018 ), .Q ( new_AGEMA_signal_8019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3536 ( .C ( clk ), .D ( new_AGEMA_signal_8024 ), .Q ( new_AGEMA_signal_8025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3542 ( .C ( clk ), .D ( new_AGEMA_signal_8030 ), .Q ( new_AGEMA_signal_8031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3548 ( .C ( clk ), .D ( new_AGEMA_signal_8036 ), .Q ( new_AGEMA_signal_8037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3556 ( .C ( clk ), .D ( new_AGEMA_signal_8044 ), .Q ( new_AGEMA_signal_8045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3564 ( .C ( clk ), .D ( new_AGEMA_signal_8052 ), .Q ( new_AGEMA_signal_8053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3572 ( .C ( clk ), .D ( new_AGEMA_signal_8060 ), .Q ( new_AGEMA_signal_8061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3574 ( .C ( clk ), .D ( new_AGEMA_signal_8062 ), .Q ( new_AGEMA_signal_8063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3576 ( .C ( clk ), .D ( new_AGEMA_signal_8064 ), .Q ( new_AGEMA_signal_8065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3578 ( .C ( clk ), .D ( new_AGEMA_signal_8066 ), .Q ( new_AGEMA_signal_8067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3584 ( .C ( clk ), .D ( new_AGEMA_signal_8072 ), .Q ( new_AGEMA_signal_8073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3590 ( .C ( clk ), .D ( new_AGEMA_signal_8078 ), .Q ( new_AGEMA_signal_8079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3596 ( .C ( clk ), .D ( new_AGEMA_signal_8084 ), .Q ( new_AGEMA_signal_8085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3598 ( .C ( clk ), .D ( new_AGEMA_signal_8086 ), .Q ( new_AGEMA_signal_8087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3600 ( .C ( clk ), .D ( new_AGEMA_signal_8088 ), .Q ( new_AGEMA_signal_8089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3602 ( .C ( clk ), .D ( new_AGEMA_signal_8090 ), .Q ( new_AGEMA_signal_8091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3604 ( .C ( clk ), .D ( new_AGEMA_signal_8092 ), .Q ( new_AGEMA_signal_8093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3606 ( .C ( clk ), .D ( new_AGEMA_signal_8094 ), .Q ( new_AGEMA_signal_8095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3608 ( .C ( clk ), .D ( new_AGEMA_signal_8096 ), .Q ( new_AGEMA_signal_8097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3614 ( .C ( clk ), .D ( new_AGEMA_signal_8102 ), .Q ( new_AGEMA_signal_8103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3620 ( .C ( clk ), .D ( new_AGEMA_signal_8108 ), .Q ( new_AGEMA_signal_8109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3626 ( .C ( clk ), .D ( new_AGEMA_signal_8114 ), .Q ( new_AGEMA_signal_8115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3632 ( .C ( clk ), .D ( new_AGEMA_signal_8120 ), .Q ( new_AGEMA_signal_8121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3638 ( .C ( clk ), .D ( new_AGEMA_signal_8126 ), .Q ( new_AGEMA_signal_8127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3644 ( .C ( clk ), .D ( new_AGEMA_signal_8132 ), .Q ( new_AGEMA_signal_8133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3652 ( .C ( clk ), .D ( new_AGEMA_signal_8140 ), .Q ( new_AGEMA_signal_8141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3660 ( .C ( clk ), .D ( new_AGEMA_signal_8148 ), .Q ( new_AGEMA_signal_8149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3668 ( .C ( clk ), .D ( new_AGEMA_signal_8156 ), .Q ( new_AGEMA_signal_8157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3676 ( .C ( clk ), .D ( new_AGEMA_signal_8164 ), .Q ( new_AGEMA_signal_8165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3684 ( .C ( clk ), .D ( new_AGEMA_signal_8172 ), .Q ( new_AGEMA_signal_8173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3692 ( .C ( clk ), .D ( new_AGEMA_signal_8180 ), .Q ( new_AGEMA_signal_8181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3698 ( .C ( clk ), .D ( new_AGEMA_signal_8186 ), .Q ( new_AGEMA_signal_8187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3704 ( .C ( clk ), .D ( new_AGEMA_signal_8192 ), .Q ( new_AGEMA_signal_8193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3710 ( .C ( clk ), .D ( new_AGEMA_signal_8198 ), .Q ( new_AGEMA_signal_8199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3716 ( .C ( clk ), .D ( new_AGEMA_signal_8204 ), .Q ( new_AGEMA_signal_8205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3722 ( .C ( clk ), .D ( new_AGEMA_signal_8210 ), .Q ( new_AGEMA_signal_8211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3728 ( .C ( clk ), .D ( new_AGEMA_signal_8216 ), .Q ( new_AGEMA_signal_8217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3730 ( .C ( clk ), .D ( new_AGEMA_signal_8218 ), .Q ( new_AGEMA_signal_8219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3732 ( .C ( clk ), .D ( new_AGEMA_signal_8220 ), .Q ( new_AGEMA_signal_8221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3734 ( .C ( clk ), .D ( new_AGEMA_signal_8222 ), .Q ( new_AGEMA_signal_8223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3738 ( .C ( clk ), .D ( new_AGEMA_signal_8226 ), .Q ( new_AGEMA_signal_8227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3742 ( .C ( clk ), .D ( new_AGEMA_signal_8230 ), .Q ( new_AGEMA_signal_8231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3746 ( .C ( clk ), .D ( new_AGEMA_signal_8234 ), .Q ( new_AGEMA_signal_8235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3750 ( .C ( clk ), .D ( new_AGEMA_signal_8238 ), .Q ( new_AGEMA_signal_8239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3754 ( .C ( clk ), .D ( new_AGEMA_signal_8242 ), .Q ( new_AGEMA_signal_8243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3758 ( .C ( clk ), .D ( new_AGEMA_signal_8246 ), .Q ( new_AGEMA_signal_8247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3762 ( .C ( clk ), .D ( new_AGEMA_signal_8250 ), .Q ( new_AGEMA_signal_8251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3766 ( .C ( clk ), .D ( new_AGEMA_signal_8254 ), .Q ( new_AGEMA_signal_8255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3770 ( .C ( clk ), .D ( new_AGEMA_signal_8258 ), .Q ( new_AGEMA_signal_8259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3772 ( .C ( clk ), .D ( new_AGEMA_signal_8260 ), .Q ( new_AGEMA_signal_8261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3774 ( .C ( clk ), .D ( new_AGEMA_signal_8262 ), .Q ( new_AGEMA_signal_8263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3776 ( .C ( clk ), .D ( new_AGEMA_signal_8264 ), .Q ( new_AGEMA_signal_8265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3780 ( .C ( clk ), .D ( new_AGEMA_signal_8268 ), .Q ( new_AGEMA_signal_8269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3786 ( .C ( clk ), .D ( new_AGEMA_signal_8274 ), .Q ( new_AGEMA_signal_8275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3792 ( .C ( clk ), .D ( new_AGEMA_signal_8280 ), .Q ( new_AGEMA_signal_8281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3802 ( .C ( clk ), .D ( new_AGEMA_signal_8290 ), .Q ( new_AGEMA_signal_8291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3806 ( .C ( clk ), .D ( new_AGEMA_signal_8294 ), .Q ( new_AGEMA_signal_8295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3810 ( .C ( clk ), .D ( new_AGEMA_signal_8298 ), .Q ( new_AGEMA_signal_8299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3818 ( .C ( clk ), .D ( new_AGEMA_signal_8306 ), .Q ( new_AGEMA_signal_8307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3826 ( .C ( clk ), .D ( new_AGEMA_signal_8314 ), .Q ( new_AGEMA_signal_8315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3834 ( .C ( clk ), .D ( new_AGEMA_signal_8322 ), .Q ( new_AGEMA_signal_8323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3842 ( .C ( clk ), .D ( new_AGEMA_signal_8330 ), .Q ( new_AGEMA_signal_8331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3850 ( .C ( clk ), .D ( new_AGEMA_signal_8338 ), .Q ( new_AGEMA_signal_8339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3858 ( .C ( clk ), .D ( new_AGEMA_signal_8346 ), .Q ( new_AGEMA_signal_8347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3866 ( .C ( clk ), .D ( new_AGEMA_signal_8354 ), .Q ( new_AGEMA_signal_8355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3874 ( .C ( clk ), .D ( new_AGEMA_signal_8362 ), .Q ( new_AGEMA_signal_8363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3882 ( .C ( clk ), .D ( new_AGEMA_signal_8370 ), .Q ( new_AGEMA_signal_8371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3890 ( .C ( clk ), .D ( new_AGEMA_signal_8378 ), .Q ( new_AGEMA_signal_8379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3898 ( .C ( clk ), .D ( new_AGEMA_signal_8386 ), .Q ( new_AGEMA_signal_8387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3906 ( .C ( clk ), .D ( new_AGEMA_signal_8394 ), .Q ( new_AGEMA_signal_8395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3912 ( .C ( clk ), .D ( new_AGEMA_signal_8400 ), .Q ( new_AGEMA_signal_8401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3918 ( .C ( clk ), .D ( new_AGEMA_signal_8406 ), .Q ( new_AGEMA_signal_8407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3924 ( .C ( clk ), .D ( new_AGEMA_signal_8412 ), .Q ( new_AGEMA_signal_8413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3934 ( .C ( clk ), .D ( new_AGEMA_signal_8422 ), .Q ( new_AGEMA_signal_8423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3944 ( .C ( clk ), .D ( new_AGEMA_signal_8432 ), .Q ( new_AGEMA_signal_8433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3954 ( .C ( clk ), .D ( new_AGEMA_signal_8442 ), .Q ( new_AGEMA_signal_8443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3962 ( .C ( clk ), .D ( new_AGEMA_signal_8450 ), .Q ( new_AGEMA_signal_8451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3970 ( .C ( clk ), .D ( new_AGEMA_signal_8458 ), .Q ( new_AGEMA_signal_8459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3978 ( .C ( clk ), .D ( new_AGEMA_signal_8466 ), .Q ( new_AGEMA_signal_8467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3986 ( .C ( clk ), .D ( new_AGEMA_signal_8474 ), .Q ( new_AGEMA_signal_8475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3994 ( .C ( clk ), .D ( new_AGEMA_signal_8482 ), .Q ( new_AGEMA_signal_8483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4002 ( .C ( clk ), .D ( new_AGEMA_signal_8490 ), .Q ( new_AGEMA_signal_8491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4010 ( .C ( clk ), .D ( new_AGEMA_signal_8498 ), .Q ( new_AGEMA_signal_8499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4018 ( .C ( clk ), .D ( new_AGEMA_signal_8506 ), .Q ( new_AGEMA_signal_8507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4026 ( .C ( clk ), .D ( new_AGEMA_signal_8514 ), .Q ( new_AGEMA_signal_8515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4036 ( .C ( clk ), .D ( new_AGEMA_signal_8524 ), .Q ( new_AGEMA_signal_8525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4040 ( .C ( clk ), .D ( new_AGEMA_signal_8528 ), .Q ( new_AGEMA_signal_8529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4044 ( .C ( clk ), .D ( new_AGEMA_signal_8532 ), .Q ( new_AGEMA_signal_8533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4050 ( .C ( clk ), .D ( new_AGEMA_signal_8538 ), .Q ( new_AGEMA_signal_8539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4056 ( .C ( clk ), .D ( new_AGEMA_signal_8544 ), .Q ( new_AGEMA_signal_8545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4062 ( .C ( clk ), .D ( new_AGEMA_signal_8550 ), .Q ( new_AGEMA_signal_8551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4066 ( .C ( clk ), .D ( new_AGEMA_signal_8554 ), .Q ( new_AGEMA_signal_8555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4070 ( .C ( clk ), .D ( new_AGEMA_signal_8558 ), .Q ( new_AGEMA_signal_8559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4074 ( .C ( clk ), .D ( new_AGEMA_signal_8562 ), .Q ( new_AGEMA_signal_8563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4084 ( .C ( clk ), .D ( new_AGEMA_signal_8572 ), .Q ( new_AGEMA_signal_8573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4094 ( .C ( clk ), .D ( new_AGEMA_signal_8582 ), .Q ( new_AGEMA_signal_8583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4104 ( .C ( clk ), .D ( new_AGEMA_signal_8592 ), .Q ( new_AGEMA_signal_8593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4112 ( .C ( clk ), .D ( new_AGEMA_signal_8600 ), .Q ( new_AGEMA_signal_8601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4120 ( .C ( clk ), .D ( new_AGEMA_signal_8608 ), .Q ( new_AGEMA_signal_8609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4128 ( .C ( clk ), .D ( new_AGEMA_signal_8616 ), .Q ( new_AGEMA_signal_8617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4132 ( .C ( clk ), .D ( new_AGEMA_signal_8620 ), .Q ( new_AGEMA_signal_8621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4136 ( .C ( clk ), .D ( new_AGEMA_signal_8624 ), .Q ( new_AGEMA_signal_8625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4140 ( .C ( clk ), .D ( new_AGEMA_signal_8628 ), .Q ( new_AGEMA_signal_8629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4154 ( .C ( clk ), .D ( new_AGEMA_signal_8642 ), .Q ( new_AGEMA_signal_8643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4162 ( .C ( clk ), .D ( new_AGEMA_signal_8650 ), .Q ( new_AGEMA_signal_8651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4170 ( .C ( clk ), .D ( new_AGEMA_signal_8658 ), .Q ( new_AGEMA_signal_8659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4178 ( .C ( clk ), .D ( new_AGEMA_signal_8666 ), .Q ( new_AGEMA_signal_8667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4186 ( .C ( clk ), .D ( new_AGEMA_signal_8674 ), .Q ( new_AGEMA_signal_8675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4194 ( .C ( clk ), .D ( new_AGEMA_signal_8682 ), .Q ( new_AGEMA_signal_8683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4200 ( .C ( clk ), .D ( new_AGEMA_signal_8688 ), .Q ( new_AGEMA_signal_8689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4206 ( .C ( clk ), .D ( new_AGEMA_signal_8694 ), .Q ( new_AGEMA_signal_8695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4212 ( .C ( clk ), .D ( new_AGEMA_signal_8700 ), .Q ( new_AGEMA_signal_8701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4216 ( .C ( clk ), .D ( new_AGEMA_signal_8704 ), .Q ( new_AGEMA_signal_8705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4220 ( .C ( clk ), .D ( new_AGEMA_signal_8708 ), .Q ( new_AGEMA_signal_8709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4224 ( .C ( clk ), .D ( new_AGEMA_signal_8712 ), .Q ( new_AGEMA_signal_8713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4232 ( .C ( clk ), .D ( new_AGEMA_signal_8720 ), .Q ( new_AGEMA_signal_8721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4240 ( .C ( clk ), .D ( new_AGEMA_signal_8728 ), .Q ( new_AGEMA_signal_8729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4248 ( .C ( clk ), .D ( new_AGEMA_signal_8736 ), .Q ( new_AGEMA_signal_8737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4258 ( .C ( clk ), .D ( new_AGEMA_signal_8746 ), .Q ( new_AGEMA_signal_8747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4264 ( .C ( clk ), .D ( new_AGEMA_signal_8752 ), .Q ( new_AGEMA_signal_8753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4270 ( .C ( clk ), .D ( new_AGEMA_signal_8758 ), .Q ( new_AGEMA_signal_8759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4276 ( .C ( clk ), .D ( new_AGEMA_signal_8764 ), .Q ( new_AGEMA_signal_8765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4282 ( .C ( clk ), .D ( new_AGEMA_signal_8770 ), .Q ( new_AGEMA_signal_8771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4288 ( .C ( clk ), .D ( new_AGEMA_signal_8776 ), .Q ( new_AGEMA_signal_8777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4294 ( .C ( clk ), .D ( new_AGEMA_signal_8782 ), .Q ( new_AGEMA_signal_8783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4300 ( .C ( clk ), .D ( new_AGEMA_signal_8788 ), .Q ( new_AGEMA_signal_8789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4306 ( .C ( clk ), .D ( new_AGEMA_signal_8794 ), .Q ( new_AGEMA_signal_8795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4326 ( .C ( clk ), .D ( new_AGEMA_signal_8814 ), .Q ( new_AGEMA_signal_8815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4334 ( .C ( clk ), .D ( new_AGEMA_signal_8822 ), .Q ( new_AGEMA_signal_8823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4342 ( .C ( clk ), .D ( new_AGEMA_signal_8830 ), .Q ( new_AGEMA_signal_8831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4348 ( .C ( clk ), .D ( new_AGEMA_signal_8836 ), .Q ( new_AGEMA_signal_8837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4354 ( .C ( clk ), .D ( new_AGEMA_signal_8842 ), .Q ( new_AGEMA_signal_8843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4360 ( .C ( clk ), .D ( new_AGEMA_signal_8848 ), .Q ( new_AGEMA_signal_8849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4380 ( .C ( clk ), .D ( new_AGEMA_signal_8868 ), .Q ( new_AGEMA_signal_8869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4388 ( .C ( clk ), .D ( new_AGEMA_signal_8876 ), .Q ( new_AGEMA_signal_8877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4396 ( .C ( clk ), .D ( new_AGEMA_signal_8884 ), .Q ( new_AGEMA_signal_8885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4404 ( .C ( clk ), .D ( new_AGEMA_signal_8892 ), .Q ( new_AGEMA_signal_8893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4412 ( .C ( clk ), .D ( new_AGEMA_signal_8900 ), .Q ( new_AGEMA_signal_8901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4420 ( .C ( clk ), .D ( new_AGEMA_signal_8908 ), .Q ( new_AGEMA_signal_8909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4430 ( .C ( clk ), .D ( new_AGEMA_signal_8918 ), .Q ( new_AGEMA_signal_8919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4440 ( .C ( clk ), .D ( new_AGEMA_signal_8928 ), .Q ( new_AGEMA_signal_8929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4450 ( .C ( clk ), .D ( new_AGEMA_signal_8938 ), .Q ( new_AGEMA_signal_8939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4458 ( .C ( clk ), .D ( new_AGEMA_signal_8946 ), .Q ( new_AGEMA_signal_8947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4466 ( .C ( clk ), .D ( new_AGEMA_signal_8954 ), .Q ( new_AGEMA_signal_8955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4474 ( .C ( clk ), .D ( new_AGEMA_signal_8962 ), .Q ( new_AGEMA_signal_8963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4480 ( .C ( clk ), .D ( new_AGEMA_signal_8968 ), .Q ( new_AGEMA_signal_8969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4486 ( .C ( clk ), .D ( new_AGEMA_signal_8974 ), .Q ( new_AGEMA_signal_8975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4492 ( .C ( clk ), .D ( new_AGEMA_signal_8980 ), .Q ( new_AGEMA_signal_8981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4510 ( .C ( clk ), .D ( new_AGEMA_signal_8998 ), .Q ( new_AGEMA_signal_8999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4516 ( .C ( clk ), .D ( new_AGEMA_signal_9004 ), .Q ( new_AGEMA_signal_9005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4522 ( .C ( clk ), .D ( new_AGEMA_signal_9010 ), .Q ( new_AGEMA_signal_9011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4530 ( .C ( clk ), .D ( new_AGEMA_signal_9018 ), .Q ( new_AGEMA_signal_9019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4538 ( .C ( clk ), .D ( new_AGEMA_signal_9026 ), .Q ( new_AGEMA_signal_9027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4546 ( .C ( clk ), .D ( new_AGEMA_signal_9034 ), .Q ( new_AGEMA_signal_9035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4552 ( .C ( clk ), .D ( new_AGEMA_signal_9040 ), .Q ( new_AGEMA_signal_9041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4558 ( .C ( clk ), .D ( new_AGEMA_signal_9046 ), .Q ( new_AGEMA_signal_9047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4564 ( .C ( clk ), .D ( new_AGEMA_signal_9052 ), .Q ( new_AGEMA_signal_9053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4578 ( .C ( clk ), .D ( new_AGEMA_signal_9066 ), .Q ( new_AGEMA_signal_9067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4586 ( .C ( clk ), .D ( new_AGEMA_signal_9074 ), .Q ( new_AGEMA_signal_9075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4594 ( .C ( clk ), .D ( new_AGEMA_signal_9082 ), .Q ( new_AGEMA_signal_9083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4612 ( .C ( clk ), .D ( new_AGEMA_signal_9100 ), .Q ( new_AGEMA_signal_9101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4618 ( .C ( clk ), .D ( new_AGEMA_signal_9106 ), .Q ( new_AGEMA_signal_9107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4624 ( .C ( clk ), .D ( new_AGEMA_signal_9112 ), .Q ( new_AGEMA_signal_9113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4630 ( .C ( clk ), .D ( new_AGEMA_signal_9118 ), .Q ( new_AGEMA_signal_9119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4636 ( .C ( clk ), .D ( new_AGEMA_signal_9124 ), .Q ( new_AGEMA_signal_9125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4642 ( .C ( clk ), .D ( new_AGEMA_signal_9130 ), .Q ( new_AGEMA_signal_9131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4710 ( .C ( clk ), .D ( new_AGEMA_signal_9198 ), .Q ( new_AGEMA_signal_9199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4720 ( .C ( clk ), .D ( new_AGEMA_signal_9208 ), .Q ( new_AGEMA_signal_9209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4730 ( .C ( clk ), .D ( new_AGEMA_signal_9218 ), .Q ( new_AGEMA_signal_9219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4798 ( .C ( clk ), .D ( new_AGEMA_signal_9286 ), .Q ( new_AGEMA_signal_9287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4806 ( .C ( clk ), .D ( new_AGEMA_signal_9294 ), .Q ( new_AGEMA_signal_9295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4814 ( .C ( clk ), .D ( new_AGEMA_signal_9302 ), .Q ( new_AGEMA_signal_9303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4840 ( .C ( clk ), .D ( new_AGEMA_signal_9328 ), .Q ( new_AGEMA_signal_9329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4848 ( .C ( clk ), .D ( new_AGEMA_signal_9336 ), .Q ( new_AGEMA_signal_9337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4856 ( .C ( clk ), .D ( new_AGEMA_signal_9344 ), .Q ( new_AGEMA_signal_9345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4864 ( .C ( clk ), .D ( new_AGEMA_signal_9352 ), .Q ( new_AGEMA_signal_9353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4872 ( .C ( clk ), .D ( new_AGEMA_signal_9360 ), .Q ( new_AGEMA_signal_9361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4880 ( .C ( clk ), .D ( new_AGEMA_signal_9368 ), .Q ( new_AGEMA_signal_9369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4918 ( .C ( clk ), .D ( new_AGEMA_signal_9406 ), .Q ( new_AGEMA_signal_9407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4926 ( .C ( clk ), .D ( new_AGEMA_signal_9414 ), .Q ( new_AGEMA_signal_9415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4934 ( .C ( clk ), .D ( new_AGEMA_signal_9422 ), .Q ( new_AGEMA_signal_9423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4980 ( .C ( clk ), .D ( new_AGEMA_signal_9468 ), .Q ( new_AGEMA_signal_9469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4992 ( .C ( clk ), .D ( new_AGEMA_signal_9480 ), .Q ( new_AGEMA_signal_9481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5004 ( .C ( clk ), .D ( new_AGEMA_signal_9492 ), .Q ( new_AGEMA_signal_9493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5018 ( .C ( clk ), .D ( new_AGEMA_signal_9506 ), .Q ( new_AGEMA_signal_9507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5032 ( .C ( clk ), .D ( new_AGEMA_signal_9520 ), .Q ( new_AGEMA_signal_9521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5046 ( .C ( clk ), .D ( new_AGEMA_signal_9534 ), .Q ( new_AGEMA_signal_9535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5084 ( .C ( clk ), .D ( new_AGEMA_signal_9572 ), .Q ( new_AGEMA_signal_9573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5098 ( .C ( clk ), .D ( new_AGEMA_signal_9586 ), .Q ( new_AGEMA_signal_9587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5112 ( .C ( clk ), .D ( new_AGEMA_signal_9600 ), .Q ( new_AGEMA_signal_9601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5192 ( .C ( clk ), .D ( new_AGEMA_signal_9680 ), .Q ( new_AGEMA_signal_9681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5208 ( .C ( clk ), .D ( new_AGEMA_signal_9696 ), .Q ( new_AGEMA_signal_9697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5224 ( .C ( clk ), .D ( new_AGEMA_signal_9712 ), .Q ( new_AGEMA_signal_9713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5258 ( .C ( clk ), .D ( new_AGEMA_signal_9746 ), .Q ( new_AGEMA_signal_9747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5274 ( .C ( clk ), .D ( new_AGEMA_signal_9762 ), .Q ( new_AGEMA_signal_9763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5290 ( .C ( clk ), .D ( new_AGEMA_signal_9778 ), .Q ( new_AGEMA_signal_9779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5406 ( .C ( clk ), .D ( new_AGEMA_signal_9894 ), .Q ( new_AGEMA_signal_9895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5422 ( .C ( clk ), .D ( new_AGEMA_signal_9910 ), .Q ( new_AGEMA_signal_9911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5438 ( .C ( clk ), .D ( new_AGEMA_signal_9926 ), .Q ( new_AGEMA_signal_9927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5486 ( .C ( clk ), .D ( new_AGEMA_signal_9974 ), .Q ( new_AGEMA_signal_9975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5504 ( .C ( clk ), .D ( new_AGEMA_signal_9992 ), .Q ( new_AGEMA_signal_9993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5522 ( .C ( clk ), .D ( new_AGEMA_signal_10010 ), .Q ( new_AGEMA_signal_10011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5636 ( .C ( clk ), .D ( new_AGEMA_signal_10124 ), .Q ( new_AGEMA_signal_10125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5656 ( .C ( clk ), .D ( new_AGEMA_signal_10144 ), .Q ( new_AGEMA_signal_10145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5676 ( .C ( clk ), .D ( new_AGEMA_signal_10164 ), .Q ( new_AGEMA_signal_10165 ) ) ;

    /* cells in depth 13 */
    buf_clk new_AGEMA_reg_buffer_3781 ( .C ( clk ), .D ( new_AGEMA_signal_8269 ), .Q ( new_AGEMA_signal_8270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3787 ( .C ( clk ), .D ( new_AGEMA_signal_8275 ), .Q ( new_AGEMA_signal_8276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3793 ( .C ( clk ), .D ( new_AGEMA_signal_8281 ), .Q ( new_AGEMA_signal_8282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3795 ( .C ( clk ), .D ( new_AGEMA_signal_8227 ), .Q ( new_AGEMA_signal_8284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3797 ( .C ( clk ), .D ( new_AGEMA_signal_8231 ), .Q ( new_AGEMA_signal_8286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3799 ( .C ( clk ), .D ( new_AGEMA_signal_8235 ), .Q ( new_AGEMA_signal_8288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3803 ( .C ( clk ), .D ( new_AGEMA_signal_8291 ), .Q ( new_AGEMA_signal_8292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3807 ( .C ( clk ), .D ( new_AGEMA_signal_8295 ), .Q ( new_AGEMA_signal_8296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3811 ( .C ( clk ), .D ( new_AGEMA_signal_8299 ), .Q ( new_AGEMA_signal_8300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3819 ( .C ( clk ), .D ( new_AGEMA_signal_8307 ), .Q ( new_AGEMA_signal_8308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3827 ( .C ( clk ), .D ( new_AGEMA_signal_8315 ), .Q ( new_AGEMA_signal_8316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3835 ( .C ( clk ), .D ( new_AGEMA_signal_8323 ), .Q ( new_AGEMA_signal_8324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3843 ( .C ( clk ), .D ( new_AGEMA_signal_8331 ), .Q ( new_AGEMA_signal_8332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3851 ( .C ( clk ), .D ( new_AGEMA_signal_8339 ), .Q ( new_AGEMA_signal_8340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3859 ( .C ( clk ), .D ( new_AGEMA_signal_8347 ), .Q ( new_AGEMA_signal_8348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3867 ( .C ( clk ), .D ( new_AGEMA_signal_8355 ), .Q ( new_AGEMA_signal_8356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3875 ( .C ( clk ), .D ( new_AGEMA_signal_8363 ), .Q ( new_AGEMA_signal_8364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3883 ( .C ( clk ), .D ( new_AGEMA_signal_8371 ), .Q ( new_AGEMA_signal_8372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3891 ( .C ( clk ), .D ( new_AGEMA_signal_8379 ), .Q ( new_AGEMA_signal_8380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3899 ( .C ( clk ), .D ( new_AGEMA_signal_8387 ), .Q ( new_AGEMA_signal_8388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3907 ( .C ( clk ), .D ( new_AGEMA_signal_8395 ), .Q ( new_AGEMA_signal_8396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3913 ( .C ( clk ), .D ( new_AGEMA_signal_8401 ), .Q ( new_AGEMA_signal_8402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3919 ( .C ( clk ), .D ( new_AGEMA_signal_8407 ), .Q ( new_AGEMA_signal_8408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3925 ( .C ( clk ), .D ( new_AGEMA_signal_8413 ), .Q ( new_AGEMA_signal_8414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3935 ( .C ( clk ), .D ( new_AGEMA_signal_8423 ), .Q ( new_AGEMA_signal_8424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3945 ( .C ( clk ), .D ( new_AGEMA_signal_8433 ), .Q ( new_AGEMA_signal_8434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3955 ( .C ( clk ), .D ( new_AGEMA_signal_8443 ), .Q ( new_AGEMA_signal_8444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3963 ( .C ( clk ), .D ( new_AGEMA_signal_8451 ), .Q ( new_AGEMA_signal_8452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3971 ( .C ( clk ), .D ( new_AGEMA_signal_8459 ), .Q ( new_AGEMA_signal_8460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3979 ( .C ( clk ), .D ( new_AGEMA_signal_8467 ), .Q ( new_AGEMA_signal_8468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3987 ( .C ( clk ), .D ( new_AGEMA_signal_8475 ), .Q ( new_AGEMA_signal_8476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3995 ( .C ( clk ), .D ( new_AGEMA_signal_8483 ), .Q ( new_AGEMA_signal_8484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4003 ( .C ( clk ), .D ( new_AGEMA_signal_8491 ), .Q ( new_AGEMA_signal_8492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4011 ( .C ( clk ), .D ( new_AGEMA_signal_8499 ), .Q ( new_AGEMA_signal_8500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4019 ( .C ( clk ), .D ( new_AGEMA_signal_8507 ), .Q ( new_AGEMA_signal_8508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4027 ( .C ( clk ), .D ( new_AGEMA_signal_8515 ), .Q ( new_AGEMA_signal_8516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4029 ( .C ( clk ), .D ( new_AGEMA_signal_7811 ), .Q ( new_AGEMA_signal_8518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4031 ( .C ( clk ), .D ( new_AGEMA_signal_7813 ), .Q ( new_AGEMA_signal_8520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4033 ( .C ( clk ), .D ( new_AGEMA_signal_7815 ), .Q ( new_AGEMA_signal_8522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4037 ( .C ( clk ), .D ( new_AGEMA_signal_8525 ), .Q ( new_AGEMA_signal_8526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4041 ( .C ( clk ), .D ( new_AGEMA_signal_8529 ), .Q ( new_AGEMA_signal_8530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4045 ( .C ( clk ), .D ( new_AGEMA_signal_8533 ), .Q ( new_AGEMA_signal_8534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4051 ( .C ( clk ), .D ( new_AGEMA_signal_8539 ), .Q ( new_AGEMA_signal_8540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4057 ( .C ( clk ), .D ( new_AGEMA_signal_8545 ), .Q ( new_AGEMA_signal_8546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4063 ( .C ( clk ), .D ( new_AGEMA_signal_8551 ), .Q ( new_AGEMA_signal_8552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4067 ( .C ( clk ), .D ( new_AGEMA_signal_8555 ), .Q ( new_AGEMA_signal_8556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4071 ( .C ( clk ), .D ( new_AGEMA_signal_8559 ), .Q ( new_AGEMA_signal_8560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4075 ( .C ( clk ), .D ( new_AGEMA_signal_8563 ), .Q ( new_AGEMA_signal_8564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4085 ( .C ( clk ), .D ( new_AGEMA_signal_8573 ), .Q ( new_AGEMA_signal_8574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4095 ( .C ( clk ), .D ( new_AGEMA_signal_8583 ), .Q ( new_AGEMA_signal_8584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4105 ( .C ( clk ), .D ( new_AGEMA_signal_8593 ), .Q ( new_AGEMA_signal_8594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4113 ( .C ( clk ), .D ( new_AGEMA_signal_8601 ), .Q ( new_AGEMA_signal_8602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4121 ( .C ( clk ), .D ( new_AGEMA_signal_8609 ), .Q ( new_AGEMA_signal_8610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4129 ( .C ( clk ), .D ( new_AGEMA_signal_8617 ), .Q ( new_AGEMA_signal_8618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4133 ( .C ( clk ), .D ( new_AGEMA_signal_8621 ), .Q ( new_AGEMA_signal_8622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4137 ( .C ( clk ), .D ( new_AGEMA_signal_8625 ), .Q ( new_AGEMA_signal_8626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4141 ( .C ( clk ), .D ( new_AGEMA_signal_8629 ), .Q ( new_AGEMA_signal_8630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4143 ( .C ( clk ), .D ( n2509 ), .Q ( new_AGEMA_signal_8632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4145 ( .C ( clk ), .D ( new_AGEMA_signal_2572 ), .Q ( new_AGEMA_signal_8634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4147 ( .C ( clk ), .D ( new_AGEMA_signal_2573 ), .Q ( new_AGEMA_signal_8636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4155 ( .C ( clk ), .D ( new_AGEMA_signal_8643 ), .Q ( new_AGEMA_signal_8644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4163 ( .C ( clk ), .D ( new_AGEMA_signal_8651 ), .Q ( new_AGEMA_signal_8652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4171 ( .C ( clk ), .D ( new_AGEMA_signal_8659 ), .Q ( new_AGEMA_signal_8660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4179 ( .C ( clk ), .D ( new_AGEMA_signal_8667 ), .Q ( new_AGEMA_signal_8668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4187 ( .C ( clk ), .D ( new_AGEMA_signal_8675 ), .Q ( new_AGEMA_signal_8676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4195 ( .C ( clk ), .D ( new_AGEMA_signal_8683 ), .Q ( new_AGEMA_signal_8684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4201 ( .C ( clk ), .D ( new_AGEMA_signal_8689 ), .Q ( new_AGEMA_signal_8690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4207 ( .C ( clk ), .D ( new_AGEMA_signal_8695 ), .Q ( new_AGEMA_signal_8696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4213 ( .C ( clk ), .D ( new_AGEMA_signal_8701 ), .Q ( new_AGEMA_signal_8702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4217 ( .C ( clk ), .D ( new_AGEMA_signal_8705 ), .Q ( new_AGEMA_signal_8706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4221 ( .C ( clk ), .D ( new_AGEMA_signal_8709 ), .Q ( new_AGEMA_signal_8710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4225 ( .C ( clk ), .D ( new_AGEMA_signal_8713 ), .Q ( new_AGEMA_signal_8714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4233 ( .C ( clk ), .D ( new_AGEMA_signal_8721 ), .Q ( new_AGEMA_signal_8722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4241 ( .C ( clk ), .D ( new_AGEMA_signal_8729 ), .Q ( new_AGEMA_signal_8730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4249 ( .C ( clk ), .D ( new_AGEMA_signal_8737 ), .Q ( new_AGEMA_signal_8738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4251 ( .C ( clk ), .D ( n2802 ), .Q ( new_AGEMA_signal_8740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4253 ( .C ( clk ), .D ( new_AGEMA_signal_2504 ), .Q ( new_AGEMA_signal_8742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4255 ( .C ( clk ), .D ( new_AGEMA_signal_2505 ), .Q ( new_AGEMA_signal_8744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4259 ( .C ( clk ), .D ( new_AGEMA_signal_8747 ), .Q ( new_AGEMA_signal_8748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4265 ( .C ( clk ), .D ( new_AGEMA_signal_8753 ), .Q ( new_AGEMA_signal_8754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4271 ( .C ( clk ), .D ( new_AGEMA_signal_8759 ), .Q ( new_AGEMA_signal_8760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4277 ( .C ( clk ), .D ( new_AGEMA_signal_8765 ), .Q ( new_AGEMA_signal_8766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4283 ( .C ( clk ), .D ( new_AGEMA_signal_8771 ), .Q ( new_AGEMA_signal_8772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4289 ( .C ( clk ), .D ( new_AGEMA_signal_8777 ), .Q ( new_AGEMA_signal_8778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4295 ( .C ( clk ), .D ( new_AGEMA_signal_8783 ), .Q ( new_AGEMA_signal_8784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4301 ( .C ( clk ), .D ( new_AGEMA_signal_8789 ), .Q ( new_AGEMA_signal_8790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4307 ( .C ( clk ), .D ( new_AGEMA_signal_8795 ), .Q ( new_AGEMA_signal_8796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4311 ( .C ( clk ), .D ( new_AGEMA_signal_8261 ), .Q ( new_AGEMA_signal_8800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4315 ( .C ( clk ), .D ( new_AGEMA_signal_8263 ), .Q ( new_AGEMA_signal_8804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4319 ( .C ( clk ), .D ( new_AGEMA_signal_8265 ), .Q ( new_AGEMA_signal_8808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4327 ( .C ( clk ), .D ( new_AGEMA_signal_8815 ), .Q ( new_AGEMA_signal_8816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4335 ( .C ( clk ), .D ( new_AGEMA_signal_8823 ), .Q ( new_AGEMA_signal_8824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4343 ( .C ( clk ), .D ( new_AGEMA_signal_8831 ), .Q ( new_AGEMA_signal_8832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4349 ( .C ( clk ), .D ( new_AGEMA_signal_8837 ), .Q ( new_AGEMA_signal_8838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4355 ( .C ( clk ), .D ( new_AGEMA_signal_8843 ), .Q ( new_AGEMA_signal_8844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4361 ( .C ( clk ), .D ( new_AGEMA_signal_8849 ), .Q ( new_AGEMA_signal_8850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4365 ( .C ( clk ), .D ( n2072 ), .Q ( new_AGEMA_signal_8854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4369 ( .C ( clk ), .D ( new_AGEMA_signal_2410 ), .Q ( new_AGEMA_signal_8858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4373 ( .C ( clk ), .D ( new_AGEMA_signal_2411 ), .Q ( new_AGEMA_signal_8862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4381 ( .C ( clk ), .D ( new_AGEMA_signal_8869 ), .Q ( new_AGEMA_signal_8870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4389 ( .C ( clk ), .D ( new_AGEMA_signal_8877 ), .Q ( new_AGEMA_signal_8878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4397 ( .C ( clk ), .D ( new_AGEMA_signal_8885 ), .Q ( new_AGEMA_signal_8886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4405 ( .C ( clk ), .D ( new_AGEMA_signal_8893 ), .Q ( new_AGEMA_signal_8894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4413 ( .C ( clk ), .D ( new_AGEMA_signal_8901 ), .Q ( new_AGEMA_signal_8902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4421 ( .C ( clk ), .D ( new_AGEMA_signal_8909 ), .Q ( new_AGEMA_signal_8910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4431 ( .C ( clk ), .D ( new_AGEMA_signal_8919 ), .Q ( new_AGEMA_signal_8920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4441 ( .C ( clk ), .D ( new_AGEMA_signal_8929 ), .Q ( new_AGEMA_signal_8930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4451 ( .C ( clk ), .D ( new_AGEMA_signal_8939 ), .Q ( new_AGEMA_signal_8940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4459 ( .C ( clk ), .D ( new_AGEMA_signal_8947 ), .Q ( new_AGEMA_signal_8948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4467 ( .C ( clk ), .D ( new_AGEMA_signal_8955 ), .Q ( new_AGEMA_signal_8956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4475 ( .C ( clk ), .D ( new_AGEMA_signal_8963 ), .Q ( new_AGEMA_signal_8964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4481 ( .C ( clk ), .D ( new_AGEMA_signal_8969 ), .Q ( new_AGEMA_signal_8970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4487 ( .C ( clk ), .D ( new_AGEMA_signal_8975 ), .Q ( new_AGEMA_signal_8976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4493 ( .C ( clk ), .D ( new_AGEMA_signal_8981 ), .Q ( new_AGEMA_signal_8982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4497 ( .C ( clk ), .D ( n2276 ), .Q ( new_AGEMA_signal_8986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4501 ( .C ( clk ), .D ( new_AGEMA_signal_2442 ), .Q ( new_AGEMA_signal_8990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4505 ( .C ( clk ), .D ( new_AGEMA_signal_2443 ), .Q ( new_AGEMA_signal_8994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4511 ( .C ( clk ), .D ( new_AGEMA_signal_8999 ), .Q ( new_AGEMA_signal_9000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4517 ( .C ( clk ), .D ( new_AGEMA_signal_9005 ), .Q ( new_AGEMA_signal_9006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4523 ( .C ( clk ), .D ( new_AGEMA_signal_9011 ), .Q ( new_AGEMA_signal_9012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4531 ( .C ( clk ), .D ( new_AGEMA_signal_9019 ), .Q ( new_AGEMA_signal_9020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4539 ( .C ( clk ), .D ( new_AGEMA_signal_9027 ), .Q ( new_AGEMA_signal_9028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4547 ( .C ( clk ), .D ( new_AGEMA_signal_9035 ), .Q ( new_AGEMA_signal_9036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4553 ( .C ( clk ), .D ( new_AGEMA_signal_9041 ), .Q ( new_AGEMA_signal_9042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4559 ( .C ( clk ), .D ( new_AGEMA_signal_9047 ), .Q ( new_AGEMA_signal_9048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4565 ( .C ( clk ), .D ( new_AGEMA_signal_9053 ), .Q ( new_AGEMA_signal_9054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4579 ( .C ( clk ), .D ( new_AGEMA_signal_9067 ), .Q ( new_AGEMA_signal_9068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4587 ( .C ( clk ), .D ( new_AGEMA_signal_9075 ), .Q ( new_AGEMA_signal_9076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4595 ( .C ( clk ), .D ( new_AGEMA_signal_9083 ), .Q ( new_AGEMA_signal_9084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4599 ( .C ( clk ), .D ( n2622 ), .Q ( new_AGEMA_signal_9088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4603 ( .C ( clk ), .D ( new_AGEMA_signal_2488 ), .Q ( new_AGEMA_signal_9092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4607 ( .C ( clk ), .D ( new_AGEMA_signal_2489 ), .Q ( new_AGEMA_signal_9096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4613 ( .C ( clk ), .D ( new_AGEMA_signal_9101 ), .Q ( new_AGEMA_signal_9102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4619 ( .C ( clk ), .D ( new_AGEMA_signal_9107 ), .Q ( new_AGEMA_signal_9108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4625 ( .C ( clk ), .D ( new_AGEMA_signal_9113 ), .Q ( new_AGEMA_signal_9114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4631 ( .C ( clk ), .D ( new_AGEMA_signal_9119 ), .Q ( new_AGEMA_signal_9120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4637 ( .C ( clk ), .D ( new_AGEMA_signal_9125 ), .Q ( new_AGEMA_signal_9126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4643 ( .C ( clk ), .D ( new_AGEMA_signal_9131 ), .Q ( new_AGEMA_signal_9132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4647 ( .C ( clk ), .D ( n2804 ), .Q ( new_AGEMA_signal_9136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4651 ( .C ( clk ), .D ( new_AGEMA_signal_2502 ), .Q ( new_AGEMA_signal_9140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4655 ( .C ( clk ), .D ( new_AGEMA_signal_2503 ), .Q ( new_AGEMA_signal_9144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4659 ( .C ( clk ), .D ( n1990 ), .Q ( new_AGEMA_signal_9148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4665 ( .C ( clk ), .D ( new_AGEMA_signal_2238 ), .Q ( new_AGEMA_signal_9154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4671 ( .C ( clk ), .D ( new_AGEMA_signal_2239 ), .Q ( new_AGEMA_signal_9160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4689 ( .C ( clk ), .D ( n2078 ), .Q ( new_AGEMA_signal_9178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4695 ( .C ( clk ), .D ( new_AGEMA_signal_2414 ), .Q ( new_AGEMA_signal_9184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4701 ( .C ( clk ), .D ( new_AGEMA_signal_2415 ), .Q ( new_AGEMA_signal_9190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4711 ( .C ( clk ), .D ( new_AGEMA_signal_9199 ), .Q ( new_AGEMA_signal_9200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4721 ( .C ( clk ), .D ( new_AGEMA_signal_9209 ), .Q ( new_AGEMA_signal_9210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4731 ( .C ( clk ), .D ( new_AGEMA_signal_9219 ), .Q ( new_AGEMA_signal_9220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4737 ( .C ( clk ), .D ( n2128 ), .Q ( new_AGEMA_signal_9226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4743 ( .C ( clk ), .D ( new_AGEMA_signal_2528 ), .Q ( new_AGEMA_signal_9232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4749 ( .C ( clk ), .D ( new_AGEMA_signal_2529 ), .Q ( new_AGEMA_signal_9238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4755 ( .C ( clk ), .D ( n2148 ), .Q ( new_AGEMA_signal_9244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4761 ( .C ( clk ), .D ( new_AGEMA_signal_2274 ), .Q ( new_AGEMA_signal_9250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4767 ( .C ( clk ), .D ( new_AGEMA_signal_2275 ), .Q ( new_AGEMA_signal_9256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4799 ( .C ( clk ), .D ( new_AGEMA_signal_9287 ), .Q ( new_AGEMA_signal_9288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4807 ( .C ( clk ), .D ( new_AGEMA_signal_9295 ), .Q ( new_AGEMA_signal_9296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4815 ( .C ( clk ), .D ( new_AGEMA_signal_9303 ), .Q ( new_AGEMA_signal_9304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4821 ( .C ( clk ), .D ( n2306 ), .Q ( new_AGEMA_signal_9310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4827 ( .C ( clk ), .D ( new_AGEMA_signal_2300 ), .Q ( new_AGEMA_signal_9316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4833 ( .C ( clk ), .D ( new_AGEMA_signal_2301 ), .Q ( new_AGEMA_signal_9322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4841 ( .C ( clk ), .D ( new_AGEMA_signal_9329 ), .Q ( new_AGEMA_signal_9330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4849 ( .C ( clk ), .D ( new_AGEMA_signal_9337 ), .Q ( new_AGEMA_signal_9338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4857 ( .C ( clk ), .D ( new_AGEMA_signal_9345 ), .Q ( new_AGEMA_signal_9346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4865 ( .C ( clk ), .D ( new_AGEMA_signal_9353 ), .Q ( new_AGEMA_signal_9354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4873 ( .C ( clk ), .D ( new_AGEMA_signal_9361 ), .Q ( new_AGEMA_signal_9362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4881 ( .C ( clk ), .D ( new_AGEMA_signal_9369 ), .Q ( new_AGEMA_signal_9370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4919 ( .C ( clk ), .D ( new_AGEMA_signal_9407 ), .Q ( new_AGEMA_signal_9408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4927 ( .C ( clk ), .D ( new_AGEMA_signal_9415 ), .Q ( new_AGEMA_signal_9416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4935 ( .C ( clk ), .D ( new_AGEMA_signal_9423 ), .Q ( new_AGEMA_signal_9424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4953 ( .C ( clk ), .D ( n1999 ), .Q ( new_AGEMA_signal_9442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4961 ( .C ( clk ), .D ( new_AGEMA_signal_2400 ), .Q ( new_AGEMA_signal_9450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4969 ( .C ( clk ), .D ( new_AGEMA_signal_2401 ), .Q ( new_AGEMA_signal_9458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4981 ( .C ( clk ), .D ( new_AGEMA_signal_9469 ), .Q ( new_AGEMA_signal_9470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4993 ( .C ( clk ), .D ( new_AGEMA_signal_9481 ), .Q ( new_AGEMA_signal_9482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5005 ( .C ( clk ), .D ( new_AGEMA_signal_9493 ), .Q ( new_AGEMA_signal_9494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5019 ( .C ( clk ), .D ( new_AGEMA_signal_9507 ), .Q ( new_AGEMA_signal_9508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5033 ( .C ( clk ), .D ( new_AGEMA_signal_9521 ), .Q ( new_AGEMA_signal_9522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5047 ( .C ( clk ), .D ( new_AGEMA_signal_9535 ), .Q ( new_AGEMA_signal_9536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5055 ( .C ( clk ), .D ( n2205 ), .Q ( new_AGEMA_signal_9544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5063 ( .C ( clk ), .D ( new_AGEMA_signal_2540 ), .Q ( new_AGEMA_signal_9552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5071 ( .C ( clk ), .D ( new_AGEMA_signal_2541 ), .Q ( new_AGEMA_signal_9560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5085 ( .C ( clk ), .D ( new_AGEMA_signal_9573 ), .Q ( new_AGEMA_signal_9574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5099 ( .C ( clk ), .D ( new_AGEMA_signal_9587 ), .Q ( new_AGEMA_signal_9588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5113 ( .C ( clk ), .D ( new_AGEMA_signal_9601 ), .Q ( new_AGEMA_signal_9602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5121 ( .C ( clk ), .D ( n2516 ), .Q ( new_AGEMA_signal_9610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5129 ( .C ( clk ), .D ( new_AGEMA_signal_2466 ), .Q ( new_AGEMA_signal_9618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5137 ( .C ( clk ), .D ( new_AGEMA_signal_2467 ), .Q ( new_AGEMA_signal_9626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5145 ( .C ( clk ), .D ( n2808 ), .Q ( new_AGEMA_signal_9634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5153 ( .C ( clk ), .D ( new_AGEMA_signal_2496 ), .Q ( new_AGEMA_signal_9642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5161 ( .C ( clk ), .D ( new_AGEMA_signal_2497 ), .Q ( new_AGEMA_signal_9650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5193 ( .C ( clk ), .D ( new_AGEMA_signal_9681 ), .Q ( new_AGEMA_signal_9682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5209 ( .C ( clk ), .D ( new_AGEMA_signal_9697 ), .Q ( new_AGEMA_signal_9698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5225 ( .C ( clk ), .D ( new_AGEMA_signal_9713 ), .Q ( new_AGEMA_signal_9714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5259 ( .C ( clk ), .D ( new_AGEMA_signal_9747 ), .Q ( new_AGEMA_signal_9748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5275 ( .C ( clk ), .D ( new_AGEMA_signal_9763 ), .Q ( new_AGEMA_signal_9764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5291 ( .C ( clk ), .D ( new_AGEMA_signal_9779 ), .Q ( new_AGEMA_signal_9780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5301 ( .C ( clk ), .D ( n2527 ), .Q ( new_AGEMA_signal_9790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5311 ( .C ( clk ), .D ( new_AGEMA_signal_2574 ), .Q ( new_AGEMA_signal_9800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5321 ( .C ( clk ), .D ( new_AGEMA_signal_2575 ), .Q ( new_AGEMA_signal_9810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5407 ( .C ( clk ), .D ( new_AGEMA_signal_9895 ), .Q ( new_AGEMA_signal_9896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5423 ( .C ( clk ), .D ( new_AGEMA_signal_9911 ), .Q ( new_AGEMA_signal_9912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5439 ( .C ( clk ), .D ( new_AGEMA_signal_9927 ), .Q ( new_AGEMA_signal_9928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5487 ( .C ( clk ), .D ( new_AGEMA_signal_9975 ), .Q ( new_AGEMA_signal_9976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5505 ( .C ( clk ), .D ( new_AGEMA_signal_9993 ), .Q ( new_AGEMA_signal_9994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5523 ( .C ( clk ), .D ( new_AGEMA_signal_10011 ), .Q ( new_AGEMA_signal_10012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5637 ( .C ( clk ), .D ( new_AGEMA_signal_10125 ), .Q ( new_AGEMA_signal_10126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5657 ( .C ( clk ), .D ( new_AGEMA_signal_10145 ), .Q ( new_AGEMA_signal_10146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5677 ( .C ( clk ), .D ( new_AGEMA_signal_10165 ), .Q ( new_AGEMA_signal_10166 ) ) ;

    /* cells in depth 14 */
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2002 ( .a ({new_AGEMA_signal_7743, new_AGEMA_signal_7741, new_AGEMA_signal_7739}), .b ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, n1933}), .clk ( clk ), .r ({Fresh[2171], Fresh[2170], Fresh[2169]}), .c ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, n1935}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2054 ( .a ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, n1958}), .b ({new_AGEMA_signal_7767, new_AGEMA_signal_7759, new_AGEMA_signal_7751}), .clk ( clk ), .r ({Fresh[2174], Fresh[2173], Fresh[2172]}), .c ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, n1959}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2109 ( .a ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, n1982}), .b ({new_AGEMA_signal_7773, new_AGEMA_signal_7771, new_AGEMA_signal_7769}), .clk ( clk ), .r ({Fresh[2177], Fresh[2176], Fresh[2175]}), .c ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, n1983}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2149 ( .a ({new_AGEMA_signal_7785, new_AGEMA_signal_7781, new_AGEMA_signal_7777}), .b ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, n2011}), .clk ( clk ), .r ({Fresh[2180], Fresh[2179], Fresh[2178]}), .c ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, n2014}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2166 ( .a ({new_AGEMA_signal_7809, new_AGEMA_signal_7801, new_AGEMA_signal_7793}), .b ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, n2025}), .clk ( clk ), .r ({Fresh[2183], Fresh[2182], Fresh[2181]}), .c ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, n2029}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2180 ( .a ({new_AGEMA_signal_7815, new_AGEMA_signal_7813, new_AGEMA_signal_7811}), .b ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, n2036}), .clk ( clk ), .r ({Fresh[2186], Fresh[2185], Fresh[2184]}), .c ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, n2037}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2197 ( .a ({new_AGEMA_signal_7833, new_AGEMA_signal_7827, new_AGEMA_signal_7821}), .b ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, n2049}), .clk ( clk ), .r ({Fresh[2189], Fresh[2188], Fresh[2187]}), .c ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, n2052}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2219 ( .a ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, n2067}), .b ({new_AGEMA_signal_7845, new_AGEMA_signal_7841, new_AGEMA_signal_7837}), .clk ( clk ), .r ({Fresh[2192], Fresh[2191], Fresh[2190]}), .c ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, n2070}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2258 ( .a ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, n2097}), .b ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, n2096}), .clk ( clk ), .r ({Fresh[2195], Fresh[2194], Fresh[2193]}), .c ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, n2098}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2287 ( .a ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, n2124}), .b ({new_AGEMA_signal_7869, new_AGEMA_signal_7861, new_AGEMA_signal_7853}), .clk ( clk ), .r ({Fresh[2198], Fresh[2197], Fresh[2196]}), .c ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, n2125}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2311 ( .a ({new_AGEMA_signal_7881, new_AGEMA_signal_7877, new_AGEMA_signal_7873}), .b ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, n2142}), .clk ( clk ), .r ({Fresh[2201], Fresh[2200], Fresh[2199]}), .c ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, n2145}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2333 ( .a ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, n2168}), .b ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, n2167}), .clk ( clk ), .r ({Fresh[2204], Fresh[2203], Fresh[2202]}), .c ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, n2169}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2350 ( .a ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, n2184}), .b ({new_AGEMA_signal_7899, new_AGEMA_signal_7893, new_AGEMA_signal_7887}), .clk ( clk ), .r ({Fresh[2207], Fresh[2206], Fresh[2205]}), .c ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, n2185}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2365 ( .a ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, n2197}), .b ({new_AGEMA_signal_7917, new_AGEMA_signal_7911, new_AGEMA_signal_7905}), .clk ( clk ), .r ({Fresh[2210], Fresh[2209], Fresh[2208]}), .c ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, n2198}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2396 ( .a ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, n2232}), .b ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, n2231}), .clk ( clk ), .r ({Fresh[2213], Fresh[2212], Fresh[2211]}), .c ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, n2312}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2404 ( .a ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, n2239}), .b ({new_AGEMA_signal_7935, new_AGEMA_signal_7929, new_AGEMA_signal_7923}), .clk ( clk ), .r ({Fresh[2216], Fresh[2215], Fresh[2214]}), .c ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, n2258}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2415 ( .a ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, n2250}), .b ({new_AGEMA_signal_7953, new_AGEMA_signal_7947, new_AGEMA_signal_7941}), .clk ( clk ), .r ({Fresh[2219], Fresh[2218], Fresh[2217]}), .c ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, n2251}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2440 ( .a ({new_AGEMA_signal_7971, new_AGEMA_signal_7965, new_AGEMA_signal_7959}), .b ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, n2272}), .clk ( clk ), .r ({Fresh[2222], Fresh[2221], Fresh[2220]}), .c ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, n2274}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2469 ( .a ({new_AGEMA_signal_7983, new_AGEMA_signal_7979, new_AGEMA_signal_7975}), .b ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, n2296}), .clk ( clk ), .r ({Fresh[2225], Fresh[2224], Fresh[2223]}), .c ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, n2302}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2490 ( .a ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, n2324}), .b ({new_AGEMA_signal_8007, new_AGEMA_signal_7999, new_AGEMA_signal_7991}), .clk ( clk ), .r ({Fresh[2228], Fresh[2227], Fresh[2226]}), .c ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, n2339}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2503 ( .a ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, n2337}), .b ({new_AGEMA_signal_8019, new_AGEMA_signal_8015, new_AGEMA_signal_8011}), .clk ( clk ), .r ({Fresh[2231], Fresh[2230], Fresh[2229]}), .c ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, n2338}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2515 ( .a ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, n2350}), .b ({new_AGEMA_signal_8037, new_AGEMA_signal_8031, new_AGEMA_signal_8025}), .clk ( clk ), .r ({Fresh[2234], Fresh[2233], Fresh[2232]}), .c ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, n2351}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2529 ( .a ({new_AGEMA_signal_8061, new_AGEMA_signal_8053, new_AGEMA_signal_8045}), .b ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, n2362}), .clk ( clk ), .r ({Fresh[2237], Fresh[2236], Fresh[2235]}), .c ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, n2365}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2551 ( .a ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, n2389}), .b ({new_AGEMA_signal_8067, new_AGEMA_signal_8065, new_AGEMA_signal_8063}), .clk ( clk ), .r ({Fresh[2240], Fresh[2239], Fresh[2238]}), .c ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, n2399}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2560 ( .a ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, n2397}), .b ({new_AGEMA_signal_8085, new_AGEMA_signal_8079, new_AGEMA_signal_8073}), .clk ( clk ), .r ({Fresh[2243], Fresh[2242], Fresh[2241]}), .c ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, n2398}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2572 ( .a ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, n2411}), .b ({new_AGEMA_signal_8091, new_AGEMA_signal_8089, new_AGEMA_signal_8087}), .clk ( clk ), .r ({Fresh[2246], Fresh[2245], Fresh[2244]}), .c ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, n2423}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2581 ( .a ({new_AGEMA_signal_8097, new_AGEMA_signal_8095, new_AGEMA_signal_8093}), .b ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, n2420}), .clk ( clk ), .r ({Fresh[2249], Fresh[2248], Fresh[2247]}), .c ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, n2422}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2596 ( .a ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, n2440}), .b ({new_AGEMA_signal_8115, new_AGEMA_signal_8109, new_AGEMA_signal_8103}), .clk ( clk ), .r ({Fresh[2252], Fresh[2251], Fresh[2250]}), .c ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, n2441}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2623 ( .a ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, n2471}), .b ({new_AGEMA_signal_8133, new_AGEMA_signal_8127, new_AGEMA_signal_8121}), .clk ( clk ), .r ({Fresh[2255], Fresh[2254], Fresh[2253]}), .c ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, n2479}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2637 ( .a ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, n2485}), .b ({new_AGEMA_signal_8157, new_AGEMA_signal_8149, new_AGEMA_signal_8141}), .clk ( clk ), .r ({Fresh[2258], Fresh[2257], Fresh[2256]}), .c ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, n2512}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2652 ( .a ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, n2502}), .b ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, n2501}), .clk ( clk ), .r ({Fresh[2261], Fresh[2260], Fresh[2259]}), .c ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, n2510}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2686 ( .a ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, n2550}), .b ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, n2549}), .clk ( clk ), .r ({Fresh[2264], Fresh[2263], Fresh[2262]}), .c ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, n2552}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2702 ( .a ({new_AGEMA_signal_8181, new_AGEMA_signal_8173, new_AGEMA_signal_8165}), .b ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, n2569}), .clk ( clk ), .r ({Fresh[2267], Fresh[2266], Fresh[2265]}), .c ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, n2593}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2713 ( .a ({new_AGEMA_signal_8199, new_AGEMA_signal_8193, new_AGEMA_signal_8187}), .b ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, n2584}), .clk ( clk ), .r ({Fresh[2270], Fresh[2269], Fresh[2268]}), .c ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, n2589}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2730 ( .a ({new_AGEMA_signal_8217, new_AGEMA_signal_8211, new_AGEMA_signal_8205}), .b ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, n2606}), .clk ( clk ), .r ({Fresh[2273], Fresh[2272], Fresh[2271]}), .c ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, n2608}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2748 ( .a ({new_AGEMA_signal_8223, new_AGEMA_signal_8221, new_AGEMA_signal_8219}), .b ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, n2634}), .clk ( clk ), .r ({Fresh[2276], Fresh[2275], Fresh[2274]}), .c ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, n2636}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2762 ( .a ({new_AGEMA_signal_8235, new_AGEMA_signal_8231, new_AGEMA_signal_8227}), .b ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, n2657}), .clk ( clk ), .r ({Fresh[2279], Fresh[2278], Fresh[2277]}), .c ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, n2659}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2784 ( .a ({new_AGEMA_signal_8247, new_AGEMA_signal_8243, new_AGEMA_signal_8239}), .b ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, n2697}), .clk ( clk ), .r ({Fresh[2282], Fresh[2281], Fresh[2280]}), .c ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, n2702}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2811 ( .a ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, n2747}), .b ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, n2746}), .clk ( clk ), .r ({Fresh[2285], Fresh[2284], Fresh[2283]}), .c ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, n2806}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2839 ( .a ({new_AGEMA_signal_8259, new_AGEMA_signal_8255, new_AGEMA_signal_8251}), .b ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, n2799}), .clk ( clk ), .r ({Fresh[2288], Fresh[2287], Fresh[2286]}), .c ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, n2801}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2853 ( .a ({new_AGEMA_signal_8265, new_AGEMA_signal_8263, new_AGEMA_signal_8261}), .b ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, n2827}), .clk ( clk ), .r ({Fresh[2291], Fresh[2290], Fresh[2289]}), .c ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, n2829}) ) ;
    buf_clk new_AGEMA_reg_buffer_3782 ( .C ( clk ), .D ( new_AGEMA_signal_8270 ), .Q ( new_AGEMA_signal_8271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3788 ( .C ( clk ), .D ( new_AGEMA_signal_8276 ), .Q ( new_AGEMA_signal_8277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3794 ( .C ( clk ), .D ( new_AGEMA_signal_8282 ), .Q ( new_AGEMA_signal_8283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3796 ( .C ( clk ), .D ( new_AGEMA_signal_8284 ), .Q ( new_AGEMA_signal_8285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3798 ( .C ( clk ), .D ( new_AGEMA_signal_8286 ), .Q ( new_AGEMA_signal_8287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3800 ( .C ( clk ), .D ( new_AGEMA_signal_8288 ), .Q ( new_AGEMA_signal_8289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3804 ( .C ( clk ), .D ( new_AGEMA_signal_8292 ), .Q ( new_AGEMA_signal_8293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3808 ( .C ( clk ), .D ( new_AGEMA_signal_8296 ), .Q ( new_AGEMA_signal_8297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3812 ( .C ( clk ), .D ( new_AGEMA_signal_8300 ), .Q ( new_AGEMA_signal_8301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3820 ( .C ( clk ), .D ( new_AGEMA_signal_8308 ), .Q ( new_AGEMA_signal_8309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3828 ( .C ( clk ), .D ( new_AGEMA_signal_8316 ), .Q ( new_AGEMA_signal_8317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3836 ( .C ( clk ), .D ( new_AGEMA_signal_8324 ), .Q ( new_AGEMA_signal_8325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3844 ( .C ( clk ), .D ( new_AGEMA_signal_8332 ), .Q ( new_AGEMA_signal_8333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3852 ( .C ( clk ), .D ( new_AGEMA_signal_8340 ), .Q ( new_AGEMA_signal_8341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3860 ( .C ( clk ), .D ( new_AGEMA_signal_8348 ), .Q ( new_AGEMA_signal_8349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3868 ( .C ( clk ), .D ( new_AGEMA_signal_8356 ), .Q ( new_AGEMA_signal_8357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3876 ( .C ( clk ), .D ( new_AGEMA_signal_8364 ), .Q ( new_AGEMA_signal_8365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3884 ( .C ( clk ), .D ( new_AGEMA_signal_8372 ), .Q ( new_AGEMA_signal_8373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3892 ( .C ( clk ), .D ( new_AGEMA_signal_8380 ), .Q ( new_AGEMA_signal_8381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3900 ( .C ( clk ), .D ( new_AGEMA_signal_8388 ), .Q ( new_AGEMA_signal_8389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3908 ( .C ( clk ), .D ( new_AGEMA_signal_8396 ), .Q ( new_AGEMA_signal_8397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3914 ( .C ( clk ), .D ( new_AGEMA_signal_8402 ), .Q ( new_AGEMA_signal_8403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3920 ( .C ( clk ), .D ( new_AGEMA_signal_8408 ), .Q ( new_AGEMA_signal_8409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3926 ( .C ( clk ), .D ( new_AGEMA_signal_8414 ), .Q ( new_AGEMA_signal_8415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3936 ( .C ( clk ), .D ( new_AGEMA_signal_8424 ), .Q ( new_AGEMA_signal_8425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3946 ( .C ( clk ), .D ( new_AGEMA_signal_8434 ), .Q ( new_AGEMA_signal_8435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3956 ( .C ( clk ), .D ( new_AGEMA_signal_8444 ), .Q ( new_AGEMA_signal_8445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3964 ( .C ( clk ), .D ( new_AGEMA_signal_8452 ), .Q ( new_AGEMA_signal_8453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3972 ( .C ( clk ), .D ( new_AGEMA_signal_8460 ), .Q ( new_AGEMA_signal_8461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3980 ( .C ( clk ), .D ( new_AGEMA_signal_8468 ), .Q ( new_AGEMA_signal_8469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3988 ( .C ( clk ), .D ( new_AGEMA_signal_8476 ), .Q ( new_AGEMA_signal_8477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3996 ( .C ( clk ), .D ( new_AGEMA_signal_8484 ), .Q ( new_AGEMA_signal_8485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4004 ( .C ( clk ), .D ( new_AGEMA_signal_8492 ), .Q ( new_AGEMA_signal_8493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4012 ( .C ( clk ), .D ( new_AGEMA_signal_8500 ), .Q ( new_AGEMA_signal_8501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4020 ( .C ( clk ), .D ( new_AGEMA_signal_8508 ), .Q ( new_AGEMA_signal_8509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4028 ( .C ( clk ), .D ( new_AGEMA_signal_8516 ), .Q ( new_AGEMA_signal_8517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4030 ( .C ( clk ), .D ( new_AGEMA_signal_8518 ), .Q ( new_AGEMA_signal_8519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4032 ( .C ( clk ), .D ( new_AGEMA_signal_8520 ), .Q ( new_AGEMA_signal_8521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4034 ( .C ( clk ), .D ( new_AGEMA_signal_8522 ), .Q ( new_AGEMA_signal_8523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4038 ( .C ( clk ), .D ( new_AGEMA_signal_8526 ), .Q ( new_AGEMA_signal_8527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4042 ( .C ( clk ), .D ( new_AGEMA_signal_8530 ), .Q ( new_AGEMA_signal_8531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4046 ( .C ( clk ), .D ( new_AGEMA_signal_8534 ), .Q ( new_AGEMA_signal_8535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4052 ( .C ( clk ), .D ( new_AGEMA_signal_8540 ), .Q ( new_AGEMA_signal_8541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4058 ( .C ( clk ), .D ( new_AGEMA_signal_8546 ), .Q ( new_AGEMA_signal_8547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4064 ( .C ( clk ), .D ( new_AGEMA_signal_8552 ), .Q ( new_AGEMA_signal_8553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4068 ( .C ( clk ), .D ( new_AGEMA_signal_8556 ), .Q ( new_AGEMA_signal_8557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4072 ( .C ( clk ), .D ( new_AGEMA_signal_8560 ), .Q ( new_AGEMA_signal_8561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4076 ( .C ( clk ), .D ( new_AGEMA_signal_8564 ), .Q ( new_AGEMA_signal_8565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4086 ( .C ( clk ), .D ( new_AGEMA_signal_8574 ), .Q ( new_AGEMA_signal_8575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4096 ( .C ( clk ), .D ( new_AGEMA_signal_8584 ), .Q ( new_AGEMA_signal_8585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4106 ( .C ( clk ), .D ( new_AGEMA_signal_8594 ), .Q ( new_AGEMA_signal_8595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4114 ( .C ( clk ), .D ( new_AGEMA_signal_8602 ), .Q ( new_AGEMA_signal_8603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4122 ( .C ( clk ), .D ( new_AGEMA_signal_8610 ), .Q ( new_AGEMA_signal_8611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4130 ( .C ( clk ), .D ( new_AGEMA_signal_8618 ), .Q ( new_AGEMA_signal_8619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4134 ( .C ( clk ), .D ( new_AGEMA_signal_8622 ), .Q ( new_AGEMA_signal_8623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4138 ( .C ( clk ), .D ( new_AGEMA_signal_8626 ), .Q ( new_AGEMA_signal_8627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4142 ( .C ( clk ), .D ( new_AGEMA_signal_8630 ), .Q ( new_AGEMA_signal_8631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4144 ( .C ( clk ), .D ( new_AGEMA_signal_8632 ), .Q ( new_AGEMA_signal_8633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4146 ( .C ( clk ), .D ( new_AGEMA_signal_8634 ), .Q ( new_AGEMA_signal_8635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4148 ( .C ( clk ), .D ( new_AGEMA_signal_8636 ), .Q ( new_AGEMA_signal_8637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4156 ( .C ( clk ), .D ( new_AGEMA_signal_8644 ), .Q ( new_AGEMA_signal_8645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4164 ( .C ( clk ), .D ( new_AGEMA_signal_8652 ), .Q ( new_AGEMA_signal_8653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4172 ( .C ( clk ), .D ( new_AGEMA_signal_8660 ), .Q ( new_AGEMA_signal_8661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4180 ( .C ( clk ), .D ( new_AGEMA_signal_8668 ), .Q ( new_AGEMA_signal_8669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4188 ( .C ( clk ), .D ( new_AGEMA_signal_8676 ), .Q ( new_AGEMA_signal_8677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4196 ( .C ( clk ), .D ( new_AGEMA_signal_8684 ), .Q ( new_AGEMA_signal_8685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4202 ( .C ( clk ), .D ( new_AGEMA_signal_8690 ), .Q ( new_AGEMA_signal_8691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4208 ( .C ( clk ), .D ( new_AGEMA_signal_8696 ), .Q ( new_AGEMA_signal_8697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4214 ( .C ( clk ), .D ( new_AGEMA_signal_8702 ), .Q ( new_AGEMA_signal_8703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4218 ( .C ( clk ), .D ( new_AGEMA_signal_8706 ), .Q ( new_AGEMA_signal_8707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4222 ( .C ( clk ), .D ( new_AGEMA_signal_8710 ), .Q ( new_AGEMA_signal_8711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4226 ( .C ( clk ), .D ( new_AGEMA_signal_8714 ), .Q ( new_AGEMA_signal_8715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4234 ( .C ( clk ), .D ( new_AGEMA_signal_8722 ), .Q ( new_AGEMA_signal_8723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4242 ( .C ( clk ), .D ( new_AGEMA_signal_8730 ), .Q ( new_AGEMA_signal_8731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4250 ( .C ( clk ), .D ( new_AGEMA_signal_8738 ), .Q ( new_AGEMA_signal_8739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4252 ( .C ( clk ), .D ( new_AGEMA_signal_8740 ), .Q ( new_AGEMA_signal_8741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4254 ( .C ( clk ), .D ( new_AGEMA_signal_8742 ), .Q ( new_AGEMA_signal_8743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4256 ( .C ( clk ), .D ( new_AGEMA_signal_8744 ), .Q ( new_AGEMA_signal_8745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4260 ( .C ( clk ), .D ( new_AGEMA_signal_8748 ), .Q ( new_AGEMA_signal_8749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4266 ( .C ( clk ), .D ( new_AGEMA_signal_8754 ), .Q ( new_AGEMA_signal_8755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4272 ( .C ( clk ), .D ( new_AGEMA_signal_8760 ), .Q ( new_AGEMA_signal_8761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4278 ( .C ( clk ), .D ( new_AGEMA_signal_8766 ), .Q ( new_AGEMA_signal_8767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4284 ( .C ( clk ), .D ( new_AGEMA_signal_8772 ), .Q ( new_AGEMA_signal_8773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4290 ( .C ( clk ), .D ( new_AGEMA_signal_8778 ), .Q ( new_AGEMA_signal_8779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4296 ( .C ( clk ), .D ( new_AGEMA_signal_8784 ), .Q ( new_AGEMA_signal_8785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4302 ( .C ( clk ), .D ( new_AGEMA_signal_8790 ), .Q ( new_AGEMA_signal_8791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4308 ( .C ( clk ), .D ( new_AGEMA_signal_8796 ), .Q ( new_AGEMA_signal_8797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4312 ( .C ( clk ), .D ( new_AGEMA_signal_8800 ), .Q ( new_AGEMA_signal_8801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4316 ( .C ( clk ), .D ( new_AGEMA_signal_8804 ), .Q ( new_AGEMA_signal_8805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4320 ( .C ( clk ), .D ( new_AGEMA_signal_8808 ), .Q ( new_AGEMA_signal_8809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4328 ( .C ( clk ), .D ( new_AGEMA_signal_8816 ), .Q ( new_AGEMA_signal_8817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4336 ( .C ( clk ), .D ( new_AGEMA_signal_8824 ), .Q ( new_AGEMA_signal_8825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4344 ( .C ( clk ), .D ( new_AGEMA_signal_8832 ), .Q ( new_AGEMA_signal_8833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4350 ( .C ( clk ), .D ( new_AGEMA_signal_8838 ), .Q ( new_AGEMA_signal_8839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4356 ( .C ( clk ), .D ( new_AGEMA_signal_8844 ), .Q ( new_AGEMA_signal_8845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4362 ( .C ( clk ), .D ( new_AGEMA_signal_8850 ), .Q ( new_AGEMA_signal_8851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4366 ( .C ( clk ), .D ( new_AGEMA_signal_8854 ), .Q ( new_AGEMA_signal_8855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4370 ( .C ( clk ), .D ( new_AGEMA_signal_8858 ), .Q ( new_AGEMA_signal_8859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4374 ( .C ( clk ), .D ( new_AGEMA_signal_8862 ), .Q ( new_AGEMA_signal_8863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4382 ( .C ( clk ), .D ( new_AGEMA_signal_8870 ), .Q ( new_AGEMA_signal_8871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4390 ( .C ( clk ), .D ( new_AGEMA_signal_8878 ), .Q ( new_AGEMA_signal_8879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4398 ( .C ( clk ), .D ( new_AGEMA_signal_8886 ), .Q ( new_AGEMA_signal_8887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4406 ( .C ( clk ), .D ( new_AGEMA_signal_8894 ), .Q ( new_AGEMA_signal_8895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4414 ( .C ( clk ), .D ( new_AGEMA_signal_8902 ), .Q ( new_AGEMA_signal_8903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4422 ( .C ( clk ), .D ( new_AGEMA_signal_8910 ), .Q ( new_AGEMA_signal_8911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4432 ( .C ( clk ), .D ( new_AGEMA_signal_8920 ), .Q ( new_AGEMA_signal_8921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4442 ( .C ( clk ), .D ( new_AGEMA_signal_8930 ), .Q ( new_AGEMA_signal_8931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4452 ( .C ( clk ), .D ( new_AGEMA_signal_8940 ), .Q ( new_AGEMA_signal_8941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4460 ( .C ( clk ), .D ( new_AGEMA_signal_8948 ), .Q ( new_AGEMA_signal_8949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4468 ( .C ( clk ), .D ( new_AGEMA_signal_8956 ), .Q ( new_AGEMA_signal_8957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4476 ( .C ( clk ), .D ( new_AGEMA_signal_8964 ), .Q ( new_AGEMA_signal_8965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4482 ( .C ( clk ), .D ( new_AGEMA_signal_8970 ), .Q ( new_AGEMA_signal_8971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4488 ( .C ( clk ), .D ( new_AGEMA_signal_8976 ), .Q ( new_AGEMA_signal_8977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4494 ( .C ( clk ), .D ( new_AGEMA_signal_8982 ), .Q ( new_AGEMA_signal_8983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4498 ( .C ( clk ), .D ( new_AGEMA_signal_8986 ), .Q ( new_AGEMA_signal_8987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4502 ( .C ( clk ), .D ( new_AGEMA_signal_8990 ), .Q ( new_AGEMA_signal_8991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4506 ( .C ( clk ), .D ( new_AGEMA_signal_8994 ), .Q ( new_AGEMA_signal_8995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4512 ( .C ( clk ), .D ( new_AGEMA_signal_9000 ), .Q ( new_AGEMA_signal_9001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4518 ( .C ( clk ), .D ( new_AGEMA_signal_9006 ), .Q ( new_AGEMA_signal_9007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4524 ( .C ( clk ), .D ( new_AGEMA_signal_9012 ), .Q ( new_AGEMA_signal_9013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4532 ( .C ( clk ), .D ( new_AGEMA_signal_9020 ), .Q ( new_AGEMA_signal_9021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4540 ( .C ( clk ), .D ( new_AGEMA_signal_9028 ), .Q ( new_AGEMA_signal_9029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4548 ( .C ( clk ), .D ( new_AGEMA_signal_9036 ), .Q ( new_AGEMA_signal_9037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4554 ( .C ( clk ), .D ( new_AGEMA_signal_9042 ), .Q ( new_AGEMA_signal_9043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4560 ( .C ( clk ), .D ( new_AGEMA_signal_9048 ), .Q ( new_AGEMA_signal_9049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4566 ( .C ( clk ), .D ( new_AGEMA_signal_9054 ), .Q ( new_AGEMA_signal_9055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4580 ( .C ( clk ), .D ( new_AGEMA_signal_9068 ), .Q ( new_AGEMA_signal_9069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4588 ( .C ( clk ), .D ( new_AGEMA_signal_9076 ), .Q ( new_AGEMA_signal_9077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4596 ( .C ( clk ), .D ( new_AGEMA_signal_9084 ), .Q ( new_AGEMA_signal_9085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4600 ( .C ( clk ), .D ( new_AGEMA_signal_9088 ), .Q ( new_AGEMA_signal_9089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4604 ( .C ( clk ), .D ( new_AGEMA_signal_9092 ), .Q ( new_AGEMA_signal_9093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4608 ( .C ( clk ), .D ( new_AGEMA_signal_9096 ), .Q ( new_AGEMA_signal_9097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4614 ( .C ( clk ), .D ( new_AGEMA_signal_9102 ), .Q ( new_AGEMA_signal_9103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4620 ( .C ( clk ), .D ( new_AGEMA_signal_9108 ), .Q ( new_AGEMA_signal_9109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4626 ( .C ( clk ), .D ( new_AGEMA_signal_9114 ), .Q ( new_AGEMA_signal_9115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4632 ( .C ( clk ), .D ( new_AGEMA_signal_9120 ), .Q ( new_AGEMA_signal_9121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4638 ( .C ( clk ), .D ( new_AGEMA_signal_9126 ), .Q ( new_AGEMA_signal_9127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4644 ( .C ( clk ), .D ( new_AGEMA_signal_9132 ), .Q ( new_AGEMA_signal_9133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4648 ( .C ( clk ), .D ( new_AGEMA_signal_9136 ), .Q ( new_AGEMA_signal_9137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4652 ( .C ( clk ), .D ( new_AGEMA_signal_9140 ), .Q ( new_AGEMA_signal_9141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4656 ( .C ( clk ), .D ( new_AGEMA_signal_9144 ), .Q ( new_AGEMA_signal_9145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4660 ( .C ( clk ), .D ( new_AGEMA_signal_9148 ), .Q ( new_AGEMA_signal_9149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4666 ( .C ( clk ), .D ( new_AGEMA_signal_9154 ), .Q ( new_AGEMA_signal_9155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4672 ( .C ( clk ), .D ( new_AGEMA_signal_9160 ), .Q ( new_AGEMA_signal_9161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4690 ( .C ( clk ), .D ( new_AGEMA_signal_9178 ), .Q ( new_AGEMA_signal_9179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4696 ( .C ( clk ), .D ( new_AGEMA_signal_9184 ), .Q ( new_AGEMA_signal_9185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4702 ( .C ( clk ), .D ( new_AGEMA_signal_9190 ), .Q ( new_AGEMA_signal_9191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4712 ( .C ( clk ), .D ( new_AGEMA_signal_9200 ), .Q ( new_AGEMA_signal_9201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4722 ( .C ( clk ), .D ( new_AGEMA_signal_9210 ), .Q ( new_AGEMA_signal_9211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4732 ( .C ( clk ), .D ( new_AGEMA_signal_9220 ), .Q ( new_AGEMA_signal_9221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4738 ( .C ( clk ), .D ( new_AGEMA_signal_9226 ), .Q ( new_AGEMA_signal_9227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4744 ( .C ( clk ), .D ( new_AGEMA_signal_9232 ), .Q ( new_AGEMA_signal_9233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4750 ( .C ( clk ), .D ( new_AGEMA_signal_9238 ), .Q ( new_AGEMA_signal_9239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4756 ( .C ( clk ), .D ( new_AGEMA_signal_9244 ), .Q ( new_AGEMA_signal_9245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4762 ( .C ( clk ), .D ( new_AGEMA_signal_9250 ), .Q ( new_AGEMA_signal_9251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4768 ( .C ( clk ), .D ( new_AGEMA_signal_9256 ), .Q ( new_AGEMA_signal_9257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4800 ( .C ( clk ), .D ( new_AGEMA_signal_9288 ), .Q ( new_AGEMA_signal_9289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4808 ( .C ( clk ), .D ( new_AGEMA_signal_9296 ), .Q ( new_AGEMA_signal_9297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4816 ( .C ( clk ), .D ( new_AGEMA_signal_9304 ), .Q ( new_AGEMA_signal_9305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4822 ( .C ( clk ), .D ( new_AGEMA_signal_9310 ), .Q ( new_AGEMA_signal_9311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4828 ( .C ( clk ), .D ( new_AGEMA_signal_9316 ), .Q ( new_AGEMA_signal_9317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4834 ( .C ( clk ), .D ( new_AGEMA_signal_9322 ), .Q ( new_AGEMA_signal_9323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4842 ( .C ( clk ), .D ( new_AGEMA_signal_9330 ), .Q ( new_AGEMA_signal_9331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4850 ( .C ( clk ), .D ( new_AGEMA_signal_9338 ), .Q ( new_AGEMA_signal_9339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4858 ( .C ( clk ), .D ( new_AGEMA_signal_9346 ), .Q ( new_AGEMA_signal_9347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4866 ( .C ( clk ), .D ( new_AGEMA_signal_9354 ), .Q ( new_AGEMA_signal_9355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4874 ( .C ( clk ), .D ( new_AGEMA_signal_9362 ), .Q ( new_AGEMA_signal_9363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4882 ( .C ( clk ), .D ( new_AGEMA_signal_9370 ), .Q ( new_AGEMA_signal_9371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4920 ( .C ( clk ), .D ( new_AGEMA_signal_9408 ), .Q ( new_AGEMA_signal_9409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4928 ( .C ( clk ), .D ( new_AGEMA_signal_9416 ), .Q ( new_AGEMA_signal_9417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4936 ( .C ( clk ), .D ( new_AGEMA_signal_9424 ), .Q ( new_AGEMA_signal_9425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4954 ( .C ( clk ), .D ( new_AGEMA_signal_9442 ), .Q ( new_AGEMA_signal_9443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4962 ( .C ( clk ), .D ( new_AGEMA_signal_9450 ), .Q ( new_AGEMA_signal_9451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4970 ( .C ( clk ), .D ( new_AGEMA_signal_9458 ), .Q ( new_AGEMA_signal_9459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4982 ( .C ( clk ), .D ( new_AGEMA_signal_9470 ), .Q ( new_AGEMA_signal_9471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4994 ( .C ( clk ), .D ( new_AGEMA_signal_9482 ), .Q ( new_AGEMA_signal_9483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5006 ( .C ( clk ), .D ( new_AGEMA_signal_9494 ), .Q ( new_AGEMA_signal_9495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5020 ( .C ( clk ), .D ( new_AGEMA_signal_9508 ), .Q ( new_AGEMA_signal_9509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5034 ( .C ( clk ), .D ( new_AGEMA_signal_9522 ), .Q ( new_AGEMA_signal_9523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5048 ( .C ( clk ), .D ( new_AGEMA_signal_9536 ), .Q ( new_AGEMA_signal_9537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5056 ( .C ( clk ), .D ( new_AGEMA_signal_9544 ), .Q ( new_AGEMA_signal_9545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5064 ( .C ( clk ), .D ( new_AGEMA_signal_9552 ), .Q ( new_AGEMA_signal_9553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5072 ( .C ( clk ), .D ( new_AGEMA_signal_9560 ), .Q ( new_AGEMA_signal_9561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5086 ( .C ( clk ), .D ( new_AGEMA_signal_9574 ), .Q ( new_AGEMA_signal_9575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5100 ( .C ( clk ), .D ( new_AGEMA_signal_9588 ), .Q ( new_AGEMA_signal_9589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5114 ( .C ( clk ), .D ( new_AGEMA_signal_9602 ), .Q ( new_AGEMA_signal_9603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5122 ( .C ( clk ), .D ( new_AGEMA_signal_9610 ), .Q ( new_AGEMA_signal_9611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5130 ( .C ( clk ), .D ( new_AGEMA_signal_9618 ), .Q ( new_AGEMA_signal_9619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5138 ( .C ( clk ), .D ( new_AGEMA_signal_9626 ), .Q ( new_AGEMA_signal_9627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5146 ( .C ( clk ), .D ( new_AGEMA_signal_9634 ), .Q ( new_AGEMA_signal_9635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5154 ( .C ( clk ), .D ( new_AGEMA_signal_9642 ), .Q ( new_AGEMA_signal_9643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5162 ( .C ( clk ), .D ( new_AGEMA_signal_9650 ), .Q ( new_AGEMA_signal_9651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5194 ( .C ( clk ), .D ( new_AGEMA_signal_9682 ), .Q ( new_AGEMA_signal_9683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5210 ( .C ( clk ), .D ( new_AGEMA_signal_9698 ), .Q ( new_AGEMA_signal_9699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5226 ( .C ( clk ), .D ( new_AGEMA_signal_9714 ), .Q ( new_AGEMA_signal_9715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5260 ( .C ( clk ), .D ( new_AGEMA_signal_9748 ), .Q ( new_AGEMA_signal_9749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5276 ( .C ( clk ), .D ( new_AGEMA_signal_9764 ), .Q ( new_AGEMA_signal_9765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5292 ( .C ( clk ), .D ( new_AGEMA_signal_9780 ), .Q ( new_AGEMA_signal_9781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5302 ( .C ( clk ), .D ( new_AGEMA_signal_9790 ), .Q ( new_AGEMA_signal_9791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5312 ( .C ( clk ), .D ( new_AGEMA_signal_9800 ), .Q ( new_AGEMA_signal_9801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5322 ( .C ( clk ), .D ( new_AGEMA_signal_9810 ), .Q ( new_AGEMA_signal_9811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5408 ( .C ( clk ), .D ( new_AGEMA_signal_9896 ), .Q ( new_AGEMA_signal_9897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5424 ( .C ( clk ), .D ( new_AGEMA_signal_9912 ), .Q ( new_AGEMA_signal_9913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5440 ( .C ( clk ), .D ( new_AGEMA_signal_9928 ), .Q ( new_AGEMA_signal_9929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5488 ( .C ( clk ), .D ( new_AGEMA_signal_9976 ), .Q ( new_AGEMA_signal_9977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5506 ( .C ( clk ), .D ( new_AGEMA_signal_9994 ), .Q ( new_AGEMA_signal_9995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5524 ( .C ( clk ), .D ( new_AGEMA_signal_10012 ), .Q ( new_AGEMA_signal_10013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5638 ( .C ( clk ), .D ( new_AGEMA_signal_10126 ), .Q ( new_AGEMA_signal_10127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5658 ( .C ( clk ), .D ( new_AGEMA_signal_10146 ), .Q ( new_AGEMA_signal_10147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5678 ( .C ( clk ), .D ( new_AGEMA_signal_10166 ), .Q ( new_AGEMA_signal_10167 ) ) ;

    /* cells in depth 15 */
    buf_clk new_AGEMA_reg_buffer_4261 ( .C ( clk ), .D ( new_AGEMA_signal_8749 ), .Q ( new_AGEMA_signal_8750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4267 ( .C ( clk ), .D ( new_AGEMA_signal_8755 ), .Q ( new_AGEMA_signal_8756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4273 ( .C ( clk ), .D ( new_AGEMA_signal_8761 ), .Q ( new_AGEMA_signal_8762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4279 ( .C ( clk ), .D ( new_AGEMA_signal_8767 ), .Q ( new_AGEMA_signal_8768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4285 ( .C ( clk ), .D ( new_AGEMA_signal_8773 ), .Q ( new_AGEMA_signal_8774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4291 ( .C ( clk ), .D ( new_AGEMA_signal_8779 ), .Q ( new_AGEMA_signal_8780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4297 ( .C ( clk ), .D ( new_AGEMA_signal_8785 ), .Q ( new_AGEMA_signal_8786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4303 ( .C ( clk ), .D ( new_AGEMA_signal_8791 ), .Q ( new_AGEMA_signal_8792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4309 ( .C ( clk ), .D ( new_AGEMA_signal_8797 ), .Q ( new_AGEMA_signal_8798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4313 ( .C ( clk ), .D ( new_AGEMA_signal_8801 ), .Q ( new_AGEMA_signal_8802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4317 ( .C ( clk ), .D ( new_AGEMA_signal_8805 ), .Q ( new_AGEMA_signal_8806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4321 ( .C ( clk ), .D ( new_AGEMA_signal_8809 ), .Q ( new_AGEMA_signal_8810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4329 ( .C ( clk ), .D ( new_AGEMA_signal_8817 ), .Q ( new_AGEMA_signal_8818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4337 ( .C ( clk ), .D ( new_AGEMA_signal_8825 ), .Q ( new_AGEMA_signal_8826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4345 ( .C ( clk ), .D ( new_AGEMA_signal_8833 ), .Q ( new_AGEMA_signal_8834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4351 ( .C ( clk ), .D ( new_AGEMA_signal_8839 ), .Q ( new_AGEMA_signal_8840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4357 ( .C ( clk ), .D ( new_AGEMA_signal_8845 ), .Q ( new_AGEMA_signal_8846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4363 ( .C ( clk ), .D ( new_AGEMA_signal_8851 ), .Q ( new_AGEMA_signal_8852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4367 ( .C ( clk ), .D ( new_AGEMA_signal_8855 ), .Q ( new_AGEMA_signal_8856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4371 ( .C ( clk ), .D ( new_AGEMA_signal_8859 ), .Q ( new_AGEMA_signal_8860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4375 ( .C ( clk ), .D ( new_AGEMA_signal_8863 ), .Q ( new_AGEMA_signal_8864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4383 ( .C ( clk ), .D ( new_AGEMA_signal_8871 ), .Q ( new_AGEMA_signal_8872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4391 ( .C ( clk ), .D ( new_AGEMA_signal_8879 ), .Q ( new_AGEMA_signal_8880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4399 ( .C ( clk ), .D ( new_AGEMA_signal_8887 ), .Q ( new_AGEMA_signal_8888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4407 ( .C ( clk ), .D ( new_AGEMA_signal_8895 ), .Q ( new_AGEMA_signal_8896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4415 ( .C ( clk ), .D ( new_AGEMA_signal_8903 ), .Q ( new_AGEMA_signal_8904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4423 ( .C ( clk ), .D ( new_AGEMA_signal_8911 ), .Q ( new_AGEMA_signal_8912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4433 ( .C ( clk ), .D ( new_AGEMA_signal_8921 ), .Q ( new_AGEMA_signal_8922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4443 ( .C ( clk ), .D ( new_AGEMA_signal_8931 ), .Q ( new_AGEMA_signal_8932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4453 ( .C ( clk ), .D ( new_AGEMA_signal_8941 ), .Q ( new_AGEMA_signal_8942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4461 ( .C ( clk ), .D ( new_AGEMA_signal_8949 ), .Q ( new_AGEMA_signal_8950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4469 ( .C ( clk ), .D ( new_AGEMA_signal_8957 ), .Q ( new_AGEMA_signal_8958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4477 ( .C ( clk ), .D ( new_AGEMA_signal_8965 ), .Q ( new_AGEMA_signal_8966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4483 ( .C ( clk ), .D ( new_AGEMA_signal_8971 ), .Q ( new_AGEMA_signal_8972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4489 ( .C ( clk ), .D ( new_AGEMA_signal_8977 ), .Q ( new_AGEMA_signal_8978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4495 ( .C ( clk ), .D ( new_AGEMA_signal_8983 ), .Q ( new_AGEMA_signal_8984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4499 ( .C ( clk ), .D ( new_AGEMA_signal_8987 ), .Q ( new_AGEMA_signal_8988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4503 ( .C ( clk ), .D ( new_AGEMA_signal_8991 ), .Q ( new_AGEMA_signal_8992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4507 ( .C ( clk ), .D ( new_AGEMA_signal_8995 ), .Q ( new_AGEMA_signal_8996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4513 ( .C ( clk ), .D ( new_AGEMA_signal_9001 ), .Q ( new_AGEMA_signal_9002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4519 ( .C ( clk ), .D ( new_AGEMA_signal_9007 ), .Q ( new_AGEMA_signal_9008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4525 ( .C ( clk ), .D ( new_AGEMA_signal_9013 ), .Q ( new_AGEMA_signal_9014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4533 ( .C ( clk ), .D ( new_AGEMA_signal_9021 ), .Q ( new_AGEMA_signal_9022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4541 ( .C ( clk ), .D ( new_AGEMA_signal_9029 ), .Q ( new_AGEMA_signal_9030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4549 ( .C ( clk ), .D ( new_AGEMA_signal_9037 ), .Q ( new_AGEMA_signal_9038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4555 ( .C ( clk ), .D ( new_AGEMA_signal_9043 ), .Q ( new_AGEMA_signal_9044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4561 ( .C ( clk ), .D ( new_AGEMA_signal_9049 ), .Q ( new_AGEMA_signal_9050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4567 ( .C ( clk ), .D ( new_AGEMA_signal_9055 ), .Q ( new_AGEMA_signal_9056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4569 ( .C ( clk ), .D ( n2512 ), .Q ( new_AGEMA_signal_9058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4571 ( .C ( clk ), .D ( new_AGEMA_signal_2568 ), .Q ( new_AGEMA_signal_9060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4573 ( .C ( clk ), .D ( new_AGEMA_signal_2569 ), .Q ( new_AGEMA_signal_9062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4581 ( .C ( clk ), .D ( new_AGEMA_signal_9069 ), .Q ( new_AGEMA_signal_9070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4589 ( .C ( clk ), .D ( new_AGEMA_signal_9077 ), .Q ( new_AGEMA_signal_9078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4597 ( .C ( clk ), .D ( new_AGEMA_signal_9085 ), .Q ( new_AGEMA_signal_9086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4601 ( .C ( clk ), .D ( new_AGEMA_signal_9089 ), .Q ( new_AGEMA_signal_9090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4605 ( .C ( clk ), .D ( new_AGEMA_signal_9093 ), .Q ( new_AGEMA_signal_9094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4609 ( .C ( clk ), .D ( new_AGEMA_signal_9097 ), .Q ( new_AGEMA_signal_9098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4615 ( .C ( clk ), .D ( new_AGEMA_signal_9103 ), .Q ( new_AGEMA_signal_9104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4621 ( .C ( clk ), .D ( new_AGEMA_signal_9109 ), .Q ( new_AGEMA_signal_9110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4627 ( .C ( clk ), .D ( new_AGEMA_signal_9115 ), .Q ( new_AGEMA_signal_9116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4633 ( .C ( clk ), .D ( new_AGEMA_signal_9121 ), .Q ( new_AGEMA_signal_9122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4639 ( .C ( clk ), .D ( new_AGEMA_signal_9127 ), .Q ( new_AGEMA_signal_9128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4645 ( .C ( clk ), .D ( new_AGEMA_signal_9133 ), .Q ( new_AGEMA_signal_9134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4649 ( .C ( clk ), .D ( new_AGEMA_signal_9137 ), .Q ( new_AGEMA_signal_9138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4653 ( .C ( clk ), .D ( new_AGEMA_signal_9141 ), .Q ( new_AGEMA_signal_9142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4657 ( .C ( clk ), .D ( new_AGEMA_signal_9145 ), .Q ( new_AGEMA_signal_9146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4661 ( .C ( clk ), .D ( new_AGEMA_signal_9149 ), .Q ( new_AGEMA_signal_9150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4667 ( .C ( clk ), .D ( new_AGEMA_signal_9155 ), .Q ( new_AGEMA_signal_9156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4673 ( .C ( clk ), .D ( new_AGEMA_signal_9161 ), .Q ( new_AGEMA_signal_9162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4677 ( .C ( clk ), .D ( n2037 ), .Q ( new_AGEMA_signal_9166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4681 ( .C ( clk ), .D ( new_AGEMA_signal_2520 ), .Q ( new_AGEMA_signal_9170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4685 ( .C ( clk ), .D ( new_AGEMA_signal_2521 ), .Q ( new_AGEMA_signal_9174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4691 ( .C ( clk ), .D ( new_AGEMA_signal_9179 ), .Q ( new_AGEMA_signal_9180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4697 ( .C ( clk ), .D ( new_AGEMA_signal_9185 ), .Q ( new_AGEMA_signal_9186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4703 ( .C ( clk ), .D ( new_AGEMA_signal_9191 ), .Q ( new_AGEMA_signal_9192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4713 ( .C ( clk ), .D ( new_AGEMA_signal_9201 ), .Q ( new_AGEMA_signal_9202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4723 ( .C ( clk ), .D ( new_AGEMA_signal_9211 ), .Q ( new_AGEMA_signal_9212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4733 ( .C ( clk ), .D ( new_AGEMA_signal_9221 ), .Q ( new_AGEMA_signal_9222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4739 ( .C ( clk ), .D ( new_AGEMA_signal_9227 ), .Q ( new_AGEMA_signal_9228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4745 ( .C ( clk ), .D ( new_AGEMA_signal_9233 ), .Q ( new_AGEMA_signal_9234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4751 ( .C ( clk ), .D ( new_AGEMA_signal_9239 ), .Q ( new_AGEMA_signal_9240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4757 ( .C ( clk ), .D ( new_AGEMA_signal_9245 ), .Q ( new_AGEMA_signal_9246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4763 ( .C ( clk ), .D ( new_AGEMA_signal_9251 ), .Q ( new_AGEMA_signal_9252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4769 ( .C ( clk ), .D ( new_AGEMA_signal_9257 ), .Q ( new_AGEMA_signal_9258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4773 ( .C ( clk ), .D ( n2198 ), .Q ( new_AGEMA_signal_9262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4777 ( .C ( clk ), .D ( new_AGEMA_signal_2538 ), .Q ( new_AGEMA_signal_9266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4781 ( .C ( clk ), .D ( new_AGEMA_signal_2539 ), .Q ( new_AGEMA_signal_9270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4785 ( .C ( clk ), .D ( n2258 ), .Q ( new_AGEMA_signal_9274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4789 ( .C ( clk ), .D ( new_AGEMA_signal_2620 ), .Q ( new_AGEMA_signal_9278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4793 ( .C ( clk ), .D ( new_AGEMA_signal_2621 ), .Q ( new_AGEMA_signal_9282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4801 ( .C ( clk ), .D ( new_AGEMA_signal_9289 ), .Q ( new_AGEMA_signal_9290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4809 ( .C ( clk ), .D ( new_AGEMA_signal_9297 ), .Q ( new_AGEMA_signal_9298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4817 ( .C ( clk ), .D ( new_AGEMA_signal_9305 ), .Q ( new_AGEMA_signal_9306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4823 ( .C ( clk ), .D ( new_AGEMA_signal_9311 ), .Q ( new_AGEMA_signal_9312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4829 ( .C ( clk ), .D ( new_AGEMA_signal_9317 ), .Q ( new_AGEMA_signal_9318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4835 ( .C ( clk ), .D ( new_AGEMA_signal_9323 ), .Q ( new_AGEMA_signal_9324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4843 ( .C ( clk ), .D ( new_AGEMA_signal_9331 ), .Q ( new_AGEMA_signal_9332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4851 ( .C ( clk ), .D ( new_AGEMA_signal_9339 ), .Q ( new_AGEMA_signal_9340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4859 ( .C ( clk ), .D ( new_AGEMA_signal_9347 ), .Q ( new_AGEMA_signal_9348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4867 ( .C ( clk ), .D ( new_AGEMA_signal_9355 ), .Q ( new_AGEMA_signal_9356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4875 ( .C ( clk ), .D ( new_AGEMA_signal_9363 ), .Q ( new_AGEMA_signal_9364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4883 ( .C ( clk ), .D ( new_AGEMA_signal_9371 ), .Q ( new_AGEMA_signal_9372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4893 ( .C ( clk ), .D ( n2593 ), .Q ( new_AGEMA_signal_9382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4897 ( .C ( clk ), .D ( new_AGEMA_signal_2578 ), .Q ( new_AGEMA_signal_9386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4901 ( .C ( clk ), .D ( new_AGEMA_signal_2579 ), .Q ( new_AGEMA_signal_9390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4905 ( .C ( clk ), .D ( n2636 ), .Q ( new_AGEMA_signal_9394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4909 ( .C ( clk ), .D ( new_AGEMA_signal_2584 ), .Q ( new_AGEMA_signal_9398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4913 ( .C ( clk ), .D ( new_AGEMA_signal_2585 ), .Q ( new_AGEMA_signal_9402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4921 ( .C ( clk ), .D ( new_AGEMA_signal_9409 ), .Q ( new_AGEMA_signal_9410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4929 ( .C ( clk ), .D ( new_AGEMA_signal_9417 ), .Q ( new_AGEMA_signal_9418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4937 ( .C ( clk ), .D ( new_AGEMA_signal_9425 ), .Q ( new_AGEMA_signal_9426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4941 ( .C ( clk ), .D ( n2806 ), .Q ( new_AGEMA_signal_9430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4945 ( .C ( clk ), .D ( new_AGEMA_signal_2590 ), .Q ( new_AGEMA_signal_9434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4949 ( .C ( clk ), .D ( new_AGEMA_signal_2591 ), .Q ( new_AGEMA_signal_9438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4955 ( .C ( clk ), .D ( new_AGEMA_signal_9443 ), .Q ( new_AGEMA_signal_9444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4963 ( .C ( clk ), .D ( new_AGEMA_signal_9451 ), .Q ( new_AGEMA_signal_9452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4971 ( .C ( clk ), .D ( new_AGEMA_signal_9459 ), .Q ( new_AGEMA_signal_9460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4983 ( .C ( clk ), .D ( new_AGEMA_signal_9471 ), .Q ( new_AGEMA_signal_9472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4995 ( .C ( clk ), .D ( new_AGEMA_signal_9483 ), .Q ( new_AGEMA_signal_9484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5007 ( .C ( clk ), .D ( new_AGEMA_signal_9495 ), .Q ( new_AGEMA_signal_9496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5021 ( .C ( clk ), .D ( new_AGEMA_signal_9509 ), .Q ( new_AGEMA_signal_9510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5035 ( .C ( clk ), .D ( new_AGEMA_signal_9523 ), .Q ( new_AGEMA_signal_9524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5049 ( .C ( clk ), .D ( new_AGEMA_signal_9537 ), .Q ( new_AGEMA_signal_9538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5057 ( .C ( clk ), .D ( new_AGEMA_signal_9545 ), .Q ( new_AGEMA_signal_9546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5065 ( .C ( clk ), .D ( new_AGEMA_signal_9553 ), .Q ( new_AGEMA_signal_9554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5073 ( .C ( clk ), .D ( new_AGEMA_signal_9561 ), .Q ( new_AGEMA_signal_9562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5087 ( .C ( clk ), .D ( new_AGEMA_signal_9575 ), .Q ( new_AGEMA_signal_9576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5101 ( .C ( clk ), .D ( new_AGEMA_signal_9589 ), .Q ( new_AGEMA_signal_9590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5115 ( .C ( clk ), .D ( new_AGEMA_signal_9603 ), .Q ( new_AGEMA_signal_9604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5123 ( .C ( clk ), .D ( new_AGEMA_signal_9611 ), .Q ( new_AGEMA_signal_9612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5131 ( .C ( clk ), .D ( new_AGEMA_signal_9619 ), .Q ( new_AGEMA_signal_9620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5139 ( .C ( clk ), .D ( new_AGEMA_signal_9627 ), .Q ( new_AGEMA_signal_9628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5147 ( .C ( clk ), .D ( new_AGEMA_signal_9635 ), .Q ( new_AGEMA_signal_9636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5155 ( .C ( clk ), .D ( new_AGEMA_signal_9643 ), .Q ( new_AGEMA_signal_9644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5163 ( .C ( clk ), .D ( new_AGEMA_signal_9651 ), .Q ( new_AGEMA_signal_9652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5195 ( .C ( clk ), .D ( new_AGEMA_signal_9683 ), .Q ( new_AGEMA_signal_9684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5211 ( .C ( clk ), .D ( new_AGEMA_signal_9699 ), .Q ( new_AGEMA_signal_9700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5227 ( .C ( clk ), .D ( new_AGEMA_signal_9715 ), .Q ( new_AGEMA_signal_9716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5261 ( .C ( clk ), .D ( new_AGEMA_signal_9749 ), .Q ( new_AGEMA_signal_9750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5277 ( .C ( clk ), .D ( new_AGEMA_signal_9765 ), .Q ( new_AGEMA_signal_9766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5293 ( .C ( clk ), .D ( new_AGEMA_signal_9781 ), .Q ( new_AGEMA_signal_9782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5303 ( .C ( clk ), .D ( new_AGEMA_signal_9791 ), .Q ( new_AGEMA_signal_9792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5313 ( .C ( clk ), .D ( new_AGEMA_signal_9801 ), .Q ( new_AGEMA_signal_9802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5323 ( .C ( clk ), .D ( new_AGEMA_signal_9811 ), .Q ( new_AGEMA_signal_9812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5343 ( .C ( clk ), .D ( n2829 ), .Q ( new_AGEMA_signal_9832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5351 ( .C ( clk ), .D ( new_AGEMA_signal_2594 ), .Q ( new_AGEMA_signal_9840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5359 ( .C ( clk ), .D ( new_AGEMA_signal_2595 ), .Q ( new_AGEMA_signal_9848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5409 ( .C ( clk ), .D ( new_AGEMA_signal_9897 ), .Q ( new_AGEMA_signal_9898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5425 ( .C ( clk ), .D ( new_AGEMA_signal_9913 ), .Q ( new_AGEMA_signal_9914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5441 ( .C ( clk ), .D ( new_AGEMA_signal_9929 ), .Q ( new_AGEMA_signal_9930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5451 ( .C ( clk ), .D ( n2312 ), .Q ( new_AGEMA_signal_9940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5461 ( .C ( clk ), .D ( new_AGEMA_signal_2542 ), .Q ( new_AGEMA_signal_9950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5471 ( .C ( clk ), .D ( new_AGEMA_signal_2543 ), .Q ( new_AGEMA_signal_9960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5489 ( .C ( clk ), .D ( new_AGEMA_signal_9977 ), .Q ( new_AGEMA_signal_9978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5507 ( .C ( clk ), .D ( new_AGEMA_signal_9995 ), .Q ( new_AGEMA_signal_9996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5525 ( .C ( clk ), .D ( new_AGEMA_signal_10013 ), .Q ( new_AGEMA_signal_10014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5639 ( .C ( clk ), .D ( new_AGEMA_signal_10127 ), .Q ( new_AGEMA_signal_10128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5659 ( .C ( clk ), .D ( new_AGEMA_signal_10147 ), .Q ( new_AGEMA_signal_10148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5679 ( .C ( clk ), .D ( new_AGEMA_signal_10167 ), .Q ( new_AGEMA_signal_10168 ) ) ;

    /* cells in depth 16 */
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2003 ( .a ({new_AGEMA_signal_8283, new_AGEMA_signal_8277, new_AGEMA_signal_8271}), .b ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, n1935}), .clk ( clk ), .r ({Fresh[2294], Fresh[2293], Fresh[2292]}), .c ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, n1941}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2059 ( .a ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, n1959}), .b ({new_AGEMA_signal_8289, new_AGEMA_signal_8287, new_AGEMA_signal_8285}), .clk ( clk ), .r ({Fresh[2297], Fresh[2296], Fresh[2295]}), .c ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, n1960}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2110 ( .a ({new_AGEMA_signal_8301, new_AGEMA_signal_8297, new_AGEMA_signal_8293}), .b ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, n1983}), .clk ( clk ), .r ({Fresh[2300], Fresh[2299], Fresh[2298]}), .c ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, n1988}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2153 ( .a ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, n2014}), .b ({new_AGEMA_signal_8325, new_AGEMA_signal_8317, new_AGEMA_signal_8309}), .clk ( clk ), .r ({Fresh[2303], Fresh[2302], Fresh[2301]}), .c ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, n2015}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2169 ( .a ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, n2029}), .b ({new_AGEMA_signal_8349, new_AGEMA_signal_8341, new_AGEMA_signal_8333}), .clk ( clk ), .r ({Fresh[2306], Fresh[2305], Fresh[2304]}), .c ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, n2030}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2200 ( .a ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, n2052}), .b ({new_AGEMA_signal_8373, new_AGEMA_signal_8365, new_AGEMA_signal_8357}), .clk ( clk ), .r ({Fresh[2309], Fresh[2308], Fresh[2307]}), .c ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, n2053}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2222 ( .a ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, n2070}), .b ({new_AGEMA_signal_8397, new_AGEMA_signal_8389, new_AGEMA_signal_8381}), .clk ( clk ), .r ({Fresh[2312], Fresh[2311], Fresh[2310]}), .c ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, n2071}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2259 ( .a ({new_AGEMA_signal_8415, new_AGEMA_signal_8409, new_AGEMA_signal_8403}), .b ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, n2098}), .clk ( clk ), .r ({Fresh[2315], Fresh[2314], Fresh[2313]}), .c ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, n2103}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2288 ( .a ({new_AGEMA_signal_8445, new_AGEMA_signal_8435, new_AGEMA_signal_8425}), .b ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, n2125}), .clk ( clk ), .r ({Fresh[2318], Fresh[2317], Fresh[2316]}), .c ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, n2126}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2314 ( .a ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, n2145}), .b ({new_AGEMA_signal_8469, new_AGEMA_signal_8461, new_AGEMA_signal_8453}), .clk ( clk ), .r ({Fresh[2321], Fresh[2320], Fresh[2319]}), .c ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, n2146}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2334 ( .a ({new_AGEMA_signal_8493, new_AGEMA_signal_8485, new_AGEMA_signal_8477}), .b ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, n2169}), .clk ( clk ), .r ({Fresh[2324], Fresh[2323], Fresh[2322]}), .c ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, n2173}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2351 ( .a ({new_AGEMA_signal_8517, new_AGEMA_signal_8509, new_AGEMA_signal_8501}), .b ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, n2185}), .clk ( clk ), .r ({Fresh[2327], Fresh[2326], Fresh[2325]}), .c ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, n2187}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2416 ( .a ({new_AGEMA_signal_8523, new_AGEMA_signal_8521, new_AGEMA_signal_8519}), .b ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, n2251}), .clk ( clk ), .r ({Fresh[2330], Fresh[2329], Fresh[2328]}), .c ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, n2256}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2441 ( .a ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, n2274}), .b ({new_AGEMA_signal_8535, new_AGEMA_signal_8531, new_AGEMA_signal_8527}), .clk ( clk ), .r ({Fresh[2333], Fresh[2332], Fresh[2331]}), .c ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, n2275}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2474 ( .a ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, n2302}), .b ({new_AGEMA_signal_8553, new_AGEMA_signal_8547, new_AGEMA_signal_8541}), .clk ( clk ), .r ({Fresh[2336], Fresh[2335], Fresh[2334]}), .c ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, n2303}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2504 ( .a ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, n2339}), .b ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, n2338}), .clk ( clk ), .r ({Fresh[2339], Fresh[2338], Fresh[2337]}), .c ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, n2382}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2516 ( .a ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, n2351}), .b ({new_AGEMA_signal_8565, new_AGEMA_signal_8561, new_AGEMA_signal_8557}), .clk ( clk ), .r ({Fresh[2342], Fresh[2341], Fresh[2340]}), .c ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, n2380}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2531 ( .a ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, n2365}), .b ({new_AGEMA_signal_8595, new_AGEMA_signal_8585, new_AGEMA_signal_8575}), .clk ( clk ), .r ({Fresh[2345], Fresh[2344], Fresh[2343]}), .c ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, n2366}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2561 ( .a ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, n2399}), .b ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, n2398}), .clk ( clk ), .r ({Fresh[2348], Fresh[2347], Fresh[2346]}), .c ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, n2425}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2582 ( .a ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, n2423}), .b ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, n2422}), .clk ( clk ), .r ({Fresh[2351], Fresh[2350], Fresh[2349]}), .c ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, n2424}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2597 ( .a ({new_AGEMA_signal_8619, new_AGEMA_signal_8611, new_AGEMA_signal_8603}), .b ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, n2441}), .clk ( clk ), .r ({Fresh[2354], Fresh[2353], Fresh[2352]}), .c ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, n2451}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2631 ( .a ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, n2479}), .b ({new_AGEMA_signal_8631, new_AGEMA_signal_8627, new_AGEMA_signal_8623}), .clk ( clk ), .r ({Fresh[2357], Fresh[2356], Fresh[2355]}), .c ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, n2514}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2658 ( .a ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, n2510}), .b ({new_AGEMA_signal_8637, new_AGEMA_signal_8635, new_AGEMA_signal_8633}), .clk ( clk ), .r ({Fresh[2360], Fresh[2359], Fresh[2358]}), .c ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, n2511}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2688 ( .a ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, n2552}), .b ({new_AGEMA_signal_8661, new_AGEMA_signal_8653, new_AGEMA_signal_8645}), .clk ( clk ), .r ({Fresh[2363], Fresh[2362], Fresh[2361]}), .c ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, n2671}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2716 ( .a ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, n2589}), .b ({new_AGEMA_signal_8685, new_AGEMA_signal_8677, new_AGEMA_signal_8669}), .clk ( clk ), .r ({Fresh[2366], Fresh[2365], Fresh[2364]}), .c ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, n2590}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2731 ( .a ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, n2608}), .b ({new_AGEMA_signal_8703, new_AGEMA_signal_8697, new_AGEMA_signal_8691}), .clk ( clk ), .r ({Fresh[2369], Fresh[2368], Fresh[2367]}), .c ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, n2623}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2763 ( .a ({new_AGEMA_signal_8715, new_AGEMA_signal_8711, new_AGEMA_signal_8707}), .b ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, n2659}), .clk ( clk ), .r ({Fresh[2372], Fresh[2371], Fresh[2370]}), .c ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, n2667}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2786 ( .a ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, n2702}), .b ({new_AGEMA_signal_8739, new_AGEMA_signal_8731, new_AGEMA_signal_8723}), .clk ( clk ), .r ({Fresh[2375], Fresh[2374], Fresh[2373]}), .c ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, n2703}) ) ;
    mux2_HPC2 #(.security_order(2), .pipeline(1)) U2840 ( .s ({new_AGEMA_signal_8535, new_AGEMA_signal_8531, new_AGEMA_signal_8527}), .b ({new_AGEMA_signal_8745, new_AGEMA_signal_8743, new_AGEMA_signal_8741}), .a ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, n2801}), .clk ( clk ), .r ({Fresh[2378], Fresh[2377], Fresh[2376]}), .c ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, n2803}) ) ;
    buf_clk new_AGEMA_reg_buffer_4262 ( .C ( clk ), .D ( new_AGEMA_signal_8750 ), .Q ( new_AGEMA_signal_8751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4268 ( .C ( clk ), .D ( new_AGEMA_signal_8756 ), .Q ( new_AGEMA_signal_8757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4274 ( .C ( clk ), .D ( new_AGEMA_signal_8762 ), .Q ( new_AGEMA_signal_8763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4280 ( .C ( clk ), .D ( new_AGEMA_signal_8768 ), .Q ( new_AGEMA_signal_8769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4286 ( .C ( clk ), .D ( new_AGEMA_signal_8774 ), .Q ( new_AGEMA_signal_8775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4292 ( .C ( clk ), .D ( new_AGEMA_signal_8780 ), .Q ( new_AGEMA_signal_8781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4298 ( .C ( clk ), .D ( new_AGEMA_signal_8786 ), .Q ( new_AGEMA_signal_8787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4304 ( .C ( clk ), .D ( new_AGEMA_signal_8792 ), .Q ( new_AGEMA_signal_8793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4310 ( .C ( clk ), .D ( new_AGEMA_signal_8798 ), .Q ( new_AGEMA_signal_8799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4314 ( .C ( clk ), .D ( new_AGEMA_signal_8802 ), .Q ( new_AGEMA_signal_8803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4318 ( .C ( clk ), .D ( new_AGEMA_signal_8806 ), .Q ( new_AGEMA_signal_8807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4322 ( .C ( clk ), .D ( new_AGEMA_signal_8810 ), .Q ( new_AGEMA_signal_8811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4330 ( .C ( clk ), .D ( new_AGEMA_signal_8818 ), .Q ( new_AGEMA_signal_8819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4338 ( .C ( clk ), .D ( new_AGEMA_signal_8826 ), .Q ( new_AGEMA_signal_8827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4346 ( .C ( clk ), .D ( new_AGEMA_signal_8834 ), .Q ( new_AGEMA_signal_8835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4352 ( .C ( clk ), .D ( new_AGEMA_signal_8840 ), .Q ( new_AGEMA_signal_8841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4358 ( .C ( clk ), .D ( new_AGEMA_signal_8846 ), .Q ( new_AGEMA_signal_8847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4364 ( .C ( clk ), .D ( new_AGEMA_signal_8852 ), .Q ( new_AGEMA_signal_8853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4368 ( .C ( clk ), .D ( new_AGEMA_signal_8856 ), .Q ( new_AGEMA_signal_8857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4372 ( .C ( clk ), .D ( new_AGEMA_signal_8860 ), .Q ( new_AGEMA_signal_8861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4376 ( .C ( clk ), .D ( new_AGEMA_signal_8864 ), .Q ( new_AGEMA_signal_8865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4384 ( .C ( clk ), .D ( new_AGEMA_signal_8872 ), .Q ( new_AGEMA_signal_8873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4392 ( .C ( clk ), .D ( new_AGEMA_signal_8880 ), .Q ( new_AGEMA_signal_8881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4400 ( .C ( clk ), .D ( new_AGEMA_signal_8888 ), .Q ( new_AGEMA_signal_8889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4408 ( .C ( clk ), .D ( new_AGEMA_signal_8896 ), .Q ( new_AGEMA_signal_8897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4416 ( .C ( clk ), .D ( new_AGEMA_signal_8904 ), .Q ( new_AGEMA_signal_8905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4424 ( .C ( clk ), .D ( new_AGEMA_signal_8912 ), .Q ( new_AGEMA_signal_8913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4434 ( .C ( clk ), .D ( new_AGEMA_signal_8922 ), .Q ( new_AGEMA_signal_8923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4444 ( .C ( clk ), .D ( new_AGEMA_signal_8932 ), .Q ( new_AGEMA_signal_8933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4454 ( .C ( clk ), .D ( new_AGEMA_signal_8942 ), .Q ( new_AGEMA_signal_8943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4462 ( .C ( clk ), .D ( new_AGEMA_signal_8950 ), .Q ( new_AGEMA_signal_8951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4470 ( .C ( clk ), .D ( new_AGEMA_signal_8958 ), .Q ( new_AGEMA_signal_8959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4478 ( .C ( clk ), .D ( new_AGEMA_signal_8966 ), .Q ( new_AGEMA_signal_8967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4484 ( .C ( clk ), .D ( new_AGEMA_signal_8972 ), .Q ( new_AGEMA_signal_8973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4490 ( .C ( clk ), .D ( new_AGEMA_signal_8978 ), .Q ( new_AGEMA_signal_8979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4496 ( .C ( clk ), .D ( new_AGEMA_signal_8984 ), .Q ( new_AGEMA_signal_8985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4500 ( .C ( clk ), .D ( new_AGEMA_signal_8988 ), .Q ( new_AGEMA_signal_8989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4504 ( .C ( clk ), .D ( new_AGEMA_signal_8992 ), .Q ( new_AGEMA_signal_8993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4508 ( .C ( clk ), .D ( new_AGEMA_signal_8996 ), .Q ( new_AGEMA_signal_8997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4514 ( .C ( clk ), .D ( new_AGEMA_signal_9002 ), .Q ( new_AGEMA_signal_9003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4520 ( .C ( clk ), .D ( new_AGEMA_signal_9008 ), .Q ( new_AGEMA_signal_9009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4526 ( .C ( clk ), .D ( new_AGEMA_signal_9014 ), .Q ( new_AGEMA_signal_9015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4534 ( .C ( clk ), .D ( new_AGEMA_signal_9022 ), .Q ( new_AGEMA_signal_9023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4542 ( .C ( clk ), .D ( new_AGEMA_signal_9030 ), .Q ( new_AGEMA_signal_9031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4550 ( .C ( clk ), .D ( new_AGEMA_signal_9038 ), .Q ( new_AGEMA_signal_9039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4556 ( .C ( clk ), .D ( new_AGEMA_signal_9044 ), .Q ( new_AGEMA_signal_9045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4562 ( .C ( clk ), .D ( new_AGEMA_signal_9050 ), .Q ( new_AGEMA_signal_9051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4568 ( .C ( clk ), .D ( new_AGEMA_signal_9056 ), .Q ( new_AGEMA_signal_9057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4570 ( .C ( clk ), .D ( new_AGEMA_signal_9058 ), .Q ( new_AGEMA_signal_9059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4572 ( .C ( clk ), .D ( new_AGEMA_signal_9060 ), .Q ( new_AGEMA_signal_9061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4574 ( .C ( clk ), .D ( new_AGEMA_signal_9062 ), .Q ( new_AGEMA_signal_9063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4582 ( .C ( clk ), .D ( new_AGEMA_signal_9070 ), .Q ( new_AGEMA_signal_9071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4590 ( .C ( clk ), .D ( new_AGEMA_signal_9078 ), .Q ( new_AGEMA_signal_9079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4598 ( .C ( clk ), .D ( new_AGEMA_signal_9086 ), .Q ( new_AGEMA_signal_9087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4602 ( .C ( clk ), .D ( new_AGEMA_signal_9090 ), .Q ( new_AGEMA_signal_9091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4606 ( .C ( clk ), .D ( new_AGEMA_signal_9094 ), .Q ( new_AGEMA_signal_9095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4610 ( .C ( clk ), .D ( new_AGEMA_signal_9098 ), .Q ( new_AGEMA_signal_9099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4616 ( .C ( clk ), .D ( new_AGEMA_signal_9104 ), .Q ( new_AGEMA_signal_9105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4622 ( .C ( clk ), .D ( new_AGEMA_signal_9110 ), .Q ( new_AGEMA_signal_9111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4628 ( .C ( clk ), .D ( new_AGEMA_signal_9116 ), .Q ( new_AGEMA_signal_9117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4634 ( .C ( clk ), .D ( new_AGEMA_signal_9122 ), .Q ( new_AGEMA_signal_9123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4640 ( .C ( clk ), .D ( new_AGEMA_signal_9128 ), .Q ( new_AGEMA_signal_9129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4646 ( .C ( clk ), .D ( new_AGEMA_signal_9134 ), .Q ( new_AGEMA_signal_9135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4650 ( .C ( clk ), .D ( new_AGEMA_signal_9138 ), .Q ( new_AGEMA_signal_9139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4654 ( .C ( clk ), .D ( new_AGEMA_signal_9142 ), .Q ( new_AGEMA_signal_9143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4658 ( .C ( clk ), .D ( new_AGEMA_signal_9146 ), .Q ( new_AGEMA_signal_9147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4662 ( .C ( clk ), .D ( new_AGEMA_signal_9150 ), .Q ( new_AGEMA_signal_9151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4668 ( .C ( clk ), .D ( new_AGEMA_signal_9156 ), .Q ( new_AGEMA_signal_9157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4674 ( .C ( clk ), .D ( new_AGEMA_signal_9162 ), .Q ( new_AGEMA_signal_9163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4678 ( .C ( clk ), .D ( new_AGEMA_signal_9166 ), .Q ( new_AGEMA_signal_9167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4682 ( .C ( clk ), .D ( new_AGEMA_signal_9170 ), .Q ( new_AGEMA_signal_9171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4686 ( .C ( clk ), .D ( new_AGEMA_signal_9174 ), .Q ( new_AGEMA_signal_9175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4692 ( .C ( clk ), .D ( new_AGEMA_signal_9180 ), .Q ( new_AGEMA_signal_9181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4698 ( .C ( clk ), .D ( new_AGEMA_signal_9186 ), .Q ( new_AGEMA_signal_9187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4704 ( .C ( clk ), .D ( new_AGEMA_signal_9192 ), .Q ( new_AGEMA_signal_9193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4714 ( .C ( clk ), .D ( new_AGEMA_signal_9202 ), .Q ( new_AGEMA_signal_9203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4724 ( .C ( clk ), .D ( new_AGEMA_signal_9212 ), .Q ( new_AGEMA_signal_9213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4734 ( .C ( clk ), .D ( new_AGEMA_signal_9222 ), .Q ( new_AGEMA_signal_9223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4740 ( .C ( clk ), .D ( new_AGEMA_signal_9228 ), .Q ( new_AGEMA_signal_9229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4746 ( .C ( clk ), .D ( new_AGEMA_signal_9234 ), .Q ( new_AGEMA_signal_9235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4752 ( .C ( clk ), .D ( new_AGEMA_signal_9240 ), .Q ( new_AGEMA_signal_9241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4758 ( .C ( clk ), .D ( new_AGEMA_signal_9246 ), .Q ( new_AGEMA_signal_9247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4764 ( .C ( clk ), .D ( new_AGEMA_signal_9252 ), .Q ( new_AGEMA_signal_9253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4770 ( .C ( clk ), .D ( new_AGEMA_signal_9258 ), .Q ( new_AGEMA_signal_9259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4774 ( .C ( clk ), .D ( new_AGEMA_signal_9262 ), .Q ( new_AGEMA_signal_9263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4778 ( .C ( clk ), .D ( new_AGEMA_signal_9266 ), .Q ( new_AGEMA_signal_9267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4782 ( .C ( clk ), .D ( new_AGEMA_signal_9270 ), .Q ( new_AGEMA_signal_9271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4786 ( .C ( clk ), .D ( new_AGEMA_signal_9274 ), .Q ( new_AGEMA_signal_9275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4790 ( .C ( clk ), .D ( new_AGEMA_signal_9278 ), .Q ( new_AGEMA_signal_9279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4794 ( .C ( clk ), .D ( new_AGEMA_signal_9282 ), .Q ( new_AGEMA_signal_9283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4802 ( .C ( clk ), .D ( new_AGEMA_signal_9290 ), .Q ( new_AGEMA_signal_9291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4810 ( .C ( clk ), .D ( new_AGEMA_signal_9298 ), .Q ( new_AGEMA_signal_9299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4818 ( .C ( clk ), .D ( new_AGEMA_signal_9306 ), .Q ( new_AGEMA_signal_9307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4824 ( .C ( clk ), .D ( new_AGEMA_signal_9312 ), .Q ( new_AGEMA_signal_9313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4830 ( .C ( clk ), .D ( new_AGEMA_signal_9318 ), .Q ( new_AGEMA_signal_9319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4836 ( .C ( clk ), .D ( new_AGEMA_signal_9324 ), .Q ( new_AGEMA_signal_9325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4844 ( .C ( clk ), .D ( new_AGEMA_signal_9332 ), .Q ( new_AGEMA_signal_9333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4852 ( .C ( clk ), .D ( new_AGEMA_signal_9340 ), .Q ( new_AGEMA_signal_9341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4860 ( .C ( clk ), .D ( new_AGEMA_signal_9348 ), .Q ( new_AGEMA_signal_9349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4868 ( .C ( clk ), .D ( new_AGEMA_signal_9356 ), .Q ( new_AGEMA_signal_9357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4876 ( .C ( clk ), .D ( new_AGEMA_signal_9364 ), .Q ( new_AGEMA_signal_9365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4884 ( .C ( clk ), .D ( new_AGEMA_signal_9372 ), .Q ( new_AGEMA_signal_9373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4894 ( .C ( clk ), .D ( new_AGEMA_signal_9382 ), .Q ( new_AGEMA_signal_9383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4898 ( .C ( clk ), .D ( new_AGEMA_signal_9386 ), .Q ( new_AGEMA_signal_9387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4902 ( .C ( clk ), .D ( new_AGEMA_signal_9390 ), .Q ( new_AGEMA_signal_9391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4906 ( .C ( clk ), .D ( new_AGEMA_signal_9394 ), .Q ( new_AGEMA_signal_9395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4910 ( .C ( clk ), .D ( new_AGEMA_signal_9398 ), .Q ( new_AGEMA_signal_9399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4914 ( .C ( clk ), .D ( new_AGEMA_signal_9402 ), .Q ( new_AGEMA_signal_9403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4922 ( .C ( clk ), .D ( new_AGEMA_signal_9410 ), .Q ( new_AGEMA_signal_9411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4930 ( .C ( clk ), .D ( new_AGEMA_signal_9418 ), .Q ( new_AGEMA_signal_9419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4938 ( .C ( clk ), .D ( new_AGEMA_signal_9426 ), .Q ( new_AGEMA_signal_9427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4942 ( .C ( clk ), .D ( new_AGEMA_signal_9430 ), .Q ( new_AGEMA_signal_9431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4946 ( .C ( clk ), .D ( new_AGEMA_signal_9434 ), .Q ( new_AGEMA_signal_9435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4950 ( .C ( clk ), .D ( new_AGEMA_signal_9438 ), .Q ( new_AGEMA_signal_9439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4956 ( .C ( clk ), .D ( new_AGEMA_signal_9444 ), .Q ( new_AGEMA_signal_9445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4964 ( .C ( clk ), .D ( new_AGEMA_signal_9452 ), .Q ( new_AGEMA_signal_9453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4972 ( .C ( clk ), .D ( new_AGEMA_signal_9460 ), .Q ( new_AGEMA_signal_9461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4984 ( .C ( clk ), .D ( new_AGEMA_signal_9472 ), .Q ( new_AGEMA_signal_9473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4996 ( .C ( clk ), .D ( new_AGEMA_signal_9484 ), .Q ( new_AGEMA_signal_9485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5008 ( .C ( clk ), .D ( new_AGEMA_signal_9496 ), .Q ( new_AGEMA_signal_9497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5022 ( .C ( clk ), .D ( new_AGEMA_signal_9510 ), .Q ( new_AGEMA_signal_9511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5036 ( .C ( clk ), .D ( new_AGEMA_signal_9524 ), .Q ( new_AGEMA_signal_9525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5050 ( .C ( clk ), .D ( new_AGEMA_signal_9538 ), .Q ( new_AGEMA_signal_9539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5058 ( .C ( clk ), .D ( new_AGEMA_signal_9546 ), .Q ( new_AGEMA_signal_9547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5066 ( .C ( clk ), .D ( new_AGEMA_signal_9554 ), .Q ( new_AGEMA_signal_9555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5074 ( .C ( clk ), .D ( new_AGEMA_signal_9562 ), .Q ( new_AGEMA_signal_9563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5088 ( .C ( clk ), .D ( new_AGEMA_signal_9576 ), .Q ( new_AGEMA_signal_9577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5102 ( .C ( clk ), .D ( new_AGEMA_signal_9590 ), .Q ( new_AGEMA_signal_9591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5116 ( .C ( clk ), .D ( new_AGEMA_signal_9604 ), .Q ( new_AGEMA_signal_9605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5124 ( .C ( clk ), .D ( new_AGEMA_signal_9612 ), .Q ( new_AGEMA_signal_9613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5132 ( .C ( clk ), .D ( new_AGEMA_signal_9620 ), .Q ( new_AGEMA_signal_9621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5140 ( .C ( clk ), .D ( new_AGEMA_signal_9628 ), .Q ( new_AGEMA_signal_9629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5148 ( .C ( clk ), .D ( new_AGEMA_signal_9636 ), .Q ( new_AGEMA_signal_9637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5156 ( .C ( clk ), .D ( new_AGEMA_signal_9644 ), .Q ( new_AGEMA_signal_9645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5164 ( .C ( clk ), .D ( new_AGEMA_signal_9652 ), .Q ( new_AGEMA_signal_9653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5196 ( .C ( clk ), .D ( new_AGEMA_signal_9684 ), .Q ( new_AGEMA_signal_9685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5212 ( .C ( clk ), .D ( new_AGEMA_signal_9700 ), .Q ( new_AGEMA_signal_9701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5228 ( .C ( clk ), .D ( new_AGEMA_signal_9716 ), .Q ( new_AGEMA_signal_9717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5262 ( .C ( clk ), .D ( new_AGEMA_signal_9750 ), .Q ( new_AGEMA_signal_9751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5278 ( .C ( clk ), .D ( new_AGEMA_signal_9766 ), .Q ( new_AGEMA_signal_9767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5294 ( .C ( clk ), .D ( new_AGEMA_signal_9782 ), .Q ( new_AGEMA_signal_9783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5304 ( .C ( clk ), .D ( new_AGEMA_signal_9792 ), .Q ( new_AGEMA_signal_9793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5314 ( .C ( clk ), .D ( new_AGEMA_signal_9802 ), .Q ( new_AGEMA_signal_9803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5324 ( .C ( clk ), .D ( new_AGEMA_signal_9812 ), .Q ( new_AGEMA_signal_9813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5344 ( .C ( clk ), .D ( new_AGEMA_signal_9832 ), .Q ( new_AGEMA_signal_9833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5352 ( .C ( clk ), .D ( new_AGEMA_signal_9840 ), .Q ( new_AGEMA_signal_9841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5360 ( .C ( clk ), .D ( new_AGEMA_signal_9848 ), .Q ( new_AGEMA_signal_9849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5410 ( .C ( clk ), .D ( new_AGEMA_signal_9898 ), .Q ( new_AGEMA_signal_9899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5426 ( .C ( clk ), .D ( new_AGEMA_signal_9914 ), .Q ( new_AGEMA_signal_9915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5442 ( .C ( clk ), .D ( new_AGEMA_signal_9930 ), .Q ( new_AGEMA_signal_9931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5452 ( .C ( clk ), .D ( new_AGEMA_signal_9940 ), .Q ( new_AGEMA_signal_9941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5462 ( .C ( clk ), .D ( new_AGEMA_signal_9950 ), .Q ( new_AGEMA_signal_9951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5472 ( .C ( clk ), .D ( new_AGEMA_signal_9960 ), .Q ( new_AGEMA_signal_9961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5490 ( .C ( clk ), .D ( new_AGEMA_signal_9978 ), .Q ( new_AGEMA_signal_9979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5508 ( .C ( clk ), .D ( new_AGEMA_signal_9996 ), .Q ( new_AGEMA_signal_9997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5526 ( .C ( clk ), .D ( new_AGEMA_signal_10014 ), .Q ( new_AGEMA_signal_10015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5640 ( .C ( clk ), .D ( new_AGEMA_signal_10128 ), .Q ( new_AGEMA_signal_10129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5660 ( .C ( clk ), .D ( new_AGEMA_signal_10148 ), .Q ( new_AGEMA_signal_10149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5680 ( .C ( clk ), .D ( new_AGEMA_signal_10168 ), .Q ( new_AGEMA_signal_10169 ) ) ;

    /* cells in depth 17 */
    buf_clk new_AGEMA_reg_buffer_4663 ( .C ( clk ), .D ( new_AGEMA_signal_9151 ), .Q ( new_AGEMA_signal_9152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4669 ( .C ( clk ), .D ( new_AGEMA_signal_9157 ), .Q ( new_AGEMA_signal_9158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4675 ( .C ( clk ), .D ( new_AGEMA_signal_9163 ), .Q ( new_AGEMA_signal_9164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4679 ( .C ( clk ), .D ( new_AGEMA_signal_9167 ), .Q ( new_AGEMA_signal_9168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4683 ( .C ( clk ), .D ( new_AGEMA_signal_9171 ), .Q ( new_AGEMA_signal_9172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4687 ( .C ( clk ), .D ( new_AGEMA_signal_9175 ), .Q ( new_AGEMA_signal_9176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4693 ( .C ( clk ), .D ( new_AGEMA_signal_9181 ), .Q ( new_AGEMA_signal_9182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4699 ( .C ( clk ), .D ( new_AGEMA_signal_9187 ), .Q ( new_AGEMA_signal_9188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4705 ( .C ( clk ), .D ( new_AGEMA_signal_9193 ), .Q ( new_AGEMA_signal_9194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4715 ( .C ( clk ), .D ( new_AGEMA_signal_9203 ), .Q ( new_AGEMA_signal_9204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4725 ( .C ( clk ), .D ( new_AGEMA_signal_9213 ), .Q ( new_AGEMA_signal_9214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4735 ( .C ( clk ), .D ( new_AGEMA_signal_9223 ), .Q ( new_AGEMA_signal_9224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4741 ( .C ( clk ), .D ( new_AGEMA_signal_9229 ), .Q ( new_AGEMA_signal_9230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4747 ( .C ( clk ), .D ( new_AGEMA_signal_9235 ), .Q ( new_AGEMA_signal_9236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4753 ( .C ( clk ), .D ( new_AGEMA_signal_9241 ), .Q ( new_AGEMA_signal_9242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4759 ( .C ( clk ), .D ( new_AGEMA_signal_9247 ), .Q ( new_AGEMA_signal_9248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4765 ( .C ( clk ), .D ( new_AGEMA_signal_9253 ), .Q ( new_AGEMA_signal_9254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4771 ( .C ( clk ), .D ( new_AGEMA_signal_9259 ), .Q ( new_AGEMA_signal_9260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4775 ( .C ( clk ), .D ( new_AGEMA_signal_9263 ), .Q ( new_AGEMA_signal_9264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4779 ( .C ( clk ), .D ( new_AGEMA_signal_9267 ), .Q ( new_AGEMA_signal_9268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4783 ( .C ( clk ), .D ( new_AGEMA_signal_9271 ), .Q ( new_AGEMA_signal_9272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4787 ( .C ( clk ), .D ( new_AGEMA_signal_9275 ), .Q ( new_AGEMA_signal_9276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4791 ( .C ( clk ), .D ( new_AGEMA_signal_9279 ), .Q ( new_AGEMA_signal_9280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4795 ( .C ( clk ), .D ( new_AGEMA_signal_9283 ), .Q ( new_AGEMA_signal_9284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4803 ( .C ( clk ), .D ( new_AGEMA_signal_9291 ), .Q ( new_AGEMA_signal_9292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4811 ( .C ( clk ), .D ( new_AGEMA_signal_9299 ), .Q ( new_AGEMA_signal_9300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4819 ( .C ( clk ), .D ( new_AGEMA_signal_9307 ), .Q ( new_AGEMA_signal_9308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4825 ( .C ( clk ), .D ( new_AGEMA_signal_9313 ), .Q ( new_AGEMA_signal_9314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4831 ( .C ( clk ), .D ( new_AGEMA_signal_9319 ), .Q ( new_AGEMA_signal_9320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4837 ( .C ( clk ), .D ( new_AGEMA_signal_9325 ), .Q ( new_AGEMA_signal_9326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4845 ( .C ( clk ), .D ( new_AGEMA_signal_9333 ), .Q ( new_AGEMA_signal_9334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4853 ( .C ( clk ), .D ( new_AGEMA_signal_9341 ), .Q ( new_AGEMA_signal_9342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4861 ( .C ( clk ), .D ( new_AGEMA_signal_9349 ), .Q ( new_AGEMA_signal_9350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4869 ( .C ( clk ), .D ( new_AGEMA_signal_9357 ), .Q ( new_AGEMA_signal_9358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4877 ( .C ( clk ), .D ( new_AGEMA_signal_9365 ), .Q ( new_AGEMA_signal_9366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4885 ( .C ( clk ), .D ( new_AGEMA_signal_9373 ), .Q ( new_AGEMA_signal_9374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4887 ( .C ( clk ), .D ( n2514 ), .Q ( new_AGEMA_signal_9376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4889 ( .C ( clk ), .D ( new_AGEMA_signal_2566 ), .Q ( new_AGEMA_signal_9378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4891 ( .C ( clk ), .D ( new_AGEMA_signal_2567 ), .Q ( new_AGEMA_signal_9380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4895 ( .C ( clk ), .D ( new_AGEMA_signal_9383 ), .Q ( new_AGEMA_signal_9384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4899 ( .C ( clk ), .D ( new_AGEMA_signal_9387 ), .Q ( new_AGEMA_signal_9388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4903 ( .C ( clk ), .D ( new_AGEMA_signal_9391 ), .Q ( new_AGEMA_signal_9392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4907 ( .C ( clk ), .D ( new_AGEMA_signal_9395 ), .Q ( new_AGEMA_signal_9396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4911 ( .C ( clk ), .D ( new_AGEMA_signal_9399 ), .Q ( new_AGEMA_signal_9400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4915 ( .C ( clk ), .D ( new_AGEMA_signal_9403 ), .Q ( new_AGEMA_signal_9404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4923 ( .C ( clk ), .D ( new_AGEMA_signal_9411 ), .Q ( new_AGEMA_signal_9412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4931 ( .C ( clk ), .D ( new_AGEMA_signal_9419 ), .Q ( new_AGEMA_signal_9420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4939 ( .C ( clk ), .D ( new_AGEMA_signal_9427 ), .Q ( new_AGEMA_signal_9428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4943 ( .C ( clk ), .D ( new_AGEMA_signal_9431 ), .Q ( new_AGEMA_signal_9432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4947 ( .C ( clk ), .D ( new_AGEMA_signal_9435 ), .Q ( new_AGEMA_signal_9436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4951 ( .C ( clk ), .D ( new_AGEMA_signal_9439 ), .Q ( new_AGEMA_signal_9440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4957 ( .C ( clk ), .D ( new_AGEMA_signal_9445 ), .Q ( new_AGEMA_signal_9446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4965 ( .C ( clk ), .D ( new_AGEMA_signal_9453 ), .Q ( new_AGEMA_signal_9454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4973 ( .C ( clk ), .D ( new_AGEMA_signal_9461 ), .Q ( new_AGEMA_signal_9462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4985 ( .C ( clk ), .D ( new_AGEMA_signal_9473 ), .Q ( new_AGEMA_signal_9474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4997 ( .C ( clk ), .D ( new_AGEMA_signal_9485 ), .Q ( new_AGEMA_signal_9486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5009 ( .C ( clk ), .D ( new_AGEMA_signal_9497 ), .Q ( new_AGEMA_signal_9498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5023 ( .C ( clk ), .D ( new_AGEMA_signal_9511 ), .Q ( new_AGEMA_signal_9512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5037 ( .C ( clk ), .D ( new_AGEMA_signal_9525 ), .Q ( new_AGEMA_signal_9526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5051 ( .C ( clk ), .D ( new_AGEMA_signal_9539 ), .Q ( new_AGEMA_signal_9540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5059 ( .C ( clk ), .D ( new_AGEMA_signal_9547 ), .Q ( new_AGEMA_signal_9548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5067 ( .C ( clk ), .D ( new_AGEMA_signal_9555 ), .Q ( new_AGEMA_signal_9556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5075 ( .C ( clk ), .D ( new_AGEMA_signal_9563 ), .Q ( new_AGEMA_signal_9564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5089 ( .C ( clk ), .D ( new_AGEMA_signal_9577 ), .Q ( new_AGEMA_signal_9578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5103 ( .C ( clk ), .D ( new_AGEMA_signal_9591 ), .Q ( new_AGEMA_signal_9592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5117 ( .C ( clk ), .D ( new_AGEMA_signal_9605 ), .Q ( new_AGEMA_signal_9606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5125 ( .C ( clk ), .D ( new_AGEMA_signal_9613 ), .Q ( new_AGEMA_signal_9614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5133 ( .C ( clk ), .D ( new_AGEMA_signal_9621 ), .Q ( new_AGEMA_signal_9622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5141 ( .C ( clk ), .D ( new_AGEMA_signal_9629 ), .Q ( new_AGEMA_signal_9630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5149 ( .C ( clk ), .D ( new_AGEMA_signal_9637 ), .Q ( new_AGEMA_signal_9638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5157 ( .C ( clk ), .D ( new_AGEMA_signal_9645 ), .Q ( new_AGEMA_signal_9646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5165 ( .C ( clk ), .D ( new_AGEMA_signal_9653 ), .Q ( new_AGEMA_signal_9654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5197 ( .C ( clk ), .D ( new_AGEMA_signal_9685 ), .Q ( new_AGEMA_signal_9686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5213 ( .C ( clk ), .D ( new_AGEMA_signal_9701 ), .Q ( new_AGEMA_signal_9702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5229 ( .C ( clk ), .D ( new_AGEMA_signal_9717 ), .Q ( new_AGEMA_signal_9718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5263 ( .C ( clk ), .D ( new_AGEMA_signal_9751 ), .Q ( new_AGEMA_signal_9752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5279 ( .C ( clk ), .D ( new_AGEMA_signal_9767 ), .Q ( new_AGEMA_signal_9768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5295 ( .C ( clk ), .D ( new_AGEMA_signal_9783 ), .Q ( new_AGEMA_signal_9784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5305 ( .C ( clk ), .D ( new_AGEMA_signal_9793 ), .Q ( new_AGEMA_signal_9794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5315 ( .C ( clk ), .D ( new_AGEMA_signal_9803 ), .Q ( new_AGEMA_signal_9804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5325 ( .C ( clk ), .D ( new_AGEMA_signal_9813 ), .Q ( new_AGEMA_signal_9814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5345 ( .C ( clk ), .D ( new_AGEMA_signal_9833 ), .Q ( new_AGEMA_signal_9834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5353 ( .C ( clk ), .D ( new_AGEMA_signal_9841 ), .Q ( new_AGEMA_signal_9842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5361 ( .C ( clk ), .D ( new_AGEMA_signal_9849 ), .Q ( new_AGEMA_signal_9850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5411 ( .C ( clk ), .D ( new_AGEMA_signal_9899 ), .Q ( new_AGEMA_signal_9900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5427 ( .C ( clk ), .D ( new_AGEMA_signal_9915 ), .Q ( new_AGEMA_signal_9916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5443 ( .C ( clk ), .D ( new_AGEMA_signal_9931 ), .Q ( new_AGEMA_signal_9932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5453 ( .C ( clk ), .D ( new_AGEMA_signal_9941 ), .Q ( new_AGEMA_signal_9942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5463 ( .C ( clk ), .D ( new_AGEMA_signal_9951 ), .Q ( new_AGEMA_signal_9952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5473 ( .C ( clk ), .D ( new_AGEMA_signal_9961 ), .Q ( new_AGEMA_signal_9962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5491 ( .C ( clk ), .D ( new_AGEMA_signal_9979 ), .Q ( new_AGEMA_signal_9980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5509 ( .C ( clk ), .D ( new_AGEMA_signal_9997 ), .Q ( new_AGEMA_signal_9998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5527 ( .C ( clk ), .D ( new_AGEMA_signal_10015 ), .Q ( new_AGEMA_signal_10016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5547 ( .C ( clk ), .D ( n2671 ), .Q ( new_AGEMA_signal_10036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5555 ( .C ( clk ), .D ( new_AGEMA_signal_2640 ), .Q ( new_AGEMA_signal_10044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5563 ( .C ( clk ), .D ( new_AGEMA_signal_2641 ), .Q ( new_AGEMA_signal_10052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5641 ( .C ( clk ), .D ( new_AGEMA_signal_10129 ), .Q ( new_AGEMA_signal_10130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5661 ( .C ( clk ), .D ( new_AGEMA_signal_10149 ), .Q ( new_AGEMA_signal_10150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5681 ( .C ( clk ), .D ( new_AGEMA_signal_10169 ), .Q ( new_AGEMA_signal_10170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5715 ( .C ( clk ), .D ( n2380 ), .Q ( new_AGEMA_signal_10204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5727 ( .C ( clk ), .D ( new_AGEMA_signal_2630 ), .Q ( new_AGEMA_signal_10216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5739 ( .C ( clk ), .D ( new_AGEMA_signal_2631 ), .Q ( new_AGEMA_signal_10228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5751 ( .C ( clk ), .D ( n2382 ), .Q ( new_AGEMA_signal_10240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5765 ( .C ( clk ), .D ( new_AGEMA_signal_2628 ), .Q ( new_AGEMA_signal_10254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5779 ( .C ( clk ), .D ( new_AGEMA_signal_2629 ), .Q ( new_AGEMA_signal_10268 ) ) ;

    /* cells in depth 18 */
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2016 ( .a ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, n1941}), .b ({new_AGEMA_signal_8763, new_AGEMA_signal_8757, new_AGEMA_signal_8751}), .clk ( clk ), .r ({Fresh[2381], Fresh[2380], Fresh[2379]}), .c ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, n2019}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2060 ( .a ({new_AGEMA_signal_8781, new_AGEMA_signal_8775, new_AGEMA_signal_8769}), .b ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, n1960}), .clk ( clk ), .r ({Fresh[2384], Fresh[2383], Fresh[2382]}), .c ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, n2002}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2116 ( .a ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, n1988}), .b ({new_AGEMA_signal_8799, new_AGEMA_signal_8793, new_AGEMA_signal_8787}), .clk ( clk ), .r ({Fresh[2387], Fresh[2386], Fresh[2385]}), .c ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, n1989}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2154 ( .a ({new_AGEMA_signal_8811, new_AGEMA_signal_8807, new_AGEMA_signal_8803}), .b ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, n2015}), .clk ( clk ), .r ({Fresh[2390], Fresh[2389], Fresh[2388]}), .c ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, n2016}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2170 ( .a ({new_AGEMA_signal_8835, new_AGEMA_signal_8827, new_AGEMA_signal_8819}), .b ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, n2030}), .clk ( clk ), .r ({Fresh[2393], Fresh[2392], Fresh[2391]}), .c ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, n2038}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2201 ( .a ({new_AGEMA_signal_8853, new_AGEMA_signal_8847, new_AGEMA_signal_8841}), .b ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, n2053}), .clk ( clk ), .r ({Fresh[2396], Fresh[2395], Fresh[2394]}), .c ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, n2111}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2223 ( .a ({new_AGEMA_signal_8865, new_AGEMA_signal_8861, new_AGEMA_signal_8857}), .b ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, n2071}), .clk ( clk ), .r ({Fresh[2399], Fresh[2398], Fresh[2397]}), .c ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, n2079}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2263 ( .a ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, n2103}), .b ({new_AGEMA_signal_8889, new_AGEMA_signal_8881, new_AGEMA_signal_8873}), .clk ( clk ), .r ({Fresh[2402], Fresh[2401], Fresh[2400]}), .c ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, n2104}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2289 ( .a ({new_AGEMA_signal_8913, new_AGEMA_signal_8905, new_AGEMA_signal_8897}), .b ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, n2126}), .clk ( clk ), .r ({Fresh[2405], Fresh[2404], Fresh[2403]}), .c ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, n2127}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2315 ( .a ({new_AGEMA_signal_8811, new_AGEMA_signal_8807, new_AGEMA_signal_8803}), .b ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, n2146}), .clk ( clk ), .r ({Fresh[2408], Fresh[2407], Fresh[2406]}), .c ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, n2147}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2336 ( .a ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, n2173}), .b ({new_AGEMA_signal_8943, new_AGEMA_signal_8933, new_AGEMA_signal_8923}), .clk ( clk ), .r ({Fresh[2411], Fresh[2410], Fresh[2409]}), .c ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, n2208}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2352 ( .a ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, n2187}), .b ({new_AGEMA_signal_8967, new_AGEMA_signal_8959, new_AGEMA_signal_8951}), .clk ( clk ), .r ({Fresh[2414], Fresh[2413], Fresh[2412]}), .c ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, n2199}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2420 ( .a ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, n2256}), .b ({new_AGEMA_signal_8985, new_AGEMA_signal_8979, new_AGEMA_signal_8973}), .clk ( clk ), .r ({Fresh[2417], Fresh[2416], Fresh[2415]}), .c ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, n2257}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2442 ( .a ({new_AGEMA_signal_8997, new_AGEMA_signal_8993, new_AGEMA_signal_8989}), .b ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, n2275}), .clk ( clk ), .r ({Fresh[2420], Fresh[2419], Fresh[2418]}), .c ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, n2281}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2475 ( .a ({new_AGEMA_signal_9015, new_AGEMA_signal_9009, new_AGEMA_signal_9003}), .b ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, n2303}), .clk ( clk ), .r ({Fresh[2423], Fresh[2422], Fresh[2421]}), .c ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, n2305}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2532 ( .a ({new_AGEMA_signal_9039, new_AGEMA_signal_9031, new_AGEMA_signal_9023}), .b ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, n2366}), .clk ( clk ), .r ({Fresh[2426], Fresh[2425], Fresh[2424]}), .c ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, n2368}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2583 ( .a ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, n2425}), .b ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, n2424}), .clk ( clk ), .r ({Fresh[2429], Fresh[2428], Fresh[2427]}), .c ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, n2426}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2605 ( .a ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, n2451}), .b ({new_AGEMA_signal_9057, new_AGEMA_signal_9051, new_AGEMA_signal_9045}), .clk ( clk ), .r ({Fresh[2432], Fresh[2431], Fresh[2430]}), .c ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, n2457}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2659 ( .a ({new_AGEMA_signal_9063, new_AGEMA_signal_9061, new_AGEMA_signal_9059}), .b ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, n2511}), .clk ( clk ), .r ({Fresh[2435], Fresh[2434], Fresh[2433]}), .c ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, n2513}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2717 ( .a ({new_AGEMA_signal_9087, new_AGEMA_signal_9079, new_AGEMA_signal_9071}), .b ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, n2590}), .clk ( clk ), .r ({Fresh[2438], Fresh[2437], Fresh[2436]}), .c ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, n2592}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2741 ( .a ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, n2623}), .b ({new_AGEMA_signal_9099, new_AGEMA_signal_9095, new_AGEMA_signal_9091}), .clk ( clk ), .r ({Fresh[2441], Fresh[2440], Fresh[2439]}), .c ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, n2637}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2767 ( .a ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, n2667}), .b ({new_AGEMA_signal_9117, new_AGEMA_signal_9111, new_AGEMA_signal_9105}), .clk ( clk ), .r ({Fresh[2444], Fresh[2443], Fresh[2442]}), .c ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, n2668}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2787 ( .a ({new_AGEMA_signal_9135, new_AGEMA_signal_9129, new_AGEMA_signal_9123}), .b ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, n2703}), .clk ( clk ), .r ({Fresh[2447], Fresh[2446], Fresh[2445]}), .c ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, n2705}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2841 ( .a ({new_AGEMA_signal_9147, new_AGEMA_signal_9143, new_AGEMA_signal_9139}), .b ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, n2803}), .clk ( clk ), .r ({Fresh[2450], Fresh[2449], Fresh[2448]}), .c ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, n2805}) ) ;
    buf_clk new_AGEMA_reg_buffer_4664 ( .C ( clk ), .D ( new_AGEMA_signal_9152 ), .Q ( new_AGEMA_signal_9153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4670 ( .C ( clk ), .D ( new_AGEMA_signal_9158 ), .Q ( new_AGEMA_signal_9159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4676 ( .C ( clk ), .D ( new_AGEMA_signal_9164 ), .Q ( new_AGEMA_signal_9165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4680 ( .C ( clk ), .D ( new_AGEMA_signal_9168 ), .Q ( new_AGEMA_signal_9169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4684 ( .C ( clk ), .D ( new_AGEMA_signal_9172 ), .Q ( new_AGEMA_signal_9173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4688 ( .C ( clk ), .D ( new_AGEMA_signal_9176 ), .Q ( new_AGEMA_signal_9177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4694 ( .C ( clk ), .D ( new_AGEMA_signal_9182 ), .Q ( new_AGEMA_signal_9183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4700 ( .C ( clk ), .D ( new_AGEMA_signal_9188 ), .Q ( new_AGEMA_signal_9189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4706 ( .C ( clk ), .D ( new_AGEMA_signal_9194 ), .Q ( new_AGEMA_signal_9195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4716 ( .C ( clk ), .D ( new_AGEMA_signal_9204 ), .Q ( new_AGEMA_signal_9205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4726 ( .C ( clk ), .D ( new_AGEMA_signal_9214 ), .Q ( new_AGEMA_signal_9215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4736 ( .C ( clk ), .D ( new_AGEMA_signal_9224 ), .Q ( new_AGEMA_signal_9225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4742 ( .C ( clk ), .D ( new_AGEMA_signal_9230 ), .Q ( new_AGEMA_signal_9231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4748 ( .C ( clk ), .D ( new_AGEMA_signal_9236 ), .Q ( new_AGEMA_signal_9237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4754 ( .C ( clk ), .D ( new_AGEMA_signal_9242 ), .Q ( new_AGEMA_signal_9243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4760 ( .C ( clk ), .D ( new_AGEMA_signal_9248 ), .Q ( new_AGEMA_signal_9249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4766 ( .C ( clk ), .D ( new_AGEMA_signal_9254 ), .Q ( new_AGEMA_signal_9255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4772 ( .C ( clk ), .D ( new_AGEMA_signal_9260 ), .Q ( new_AGEMA_signal_9261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4776 ( .C ( clk ), .D ( new_AGEMA_signal_9264 ), .Q ( new_AGEMA_signal_9265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4780 ( .C ( clk ), .D ( new_AGEMA_signal_9268 ), .Q ( new_AGEMA_signal_9269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4784 ( .C ( clk ), .D ( new_AGEMA_signal_9272 ), .Q ( new_AGEMA_signal_9273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4788 ( .C ( clk ), .D ( new_AGEMA_signal_9276 ), .Q ( new_AGEMA_signal_9277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4792 ( .C ( clk ), .D ( new_AGEMA_signal_9280 ), .Q ( new_AGEMA_signal_9281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4796 ( .C ( clk ), .D ( new_AGEMA_signal_9284 ), .Q ( new_AGEMA_signal_9285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4804 ( .C ( clk ), .D ( new_AGEMA_signal_9292 ), .Q ( new_AGEMA_signal_9293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4812 ( .C ( clk ), .D ( new_AGEMA_signal_9300 ), .Q ( new_AGEMA_signal_9301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4820 ( .C ( clk ), .D ( new_AGEMA_signal_9308 ), .Q ( new_AGEMA_signal_9309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4826 ( .C ( clk ), .D ( new_AGEMA_signal_9314 ), .Q ( new_AGEMA_signal_9315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4832 ( .C ( clk ), .D ( new_AGEMA_signal_9320 ), .Q ( new_AGEMA_signal_9321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4838 ( .C ( clk ), .D ( new_AGEMA_signal_9326 ), .Q ( new_AGEMA_signal_9327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4846 ( .C ( clk ), .D ( new_AGEMA_signal_9334 ), .Q ( new_AGEMA_signal_9335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4854 ( .C ( clk ), .D ( new_AGEMA_signal_9342 ), .Q ( new_AGEMA_signal_9343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4862 ( .C ( clk ), .D ( new_AGEMA_signal_9350 ), .Q ( new_AGEMA_signal_9351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4870 ( .C ( clk ), .D ( new_AGEMA_signal_9358 ), .Q ( new_AGEMA_signal_9359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4878 ( .C ( clk ), .D ( new_AGEMA_signal_9366 ), .Q ( new_AGEMA_signal_9367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4886 ( .C ( clk ), .D ( new_AGEMA_signal_9374 ), .Q ( new_AGEMA_signal_9375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4888 ( .C ( clk ), .D ( new_AGEMA_signal_9376 ), .Q ( new_AGEMA_signal_9377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4890 ( .C ( clk ), .D ( new_AGEMA_signal_9378 ), .Q ( new_AGEMA_signal_9379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4892 ( .C ( clk ), .D ( new_AGEMA_signal_9380 ), .Q ( new_AGEMA_signal_9381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4896 ( .C ( clk ), .D ( new_AGEMA_signal_9384 ), .Q ( new_AGEMA_signal_9385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4900 ( .C ( clk ), .D ( new_AGEMA_signal_9388 ), .Q ( new_AGEMA_signal_9389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4904 ( .C ( clk ), .D ( new_AGEMA_signal_9392 ), .Q ( new_AGEMA_signal_9393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4908 ( .C ( clk ), .D ( new_AGEMA_signal_9396 ), .Q ( new_AGEMA_signal_9397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4912 ( .C ( clk ), .D ( new_AGEMA_signal_9400 ), .Q ( new_AGEMA_signal_9401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4916 ( .C ( clk ), .D ( new_AGEMA_signal_9404 ), .Q ( new_AGEMA_signal_9405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4924 ( .C ( clk ), .D ( new_AGEMA_signal_9412 ), .Q ( new_AGEMA_signal_9413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4932 ( .C ( clk ), .D ( new_AGEMA_signal_9420 ), .Q ( new_AGEMA_signal_9421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4940 ( .C ( clk ), .D ( new_AGEMA_signal_9428 ), .Q ( new_AGEMA_signal_9429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4944 ( .C ( clk ), .D ( new_AGEMA_signal_9432 ), .Q ( new_AGEMA_signal_9433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4948 ( .C ( clk ), .D ( new_AGEMA_signal_9436 ), .Q ( new_AGEMA_signal_9437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4952 ( .C ( clk ), .D ( new_AGEMA_signal_9440 ), .Q ( new_AGEMA_signal_9441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4958 ( .C ( clk ), .D ( new_AGEMA_signal_9446 ), .Q ( new_AGEMA_signal_9447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4966 ( .C ( clk ), .D ( new_AGEMA_signal_9454 ), .Q ( new_AGEMA_signal_9455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4974 ( .C ( clk ), .D ( new_AGEMA_signal_9462 ), .Q ( new_AGEMA_signal_9463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4986 ( .C ( clk ), .D ( new_AGEMA_signal_9474 ), .Q ( new_AGEMA_signal_9475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4998 ( .C ( clk ), .D ( new_AGEMA_signal_9486 ), .Q ( new_AGEMA_signal_9487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5010 ( .C ( clk ), .D ( new_AGEMA_signal_9498 ), .Q ( new_AGEMA_signal_9499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5024 ( .C ( clk ), .D ( new_AGEMA_signal_9512 ), .Q ( new_AGEMA_signal_9513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5038 ( .C ( clk ), .D ( new_AGEMA_signal_9526 ), .Q ( new_AGEMA_signal_9527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5052 ( .C ( clk ), .D ( new_AGEMA_signal_9540 ), .Q ( new_AGEMA_signal_9541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5060 ( .C ( clk ), .D ( new_AGEMA_signal_9548 ), .Q ( new_AGEMA_signal_9549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5068 ( .C ( clk ), .D ( new_AGEMA_signal_9556 ), .Q ( new_AGEMA_signal_9557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5076 ( .C ( clk ), .D ( new_AGEMA_signal_9564 ), .Q ( new_AGEMA_signal_9565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5090 ( .C ( clk ), .D ( new_AGEMA_signal_9578 ), .Q ( new_AGEMA_signal_9579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5104 ( .C ( clk ), .D ( new_AGEMA_signal_9592 ), .Q ( new_AGEMA_signal_9593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5118 ( .C ( clk ), .D ( new_AGEMA_signal_9606 ), .Q ( new_AGEMA_signal_9607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5126 ( .C ( clk ), .D ( new_AGEMA_signal_9614 ), .Q ( new_AGEMA_signal_9615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5134 ( .C ( clk ), .D ( new_AGEMA_signal_9622 ), .Q ( new_AGEMA_signal_9623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5142 ( .C ( clk ), .D ( new_AGEMA_signal_9630 ), .Q ( new_AGEMA_signal_9631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5150 ( .C ( clk ), .D ( new_AGEMA_signal_9638 ), .Q ( new_AGEMA_signal_9639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5158 ( .C ( clk ), .D ( new_AGEMA_signal_9646 ), .Q ( new_AGEMA_signal_9647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5166 ( .C ( clk ), .D ( new_AGEMA_signal_9654 ), .Q ( new_AGEMA_signal_9655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5198 ( .C ( clk ), .D ( new_AGEMA_signal_9686 ), .Q ( new_AGEMA_signal_9687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5214 ( .C ( clk ), .D ( new_AGEMA_signal_9702 ), .Q ( new_AGEMA_signal_9703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5230 ( .C ( clk ), .D ( new_AGEMA_signal_9718 ), .Q ( new_AGEMA_signal_9719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5264 ( .C ( clk ), .D ( new_AGEMA_signal_9752 ), .Q ( new_AGEMA_signal_9753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5280 ( .C ( clk ), .D ( new_AGEMA_signal_9768 ), .Q ( new_AGEMA_signal_9769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5296 ( .C ( clk ), .D ( new_AGEMA_signal_9784 ), .Q ( new_AGEMA_signal_9785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5306 ( .C ( clk ), .D ( new_AGEMA_signal_9794 ), .Q ( new_AGEMA_signal_9795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5316 ( .C ( clk ), .D ( new_AGEMA_signal_9804 ), .Q ( new_AGEMA_signal_9805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5326 ( .C ( clk ), .D ( new_AGEMA_signal_9814 ), .Q ( new_AGEMA_signal_9815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5346 ( .C ( clk ), .D ( new_AGEMA_signal_9834 ), .Q ( new_AGEMA_signal_9835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5354 ( .C ( clk ), .D ( new_AGEMA_signal_9842 ), .Q ( new_AGEMA_signal_9843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5362 ( .C ( clk ), .D ( new_AGEMA_signal_9850 ), .Q ( new_AGEMA_signal_9851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5412 ( .C ( clk ), .D ( new_AGEMA_signal_9900 ), .Q ( new_AGEMA_signal_9901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5428 ( .C ( clk ), .D ( new_AGEMA_signal_9916 ), .Q ( new_AGEMA_signal_9917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5444 ( .C ( clk ), .D ( new_AGEMA_signal_9932 ), .Q ( new_AGEMA_signal_9933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5454 ( .C ( clk ), .D ( new_AGEMA_signal_9942 ), .Q ( new_AGEMA_signal_9943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5464 ( .C ( clk ), .D ( new_AGEMA_signal_9952 ), .Q ( new_AGEMA_signal_9953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5474 ( .C ( clk ), .D ( new_AGEMA_signal_9962 ), .Q ( new_AGEMA_signal_9963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5492 ( .C ( clk ), .D ( new_AGEMA_signal_9980 ), .Q ( new_AGEMA_signal_9981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5510 ( .C ( clk ), .D ( new_AGEMA_signal_9998 ), .Q ( new_AGEMA_signal_9999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5528 ( .C ( clk ), .D ( new_AGEMA_signal_10016 ), .Q ( new_AGEMA_signal_10017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5548 ( .C ( clk ), .D ( new_AGEMA_signal_10036 ), .Q ( new_AGEMA_signal_10037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5556 ( .C ( clk ), .D ( new_AGEMA_signal_10044 ), .Q ( new_AGEMA_signal_10045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5564 ( .C ( clk ), .D ( new_AGEMA_signal_10052 ), .Q ( new_AGEMA_signal_10053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5642 ( .C ( clk ), .D ( new_AGEMA_signal_10130 ), .Q ( new_AGEMA_signal_10131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5662 ( .C ( clk ), .D ( new_AGEMA_signal_10150 ), .Q ( new_AGEMA_signal_10151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5682 ( .C ( clk ), .D ( new_AGEMA_signal_10170 ), .Q ( new_AGEMA_signal_10171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5716 ( .C ( clk ), .D ( new_AGEMA_signal_10204 ), .Q ( new_AGEMA_signal_10205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5728 ( .C ( clk ), .D ( new_AGEMA_signal_10216 ), .Q ( new_AGEMA_signal_10217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5740 ( .C ( clk ), .D ( new_AGEMA_signal_10228 ), .Q ( new_AGEMA_signal_10229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5752 ( .C ( clk ), .D ( new_AGEMA_signal_10240 ), .Q ( new_AGEMA_signal_10241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5766 ( .C ( clk ), .D ( new_AGEMA_signal_10254 ), .Q ( new_AGEMA_signal_10255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5780 ( .C ( clk ), .D ( new_AGEMA_signal_10268 ), .Q ( new_AGEMA_signal_10269 ) ) ;

    /* cells in depth 19 */
    buf_clk new_AGEMA_reg_buffer_4959 ( .C ( clk ), .D ( new_AGEMA_signal_9447 ), .Q ( new_AGEMA_signal_9448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4967 ( .C ( clk ), .D ( new_AGEMA_signal_9455 ), .Q ( new_AGEMA_signal_9456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4975 ( .C ( clk ), .D ( new_AGEMA_signal_9463 ), .Q ( new_AGEMA_signal_9464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4987 ( .C ( clk ), .D ( new_AGEMA_signal_9475 ), .Q ( new_AGEMA_signal_9476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4999 ( .C ( clk ), .D ( new_AGEMA_signal_9487 ), .Q ( new_AGEMA_signal_9488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5011 ( .C ( clk ), .D ( new_AGEMA_signal_9499 ), .Q ( new_AGEMA_signal_9500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5025 ( .C ( clk ), .D ( new_AGEMA_signal_9513 ), .Q ( new_AGEMA_signal_9514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5039 ( .C ( clk ), .D ( new_AGEMA_signal_9527 ), .Q ( new_AGEMA_signal_9528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5053 ( .C ( clk ), .D ( new_AGEMA_signal_9541 ), .Q ( new_AGEMA_signal_9542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5061 ( .C ( clk ), .D ( new_AGEMA_signal_9549 ), .Q ( new_AGEMA_signal_9550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5069 ( .C ( clk ), .D ( new_AGEMA_signal_9557 ), .Q ( new_AGEMA_signal_9558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5077 ( .C ( clk ), .D ( new_AGEMA_signal_9565 ), .Q ( new_AGEMA_signal_9566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5091 ( .C ( clk ), .D ( new_AGEMA_signal_9579 ), .Q ( new_AGEMA_signal_9580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5105 ( .C ( clk ), .D ( new_AGEMA_signal_9593 ), .Q ( new_AGEMA_signal_9594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5119 ( .C ( clk ), .D ( new_AGEMA_signal_9607 ), .Q ( new_AGEMA_signal_9608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5127 ( .C ( clk ), .D ( new_AGEMA_signal_9615 ), .Q ( new_AGEMA_signal_9616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5135 ( .C ( clk ), .D ( new_AGEMA_signal_9623 ), .Q ( new_AGEMA_signal_9624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5143 ( .C ( clk ), .D ( new_AGEMA_signal_9631 ), .Q ( new_AGEMA_signal_9632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5151 ( .C ( clk ), .D ( new_AGEMA_signal_9639 ), .Q ( new_AGEMA_signal_9640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5159 ( .C ( clk ), .D ( new_AGEMA_signal_9647 ), .Q ( new_AGEMA_signal_9648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5167 ( .C ( clk ), .D ( new_AGEMA_signal_9655 ), .Q ( new_AGEMA_signal_9656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5169 ( .C ( clk ), .D ( n2002 ), .Q ( new_AGEMA_signal_9658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5173 ( .C ( clk ), .D ( new_AGEMA_signal_2654 ), .Q ( new_AGEMA_signal_9662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5177 ( .C ( clk ), .D ( new_AGEMA_signal_2655 ), .Q ( new_AGEMA_signal_9666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5199 ( .C ( clk ), .D ( new_AGEMA_signal_9687 ), .Q ( new_AGEMA_signal_9688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5215 ( .C ( clk ), .D ( new_AGEMA_signal_9703 ), .Q ( new_AGEMA_signal_9704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5231 ( .C ( clk ), .D ( new_AGEMA_signal_9719 ), .Q ( new_AGEMA_signal_9720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5235 ( .C ( clk ), .D ( n2208 ), .Q ( new_AGEMA_signal_9724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5239 ( .C ( clk ), .D ( new_AGEMA_signal_2672 ), .Q ( new_AGEMA_signal_9728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5243 ( .C ( clk ), .D ( new_AGEMA_signal_2673 ), .Q ( new_AGEMA_signal_9732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5265 ( .C ( clk ), .D ( new_AGEMA_signal_9753 ), .Q ( new_AGEMA_signal_9754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5281 ( .C ( clk ), .D ( new_AGEMA_signal_9769 ), .Q ( new_AGEMA_signal_9770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5297 ( .C ( clk ), .D ( new_AGEMA_signal_9785 ), .Q ( new_AGEMA_signal_9786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5307 ( .C ( clk ), .D ( new_AGEMA_signal_9795 ), .Q ( new_AGEMA_signal_9796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5317 ( .C ( clk ), .D ( new_AGEMA_signal_9805 ), .Q ( new_AGEMA_signal_9806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5327 ( .C ( clk ), .D ( new_AGEMA_signal_9815 ), .Q ( new_AGEMA_signal_9816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5331 ( .C ( clk ), .D ( n2668 ), .Q ( new_AGEMA_signal_9820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5335 ( .C ( clk ), .D ( new_AGEMA_signal_2694 ), .Q ( new_AGEMA_signal_9824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5339 ( .C ( clk ), .D ( new_AGEMA_signal_2695 ), .Q ( new_AGEMA_signal_9828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5347 ( .C ( clk ), .D ( new_AGEMA_signal_9835 ), .Q ( new_AGEMA_signal_9836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5355 ( .C ( clk ), .D ( new_AGEMA_signal_9843 ), .Q ( new_AGEMA_signal_9844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5363 ( .C ( clk ), .D ( new_AGEMA_signal_9851 ), .Q ( new_AGEMA_signal_9852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5367 ( .C ( clk ), .D ( n2016 ), .Q ( new_AGEMA_signal_9856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5373 ( .C ( clk ), .D ( new_AGEMA_signal_2658 ), .Q ( new_AGEMA_signal_9862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5379 ( .C ( clk ), .D ( new_AGEMA_signal_2659 ), .Q ( new_AGEMA_signal_9868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5385 ( .C ( clk ), .D ( n2111 ), .Q ( new_AGEMA_signal_9874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5391 ( .C ( clk ), .D ( new_AGEMA_signal_2662 ), .Q ( new_AGEMA_signal_9880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5397 ( .C ( clk ), .D ( new_AGEMA_signal_2663 ), .Q ( new_AGEMA_signal_9886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5413 ( .C ( clk ), .D ( new_AGEMA_signal_9901 ), .Q ( new_AGEMA_signal_9902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5429 ( .C ( clk ), .D ( new_AGEMA_signal_9917 ), .Q ( new_AGEMA_signal_9918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5445 ( .C ( clk ), .D ( new_AGEMA_signal_9933 ), .Q ( new_AGEMA_signal_9934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5455 ( .C ( clk ), .D ( new_AGEMA_signal_9943 ), .Q ( new_AGEMA_signal_9944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5465 ( .C ( clk ), .D ( new_AGEMA_signal_9953 ), .Q ( new_AGEMA_signal_9954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5475 ( .C ( clk ), .D ( new_AGEMA_signal_9963 ), .Q ( new_AGEMA_signal_9964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5493 ( .C ( clk ), .D ( new_AGEMA_signal_9981 ), .Q ( new_AGEMA_signal_9982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5511 ( .C ( clk ), .D ( new_AGEMA_signal_9999 ), .Q ( new_AGEMA_signal_10000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5529 ( .C ( clk ), .D ( new_AGEMA_signal_10017 ), .Q ( new_AGEMA_signal_10018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5549 ( .C ( clk ), .D ( new_AGEMA_signal_10037 ), .Q ( new_AGEMA_signal_10038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5557 ( .C ( clk ), .D ( new_AGEMA_signal_10045 ), .Q ( new_AGEMA_signal_10046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5565 ( .C ( clk ), .D ( new_AGEMA_signal_10053 ), .Q ( new_AGEMA_signal_10054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5583 ( .C ( clk ), .D ( n2019 ), .Q ( new_AGEMA_signal_10072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5591 ( .C ( clk ), .D ( new_AGEMA_signal_2652 ), .Q ( new_AGEMA_signal_10080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5599 ( .C ( clk ), .D ( new_AGEMA_signal_2653 ), .Q ( new_AGEMA_signal_10088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5643 ( .C ( clk ), .D ( new_AGEMA_signal_10131 ), .Q ( new_AGEMA_signal_10132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5663 ( .C ( clk ), .D ( new_AGEMA_signal_10151 ), .Q ( new_AGEMA_signal_10152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5683 ( .C ( clk ), .D ( new_AGEMA_signal_10171 ), .Q ( new_AGEMA_signal_10172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5717 ( .C ( clk ), .D ( new_AGEMA_signal_10205 ), .Q ( new_AGEMA_signal_10206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5729 ( .C ( clk ), .D ( new_AGEMA_signal_10217 ), .Q ( new_AGEMA_signal_10218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5741 ( .C ( clk ), .D ( new_AGEMA_signal_10229 ), .Q ( new_AGEMA_signal_10230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5753 ( .C ( clk ), .D ( new_AGEMA_signal_10241 ), .Q ( new_AGEMA_signal_10242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5767 ( .C ( clk ), .D ( new_AGEMA_signal_10255 ), .Q ( new_AGEMA_signal_10256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5781 ( .C ( clk ), .D ( new_AGEMA_signal_10269 ), .Q ( new_AGEMA_signal_10270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5793 ( .C ( clk ), .D ( n2426 ), .Q ( new_AGEMA_signal_10282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5807 ( .C ( clk ), .D ( new_AGEMA_signal_2684 ), .Q ( new_AGEMA_signal_10296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5821 ( .C ( clk ), .D ( new_AGEMA_signal_2685 ), .Q ( new_AGEMA_signal_10310 ) ) ;

    /* cells in depth 20 */
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2117 ( .a ({new_AGEMA_signal_9165, new_AGEMA_signal_9159, new_AGEMA_signal_9153}), .b ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, n1989}), .clk ( clk ), .r ({Fresh[2453], Fresh[2452], Fresh[2451]}), .c ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, n2000}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2181 ( .a ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, n2038}), .b ({new_AGEMA_signal_9177, new_AGEMA_signal_9173, new_AGEMA_signal_9169}), .clk ( clk ), .r ({Fresh[2456], Fresh[2455], Fresh[2454]}), .c ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, n2113}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2231 ( .a ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, n2079}), .b ({new_AGEMA_signal_9195, new_AGEMA_signal_9189, new_AGEMA_signal_9183}), .clk ( clk ), .r ({Fresh[2459], Fresh[2458], Fresh[2457]}), .c ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, n2109}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2264 ( .a ({new_AGEMA_signal_9225, new_AGEMA_signal_9215, new_AGEMA_signal_9205}), .b ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, n2104}), .clk ( clk ), .r ({Fresh[2462], Fresh[2461], Fresh[2460]}), .c ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, n2107}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2290 ( .a ({new_AGEMA_signal_9243, new_AGEMA_signal_9237, new_AGEMA_signal_9231}), .b ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, n2127}), .clk ( clk ), .r ({Fresh[2465], Fresh[2464], Fresh[2463]}), .c ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, n2212}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2316 ( .a ({new_AGEMA_signal_9261, new_AGEMA_signal_9255, new_AGEMA_signal_9249}), .b ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, n2147}), .clk ( clk ), .r ({Fresh[2468], Fresh[2467], Fresh[2466]}), .c ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, n2149}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2366 ( .a ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, n2199}), .b ({new_AGEMA_signal_9273, new_AGEMA_signal_9269, new_AGEMA_signal_9265}), .clk ( clk ), .r ({Fresh[2471], Fresh[2470], Fresh[2469]}), .c ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, n2206}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2421 ( .a ({new_AGEMA_signal_9285, new_AGEMA_signal_9281, new_AGEMA_signal_9277}), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, n2257}), .clk ( clk ), .r ({Fresh[2474], Fresh[2473], Fresh[2472]}), .c ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, n2310}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2447 ( .a ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, n2281}), .b ({new_AGEMA_signal_9309, new_AGEMA_signal_9301, new_AGEMA_signal_9293}), .clk ( clk ), .r ({Fresh[2477], Fresh[2476], Fresh[2475]}), .c ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, n2308}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2476 ( .a ({new_AGEMA_signal_9327, new_AGEMA_signal_9321, new_AGEMA_signal_9315}), .b ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, n2305}), .clk ( clk ), .r ({Fresh[2480], Fresh[2479], Fresh[2478]}), .c ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, n2307}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2533 ( .a ({new_AGEMA_signal_9351, new_AGEMA_signal_9343, new_AGEMA_signal_9335}), .b ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, n2368}), .clk ( clk ), .r ({Fresh[2483], Fresh[2482], Fresh[2481]}), .c ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, n2370}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2611 ( .a ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, n2457}), .b ({new_AGEMA_signal_9375, new_AGEMA_signal_9367, new_AGEMA_signal_9359}), .clk ( clk ), .r ({Fresh[2486], Fresh[2485], Fresh[2484]}), .c ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, n2530}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2660 ( .a ({new_AGEMA_signal_9381, new_AGEMA_signal_9379, new_AGEMA_signal_9377}), .b ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, n2513}), .clk ( clk ), .r ({Fresh[2489], Fresh[2488], Fresh[2487]}), .c ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, n2515}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2718 ( .a ({new_AGEMA_signal_9393, new_AGEMA_signal_9389, new_AGEMA_signal_9385}), .b ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, n2592}), .clk ( clk ), .r ({Fresh[2492], Fresh[2491], Fresh[2490]}), .c ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, n2639}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2749 ( .a ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, n2637}), .b ({new_AGEMA_signal_9405, new_AGEMA_signal_9401, new_AGEMA_signal_9397}), .clk ( clk ), .r ({Fresh[2495], Fresh[2494], Fresh[2493]}), .c ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, n2638}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2788 ( .a ({new_AGEMA_signal_9429, new_AGEMA_signal_9421, new_AGEMA_signal_9413}), .b ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, n2705}), .clk ( clk ), .r ({Fresh[2498], Fresh[2497], Fresh[2496]}), .c ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, n2832}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2842 ( .a ({new_AGEMA_signal_9441, new_AGEMA_signal_9437, new_AGEMA_signal_9433}), .b ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, n2805}), .clk ( clk ), .r ({Fresh[2501], Fresh[2500], Fresh[2499]}), .c ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, n2807}) ) ;
    buf_clk new_AGEMA_reg_buffer_4960 ( .C ( clk ), .D ( new_AGEMA_signal_9448 ), .Q ( new_AGEMA_signal_9449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4968 ( .C ( clk ), .D ( new_AGEMA_signal_9456 ), .Q ( new_AGEMA_signal_9457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4976 ( .C ( clk ), .D ( new_AGEMA_signal_9464 ), .Q ( new_AGEMA_signal_9465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4988 ( .C ( clk ), .D ( new_AGEMA_signal_9476 ), .Q ( new_AGEMA_signal_9477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5000 ( .C ( clk ), .D ( new_AGEMA_signal_9488 ), .Q ( new_AGEMA_signal_9489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5012 ( .C ( clk ), .D ( new_AGEMA_signal_9500 ), .Q ( new_AGEMA_signal_9501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5026 ( .C ( clk ), .D ( new_AGEMA_signal_9514 ), .Q ( new_AGEMA_signal_9515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5040 ( .C ( clk ), .D ( new_AGEMA_signal_9528 ), .Q ( new_AGEMA_signal_9529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5054 ( .C ( clk ), .D ( new_AGEMA_signal_9542 ), .Q ( new_AGEMA_signal_9543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5062 ( .C ( clk ), .D ( new_AGEMA_signal_9550 ), .Q ( new_AGEMA_signal_9551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5070 ( .C ( clk ), .D ( new_AGEMA_signal_9558 ), .Q ( new_AGEMA_signal_9559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5078 ( .C ( clk ), .D ( new_AGEMA_signal_9566 ), .Q ( new_AGEMA_signal_9567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5092 ( .C ( clk ), .D ( new_AGEMA_signal_9580 ), .Q ( new_AGEMA_signal_9581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5106 ( .C ( clk ), .D ( new_AGEMA_signal_9594 ), .Q ( new_AGEMA_signal_9595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5120 ( .C ( clk ), .D ( new_AGEMA_signal_9608 ), .Q ( new_AGEMA_signal_9609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5128 ( .C ( clk ), .D ( new_AGEMA_signal_9616 ), .Q ( new_AGEMA_signal_9617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5136 ( .C ( clk ), .D ( new_AGEMA_signal_9624 ), .Q ( new_AGEMA_signal_9625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5144 ( .C ( clk ), .D ( new_AGEMA_signal_9632 ), .Q ( new_AGEMA_signal_9633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5152 ( .C ( clk ), .D ( new_AGEMA_signal_9640 ), .Q ( new_AGEMA_signal_9641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5160 ( .C ( clk ), .D ( new_AGEMA_signal_9648 ), .Q ( new_AGEMA_signal_9649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5168 ( .C ( clk ), .D ( new_AGEMA_signal_9656 ), .Q ( new_AGEMA_signal_9657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5170 ( .C ( clk ), .D ( new_AGEMA_signal_9658 ), .Q ( new_AGEMA_signal_9659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5174 ( .C ( clk ), .D ( new_AGEMA_signal_9662 ), .Q ( new_AGEMA_signal_9663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5178 ( .C ( clk ), .D ( new_AGEMA_signal_9666 ), .Q ( new_AGEMA_signal_9667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5200 ( .C ( clk ), .D ( new_AGEMA_signal_9688 ), .Q ( new_AGEMA_signal_9689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5216 ( .C ( clk ), .D ( new_AGEMA_signal_9704 ), .Q ( new_AGEMA_signal_9705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5232 ( .C ( clk ), .D ( new_AGEMA_signal_9720 ), .Q ( new_AGEMA_signal_9721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5236 ( .C ( clk ), .D ( new_AGEMA_signal_9724 ), .Q ( new_AGEMA_signal_9725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5240 ( .C ( clk ), .D ( new_AGEMA_signal_9728 ), .Q ( new_AGEMA_signal_9729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5244 ( .C ( clk ), .D ( new_AGEMA_signal_9732 ), .Q ( new_AGEMA_signal_9733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5266 ( .C ( clk ), .D ( new_AGEMA_signal_9754 ), .Q ( new_AGEMA_signal_9755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5282 ( .C ( clk ), .D ( new_AGEMA_signal_9770 ), .Q ( new_AGEMA_signal_9771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5298 ( .C ( clk ), .D ( new_AGEMA_signal_9786 ), .Q ( new_AGEMA_signal_9787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5308 ( .C ( clk ), .D ( new_AGEMA_signal_9796 ), .Q ( new_AGEMA_signal_9797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5318 ( .C ( clk ), .D ( new_AGEMA_signal_9806 ), .Q ( new_AGEMA_signal_9807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5328 ( .C ( clk ), .D ( new_AGEMA_signal_9816 ), .Q ( new_AGEMA_signal_9817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5332 ( .C ( clk ), .D ( new_AGEMA_signal_9820 ), .Q ( new_AGEMA_signal_9821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5336 ( .C ( clk ), .D ( new_AGEMA_signal_9824 ), .Q ( new_AGEMA_signal_9825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5340 ( .C ( clk ), .D ( new_AGEMA_signal_9828 ), .Q ( new_AGEMA_signal_9829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5348 ( .C ( clk ), .D ( new_AGEMA_signal_9836 ), .Q ( new_AGEMA_signal_9837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5356 ( .C ( clk ), .D ( new_AGEMA_signal_9844 ), .Q ( new_AGEMA_signal_9845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5364 ( .C ( clk ), .D ( new_AGEMA_signal_9852 ), .Q ( new_AGEMA_signal_9853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5368 ( .C ( clk ), .D ( new_AGEMA_signal_9856 ), .Q ( new_AGEMA_signal_9857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5374 ( .C ( clk ), .D ( new_AGEMA_signal_9862 ), .Q ( new_AGEMA_signal_9863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5380 ( .C ( clk ), .D ( new_AGEMA_signal_9868 ), .Q ( new_AGEMA_signal_9869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5386 ( .C ( clk ), .D ( new_AGEMA_signal_9874 ), .Q ( new_AGEMA_signal_9875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5392 ( .C ( clk ), .D ( new_AGEMA_signal_9880 ), .Q ( new_AGEMA_signal_9881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5398 ( .C ( clk ), .D ( new_AGEMA_signal_9886 ), .Q ( new_AGEMA_signal_9887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5414 ( .C ( clk ), .D ( new_AGEMA_signal_9902 ), .Q ( new_AGEMA_signal_9903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5430 ( .C ( clk ), .D ( new_AGEMA_signal_9918 ), .Q ( new_AGEMA_signal_9919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5446 ( .C ( clk ), .D ( new_AGEMA_signal_9934 ), .Q ( new_AGEMA_signal_9935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5456 ( .C ( clk ), .D ( new_AGEMA_signal_9944 ), .Q ( new_AGEMA_signal_9945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5466 ( .C ( clk ), .D ( new_AGEMA_signal_9954 ), .Q ( new_AGEMA_signal_9955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5476 ( .C ( clk ), .D ( new_AGEMA_signal_9964 ), .Q ( new_AGEMA_signal_9965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5494 ( .C ( clk ), .D ( new_AGEMA_signal_9982 ), .Q ( new_AGEMA_signal_9983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5512 ( .C ( clk ), .D ( new_AGEMA_signal_10000 ), .Q ( new_AGEMA_signal_10001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5530 ( .C ( clk ), .D ( new_AGEMA_signal_10018 ), .Q ( new_AGEMA_signal_10019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5550 ( .C ( clk ), .D ( new_AGEMA_signal_10038 ), .Q ( new_AGEMA_signal_10039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5558 ( .C ( clk ), .D ( new_AGEMA_signal_10046 ), .Q ( new_AGEMA_signal_10047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5566 ( .C ( clk ), .D ( new_AGEMA_signal_10054 ), .Q ( new_AGEMA_signal_10055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5584 ( .C ( clk ), .D ( new_AGEMA_signal_10072 ), .Q ( new_AGEMA_signal_10073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5592 ( .C ( clk ), .D ( new_AGEMA_signal_10080 ), .Q ( new_AGEMA_signal_10081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5600 ( .C ( clk ), .D ( new_AGEMA_signal_10088 ), .Q ( new_AGEMA_signal_10089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5644 ( .C ( clk ), .D ( new_AGEMA_signal_10132 ), .Q ( new_AGEMA_signal_10133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5664 ( .C ( clk ), .D ( new_AGEMA_signal_10152 ), .Q ( new_AGEMA_signal_10153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5684 ( .C ( clk ), .D ( new_AGEMA_signal_10172 ), .Q ( new_AGEMA_signal_10173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5718 ( .C ( clk ), .D ( new_AGEMA_signal_10206 ), .Q ( new_AGEMA_signal_10207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5730 ( .C ( clk ), .D ( new_AGEMA_signal_10218 ), .Q ( new_AGEMA_signal_10219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5742 ( .C ( clk ), .D ( new_AGEMA_signal_10230 ), .Q ( new_AGEMA_signal_10231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5754 ( .C ( clk ), .D ( new_AGEMA_signal_10242 ), .Q ( new_AGEMA_signal_10243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5768 ( .C ( clk ), .D ( new_AGEMA_signal_10256 ), .Q ( new_AGEMA_signal_10257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5782 ( .C ( clk ), .D ( new_AGEMA_signal_10270 ), .Q ( new_AGEMA_signal_10271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5794 ( .C ( clk ), .D ( new_AGEMA_signal_10282 ), .Q ( new_AGEMA_signal_10283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5808 ( .C ( clk ), .D ( new_AGEMA_signal_10296 ), .Q ( new_AGEMA_signal_10297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5822 ( .C ( clk ), .D ( new_AGEMA_signal_10310 ), .Q ( new_AGEMA_signal_10311 ) ) ;

    /* cells in depth 21 */
    buf_clk new_AGEMA_reg_buffer_5171 ( .C ( clk ), .D ( new_AGEMA_signal_9659 ), .Q ( new_AGEMA_signal_9660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5175 ( .C ( clk ), .D ( new_AGEMA_signal_9663 ), .Q ( new_AGEMA_signal_9664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5179 ( .C ( clk ), .D ( new_AGEMA_signal_9667 ), .Q ( new_AGEMA_signal_9668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5181 ( .C ( clk ), .D ( n2109 ), .Q ( new_AGEMA_signal_9670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5183 ( .C ( clk ), .D ( new_AGEMA_signal_2702 ), .Q ( new_AGEMA_signal_9672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5185 ( .C ( clk ), .D ( new_AGEMA_signal_2703 ), .Q ( new_AGEMA_signal_9674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5201 ( .C ( clk ), .D ( new_AGEMA_signal_9689 ), .Q ( new_AGEMA_signal_9690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5217 ( .C ( clk ), .D ( new_AGEMA_signal_9705 ), .Q ( new_AGEMA_signal_9706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5233 ( .C ( clk ), .D ( new_AGEMA_signal_9721 ), .Q ( new_AGEMA_signal_9722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5237 ( .C ( clk ), .D ( new_AGEMA_signal_9725 ), .Q ( new_AGEMA_signal_9726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5241 ( .C ( clk ), .D ( new_AGEMA_signal_9729 ), .Q ( new_AGEMA_signal_9730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5245 ( .C ( clk ), .D ( new_AGEMA_signal_9733 ), .Q ( new_AGEMA_signal_9734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5247 ( .C ( clk ), .D ( n2310 ), .Q ( new_AGEMA_signal_9736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5249 ( .C ( clk ), .D ( new_AGEMA_signal_2712 ), .Q ( new_AGEMA_signal_9738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5251 ( .C ( clk ), .D ( new_AGEMA_signal_2713 ), .Q ( new_AGEMA_signal_9740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5267 ( .C ( clk ), .D ( new_AGEMA_signal_9755 ), .Q ( new_AGEMA_signal_9756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5283 ( .C ( clk ), .D ( new_AGEMA_signal_9771 ), .Q ( new_AGEMA_signal_9772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5299 ( .C ( clk ), .D ( new_AGEMA_signal_9787 ), .Q ( new_AGEMA_signal_9788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5309 ( .C ( clk ), .D ( new_AGEMA_signal_9797 ), .Q ( new_AGEMA_signal_9798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5319 ( .C ( clk ), .D ( new_AGEMA_signal_9807 ), .Q ( new_AGEMA_signal_9808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5329 ( .C ( clk ), .D ( new_AGEMA_signal_9817 ), .Q ( new_AGEMA_signal_9818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5333 ( .C ( clk ), .D ( new_AGEMA_signal_9821 ), .Q ( new_AGEMA_signal_9822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5337 ( .C ( clk ), .D ( new_AGEMA_signal_9825 ), .Q ( new_AGEMA_signal_9826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5341 ( .C ( clk ), .D ( new_AGEMA_signal_9829 ), .Q ( new_AGEMA_signal_9830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5349 ( .C ( clk ), .D ( new_AGEMA_signal_9837 ), .Q ( new_AGEMA_signal_9838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5357 ( .C ( clk ), .D ( new_AGEMA_signal_9845 ), .Q ( new_AGEMA_signal_9846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5365 ( .C ( clk ), .D ( new_AGEMA_signal_9853 ), .Q ( new_AGEMA_signal_9854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5369 ( .C ( clk ), .D ( new_AGEMA_signal_9857 ), .Q ( new_AGEMA_signal_9858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5375 ( .C ( clk ), .D ( new_AGEMA_signal_9863 ), .Q ( new_AGEMA_signal_9864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5381 ( .C ( clk ), .D ( new_AGEMA_signal_9869 ), .Q ( new_AGEMA_signal_9870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5387 ( .C ( clk ), .D ( new_AGEMA_signal_9875 ), .Q ( new_AGEMA_signal_9876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5393 ( .C ( clk ), .D ( new_AGEMA_signal_9881 ), .Q ( new_AGEMA_signal_9882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5399 ( .C ( clk ), .D ( new_AGEMA_signal_9887 ), .Q ( new_AGEMA_signal_9888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5415 ( .C ( clk ), .D ( new_AGEMA_signal_9903 ), .Q ( new_AGEMA_signal_9904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5431 ( .C ( clk ), .D ( new_AGEMA_signal_9919 ), .Q ( new_AGEMA_signal_9920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5447 ( .C ( clk ), .D ( new_AGEMA_signal_9935 ), .Q ( new_AGEMA_signal_9936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5457 ( .C ( clk ), .D ( new_AGEMA_signal_9945 ), .Q ( new_AGEMA_signal_9946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5467 ( .C ( clk ), .D ( new_AGEMA_signal_9955 ), .Q ( new_AGEMA_signal_9956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5477 ( .C ( clk ), .D ( new_AGEMA_signal_9965 ), .Q ( new_AGEMA_signal_9966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5495 ( .C ( clk ), .D ( new_AGEMA_signal_9983 ), .Q ( new_AGEMA_signal_9984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5513 ( .C ( clk ), .D ( new_AGEMA_signal_10001 ), .Q ( new_AGEMA_signal_10002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5531 ( .C ( clk ), .D ( new_AGEMA_signal_10019 ), .Q ( new_AGEMA_signal_10020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5535 ( .C ( clk ), .D ( n2530 ), .Q ( new_AGEMA_signal_10024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5539 ( .C ( clk ), .D ( new_AGEMA_signal_2720 ), .Q ( new_AGEMA_signal_10028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5543 ( .C ( clk ), .D ( new_AGEMA_signal_2721 ), .Q ( new_AGEMA_signal_10032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5551 ( .C ( clk ), .D ( new_AGEMA_signal_10039 ), .Q ( new_AGEMA_signal_10040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5559 ( .C ( clk ), .D ( new_AGEMA_signal_10047 ), .Q ( new_AGEMA_signal_10048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5567 ( .C ( clk ), .D ( new_AGEMA_signal_10055 ), .Q ( new_AGEMA_signal_10056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5571 ( .C ( clk ), .D ( n2832 ), .Q ( new_AGEMA_signal_10060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5575 ( .C ( clk ), .D ( new_AGEMA_signal_2726 ), .Q ( new_AGEMA_signal_10064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5579 ( .C ( clk ), .D ( new_AGEMA_signal_2727 ), .Q ( new_AGEMA_signal_10068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5585 ( .C ( clk ), .D ( new_AGEMA_signal_10073 ), .Q ( new_AGEMA_signal_10074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5593 ( .C ( clk ), .D ( new_AGEMA_signal_10081 ), .Q ( new_AGEMA_signal_10082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5601 ( .C ( clk ), .D ( new_AGEMA_signal_10089 ), .Q ( new_AGEMA_signal_10090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5607 ( .C ( clk ), .D ( n2113 ), .Q ( new_AGEMA_signal_10096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5613 ( .C ( clk ), .D ( new_AGEMA_signal_2660 ), .Q ( new_AGEMA_signal_10102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5619 ( .C ( clk ), .D ( new_AGEMA_signal_2661 ), .Q ( new_AGEMA_signal_10108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5645 ( .C ( clk ), .D ( new_AGEMA_signal_10133 ), .Q ( new_AGEMA_signal_10134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5665 ( .C ( clk ), .D ( new_AGEMA_signal_10153 ), .Q ( new_AGEMA_signal_10154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5685 ( .C ( clk ), .D ( new_AGEMA_signal_10173 ), .Q ( new_AGEMA_signal_10174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5691 ( .C ( clk ), .D ( n2212 ), .Q ( new_AGEMA_signal_10180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5699 ( .C ( clk ), .D ( new_AGEMA_signal_2706 ), .Q ( new_AGEMA_signal_10188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5707 ( .C ( clk ), .D ( new_AGEMA_signal_2707 ), .Q ( new_AGEMA_signal_10196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5719 ( .C ( clk ), .D ( new_AGEMA_signal_10207 ), .Q ( new_AGEMA_signal_10208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5731 ( .C ( clk ), .D ( new_AGEMA_signal_10219 ), .Q ( new_AGEMA_signal_10220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5743 ( .C ( clk ), .D ( new_AGEMA_signal_10231 ), .Q ( new_AGEMA_signal_10232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5755 ( .C ( clk ), .D ( new_AGEMA_signal_10243 ), .Q ( new_AGEMA_signal_10244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5769 ( .C ( clk ), .D ( new_AGEMA_signal_10257 ), .Q ( new_AGEMA_signal_10258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5783 ( .C ( clk ), .D ( new_AGEMA_signal_10271 ), .Q ( new_AGEMA_signal_10272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5795 ( .C ( clk ), .D ( new_AGEMA_signal_10283 ), .Q ( new_AGEMA_signal_10284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5809 ( .C ( clk ), .D ( new_AGEMA_signal_10297 ), .Q ( new_AGEMA_signal_10298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5823 ( .C ( clk ), .D ( new_AGEMA_signal_10311 ), .Q ( new_AGEMA_signal_10312 ) ) ;

    /* cells in depth 22 */
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2129 ( .a ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, n2000}), .b ({new_AGEMA_signal_9465, new_AGEMA_signal_9457, new_AGEMA_signal_9449}), .clk ( clk ), .r ({Fresh[2504], Fresh[2503], Fresh[2502]}), .c ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, n2001}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2267 ( .a ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, n2107}), .b ({new_AGEMA_signal_9501, new_AGEMA_signal_9489, new_AGEMA_signal_9477}), .clk ( clk ), .r ({Fresh[2507], Fresh[2506], Fresh[2505]}), .c ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, n2108}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2317 ( .a ({new_AGEMA_signal_9543, new_AGEMA_signal_9529, new_AGEMA_signal_9515}), .b ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, n2149}), .clk ( clk ), .r ({Fresh[2510], Fresh[2509], Fresh[2508]}), .c ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, n2153}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2374 ( .a ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, n2206}), .b ({new_AGEMA_signal_9567, new_AGEMA_signal_9559, new_AGEMA_signal_9551}), .clk ( clk ), .r ({Fresh[2513], Fresh[2512], Fresh[2511]}), .c ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, n2207}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2477 ( .a ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, n2308}), .b ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, n2307}), .clk ( clk ), .r ({Fresh[2516], Fresh[2515], Fresh[2514]}), .c ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, n2309}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2535 ( .a ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, n2370}), .b ({new_AGEMA_signal_9609, new_AGEMA_signal_9595, new_AGEMA_signal_9581}), .clk ( clk ), .r ({Fresh[2519], Fresh[2518], Fresh[2517]}), .c ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, n2373}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2661 ( .a ({new_AGEMA_signal_9633, new_AGEMA_signal_9625, new_AGEMA_signal_9617}), .b ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, n2515}), .clk ( clk ), .r ({Fresh[2522], Fresh[2521], Fresh[2520]}), .c ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, n2528}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2750 ( .a ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, n2639}), .b ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, n2638}), .clk ( clk ), .r ({Fresh[2525], Fresh[2524], Fresh[2523]}), .c ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, n2669}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2843 ( .a ({new_AGEMA_signal_9657, new_AGEMA_signal_9649, new_AGEMA_signal_9641}), .b ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, n2807}), .clk ( clk ), .r ({Fresh[2528], Fresh[2527], Fresh[2526]}), .c ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, n2830}) ) ;
    buf_clk new_AGEMA_reg_buffer_5172 ( .C ( clk ), .D ( new_AGEMA_signal_9660 ), .Q ( new_AGEMA_signal_9661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5176 ( .C ( clk ), .D ( new_AGEMA_signal_9664 ), .Q ( new_AGEMA_signal_9665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5180 ( .C ( clk ), .D ( new_AGEMA_signal_9668 ), .Q ( new_AGEMA_signal_9669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5182 ( .C ( clk ), .D ( new_AGEMA_signal_9670 ), .Q ( new_AGEMA_signal_9671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5184 ( .C ( clk ), .D ( new_AGEMA_signal_9672 ), .Q ( new_AGEMA_signal_9673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5186 ( .C ( clk ), .D ( new_AGEMA_signal_9674 ), .Q ( new_AGEMA_signal_9675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5202 ( .C ( clk ), .D ( new_AGEMA_signal_9690 ), .Q ( new_AGEMA_signal_9691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5218 ( .C ( clk ), .D ( new_AGEMA_signal_9706 ), .Q ( new_AGEMA_signal_9707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5234 ( .C ( clk ), .D ( new_AGEMA_signal_9722 ), .Q ( new_AGEMA_signal_9723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5238 ( .C ( clk ), .D ( new_AGEMA_signal_9726 ), .Q ( new_AGEMA_signal_9727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5242 ( .C ( clk ), .D ( new_AGEMA_signal_9730 ), .Q ( new_AGEMA_signal_9731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5246 ( .C ( clk ), .D ( new_AGEMA_signal_9734 ), .Q ( new_AGEMA_signal_9735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5248 ( .C ( clk ), .D ( new_AGEMA_signal_9736 ), .Q ( new_AGEMA_signal_9737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5250 ( .C ( clk ), .D ( new_AGEMA_signal_9738 ), .Q ( new_AGEMA_signal_9739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5252 ( .C ( clk ), .D ( new_AGEMA_signal_9740 ), .Q ( new_AGEMA_signal_9741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5268 ( .C ( clk ), .D ( new_AGEMA_signal_9756 ), .Q ( new_AGEMA_signal_9757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5284 ( .C ( clk ), .D ( new_AGEMA_signal_9772 ), .Q ( new_AGEMA_signal_9773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5300 ( .C ( clk ), .D ( new_AGEMA_signal_9788 ), .Q ( new_AGEMA_signal_9789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5310 ( .C ( clk ), .D ( new_AGEMA_signal_9798 ), .Q ( new_AGEMA_signal_9799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5320 ( .C ( clk ), .D ( new_AGEMA_signal_9808 ), .Q ( new_AGEMA_signal_9809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5330 ( .C ( clk ), .D ( new_AGEMA_signal_9818 ), .Q ( new_AGEMA_signal_9819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5334 ( .C ( clk ), .D ( new_AGEMA_signal_9822 ), .Q ( new_AGEMA_signal_9823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5338 ( .C ( clk ), .D ( new_AGEMA_signal_9826 ), .Q ( new_AGEMA_signal_9827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5342 ( .C ( clk ), .D ( new_AGEMA_signal_9830 ), .Q ( new_AGEMA_signal_9831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5350 ( .C ( clk ), .D ( new_AGEMA_signal_9838 ), .Q ( new_AGEMA_signal_9839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5358 ( .C ( clk ), .D ( new_AGEMA_signal_9846 ), .Q ( new_AGEMA_signal_9847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5366 ( .C ( clk ), .D ( new_AGEMA_signal_9854 ), .Q ( new_AGEMA_signal_9855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5370 ( .C ( clk ), .D ( new_AGEMA_signal_9858 ), .Q ( new_AGEMA_signal_9859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5376 ( .C ( clk ), .D ( new_AGEMA_signal_9864 ), .Q ( new_AGEMA_signal_9865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5382 ( .C ( clk ), .D ( new_AGEMA_signal_9870 ), .Q ( new_AGEMA_signal_9871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5388 ( .C ( clk ), .D ( new_AGEMA_signal_9876 ), .Q ( new_AGEMA_signal_9877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5394 ( .C ( clk ), .D ( new_AGEMA_signal_9882 ), .Q ( new_AGEMA_signal_9883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5400 ( .C ( clk ), .D ( new_AGEMA_signal_9888 ), .Q ( new_AGEMA_signal_9889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5416 ( .C ( clk ), .D ( new_AGEMA_signal_9904 ), .Q ( new_AGEMA_signal_9905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5432 ( .C ( clk ), .D ( new_AGEMA_signal_9920 ), .Q ( new_AGEMA_signal_9921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5448 ( .C ( clk ), .D ( new_AGEMA_signal_9936 ), .Q ( new_AGEMA_signal_9937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5458 ( .C ( clk ), .D ( new_AGEMA_signal_9946 ), .Q ( new_AGEMA_signal_9947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5468 ( .C ( clk ), .D ( new_AGEMA_signal_9956 ), .Q ( new_AGEMA_signal_9957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5478 ( .C ( clk ), .D ( new_AGEMA_signal_9966 ), .Q ( new_AGEMA_signal_9967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5496 ( .C ( clk ), .D ( new_AGEMA_signal_9984 ), .Q ( new_AGEMA_signal_9985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5514 ( .C ( clk ), .D ( new_AGEMA_signal_10002 ), .Q ( new_AGEMA_signal_10003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5532 ( .C ( clk ), .D ( new_AGEMA_signal_10020 ), .Q ( new_AGEMA_signal_10021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5536 ( .C ( clk ), .D ( new_AGEMA_signal_10024 ), .Q ( new_AGEMA_signal_10025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5540 ( .C ( clk ), .D ( new_AGEMA_signal_10028 ), .Q ( new_AGEMA_signal_10029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5544 ( .C ( clk ), .D ( new_AGEMA_signal_10032 ), .Q ( new_AGEMA_signal_10033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5552 ( .C ( clk ), .D ( new_AGEMA_signal_10040 ), .Q ( new_AGEMA_signal_10041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5560 ( .C ( clk ), .D ( new_AGEMA_signal_10048 ), .Q ( new_AGEMA_signal_10049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5568 ( .C ( clk ), .D ( new_AGEMA_signal_10056 ), .Q ( new_AGEMA_signal_10057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5572 ( .C ( clk ), .D ( new_AGEMA_signal_10060 ), .Q ( new_AGEMA_signal_10061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5576 ( .C ( clk ), .D ( new_AGEMA_signal_10064 ), .Q ( new_AGEMA_signal_10065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5580 ( .C ( clk ), .D ( new_AGEMA_signal_10068 ), .Q ( new_AGEMA_signal_10069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5586 ( .C ( clk ), .D ( new_AGEMA_signal_10074 ), .Q ( new_AGEMA_signal_10075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5594 ( .C ( clk ), .D ( new_AGEMA_signal_10082 ), .Q ( new_AGEMA_signal_10083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5602 ( .C ( clk ), .D ( new_AGEMA_signal_10090 ), .Q ( new_AGEMA_signal_10091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5608 ( .C ( clk ), .D ( new_AGEMA_signal_10096 ), .Q ( new_AGEMA_signal_10097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5614 ( .C ( clk ), .D ( new_AGEMA_signal_10102 ), .Q ( new_AGEMA_signal_10103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5620 ( .C ( clk ), .D ( new_AGEMA_signal_10108 ), .Q ( new_AGEMA_signal_10109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5646 ( .C ( clk ), .D ( new_AGEMA_signal_10134 ), .Q ( new_AGEMA_signal_10135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5666 ( .C ( clk ), .D ( new_AGEMA_signal_10154 ), .Q ( new_AGEMA_signal_10155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5686 ( .C ( clk ), .D ( new_AGEMA_signal_10174 ), .Q ( new_AGEMA_signal_10175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5692 ( .C ( clk ), .D ( new_AGEMA_signal_10180 ), .Q ( new_AGEMA_signal_10181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5700 ( .C ( clk ), .D ( new_AGEMA_signal_10188 ), .Q ( new_AGEMA_signal_10189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5708 ( .C ( clk ), .D ( new_AGEMA_signal_10196 ), .Q ( new_AGEMA_signal_10197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5720 ( .C ( clk ), .D ( new_AGEMA_signal_10208 ), .Q ( new_AGEMA_signal_10209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5732 ( .C ( clk ), .D ( new_AGEMA_signal_10220 ), .Q ( new_AGEMA_signal_10221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5744 ( .C ( clk ), .D ( new_AGEMA_signal_10232 ), .Q ( new_AGEMA_signal_10233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5756 ( .C ( clk ), .D ( new_AGEMA_signal_10244 ), .Q ( new_AGEMA_signal_10245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5770 ( .C ( clk ), .D ( new_AGEMA_signal_10258 ), .Q ( new_AGEMA_signal_10259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5784 ( .C ( clk ), .D ( new_AGEMA_signal_10272 ), .Q ( new_AGEMA_signal_10273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5796 ( .C ( clk ), .D ( new_AGEMA_signal_10284 ), .Q ( new_AGEMA_signal_10285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5810 ( .C ( clk ), .D ( new_AGEMA_signal_10298 ), .Q ( new_AGEMA_signal_10299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5824 ( .C ( clk ), .D ( new_AGEMA_signal_10312 ), .Q ( new_AGEMA_signal_10313 ) ) ;

    /* cells in depth 23 */
    buf_clk new_AGEMA_reg_buffer_5371 ( .C ( clk ), .D ( new_AGEMA_signal_9859 ), .Q ( new_AGEMA_signal_9860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5377 ( .C ( clk ), .D ( new_AGEMA_signal_9865 ), .Q ( new_AGEMA_signal_9866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5383 ( .C ( clk ), .D ( new_AGEMA_signal_9871 ), .Q ( new_AGEMA_signal_9872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5389 ( .C ( clk ), .D ( new_AGEMA_signal_9877 ), .Q ( new_AGEMA_signal_9878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5395 ( .C ( clk ), .D ( new_AGEMA_signal_9883 ), .Q ( new_AGEMA_signal_9884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5401 ( .C ( clk ), .D ( new_AGEMA_signal_9889 ), .Q ( new_AGEMA_signal_9890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5417 ( .C ( clk ), .D ( new_AGEMA_signal_9905 ), .Q ( new_AGEMA_signal_9906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5433 ( .C ( clk ), .D ( new_AGEMA_signal_9921 ), .Q ( new_AGEMA_signal_9922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5449 ( .C ( clk ), .D ( new_AGEMA_signal_9937 ), .Q ( new_AGEMA_signal_9938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5459 ( .C ( clk ), .D ( new_AGEMA_signal_9947 ), .Q ( new_AGEMA_signal_9948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5469 ( .C ( clk ), .D ( new_AGEMA_signal_9957 ), .Q ( new_AGEMA_signal_9958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5479 ( .C ( clk ), .D ( new_AGEMA_signal_9967 ), .Q ( new_AGEMA_signal_9968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5497 ( .C ( clk ), .D ( new_AGEMA_signal_9985 ), .Q ( new_AGEMA_signal_9986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5515 ( .C ( clk ), .D ( new_AGEMA_signal_10003 ), .Q ( new_AGEMA_signal_10004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5533 ( .C ( clk ), .D ( new_AGEMA_signal_10021 ), .Q ( new_AGEMA_signal_10022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5537 ( .C ( clk ), .D ( new_AGEMA_signal_10025 ), .Q ( new_AGEMA_signal_10026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5541 ( .C ( clk ), .D ( new_AGEMA_signal_10029 ), .Q ( new_AGEMA_signal_10030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5545 ( .C ( clk ), .D ( new_AGEMA_signal_10033 ), .Q ( new_AGEMA_signal_10034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5553 ( .C ( clk ), .D ( new_AGEMA_signal_10041 ), .Q ( new_AGEMA_signal_10042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5561 ( .C ( clk ), .D ( new_AGEMA_signal_10049 ), .Q ( new_AGEMA_signal_10050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5569 ( .C ( clk ), .D ( new_AGEMA_signal_10057 ), .Q ( new_AGEMA_signal_10058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5573 ( .C ( clk ), .D ( new_AGEMA_signal_10061 ), .Q ( new_AGEMA_signal_10062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5577 ( .C ( clk ), .D ( new_AGEMA_signal_10065 ), .Q ( new_AGEMA_signal_10066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5581 ( .C ( clk ), .D ( new_AGEMA_signal_10069 ), .Q ( new_AGEMA_signal_10070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5587 ( .C ( clk ), .D ( new_AGEMA_signal_10075 ), .Q ( new_AGEMA_signal_10076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5595 ( .C ( clk ), .D ( new_AGEMA_signal_10083 ), .Q ( new_AGEMA_signal_10084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5603 ( .C ( clk ), .D ( new_AGEMA_signal_10091 ), .Q ( new_AGEMA_signal_10092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5609 ( .C ( clk ), .D ( new_AGEMA_signal_10097 ), .Q ( new_AGEMA_signal_10098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5615 ( .C ( clk ), .D ( new_AGEMA_signal_10103 ), .Q ( new_AGEMA_signal_10104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5621 ( .C ( clk ), .D ( new_AGEMA_signal_10109 ), .Q ( new_AGEMA_signal_10110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5647 ( .C ( clk ), .D ( new_AGEMA_signal_10135 ), .Q ( new_AGEMA_signal_10136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5667 ( .C ( clk ), .D ( new_AGEMA_signal_10155 ), .Q ( new_AGEMA_signal_10156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5687 ( .C ( clk ), .D ( new_AGEMA_signal_10175 ), .Q ( new_AGEMA_signal_10176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5693 ( .C ( clk ), .D ( new_AGEMA_signal_10181 ), .Q ( new_AGEMA_signal_10182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5701 ( .C ( clk ), .D ( new_AGEMA_signal_10189 ), .Q ( new_AGEMA_signal_10190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5709 ( .C ( clk ), .D ( new_AGEMA_signal_10197 ), .Q ( new_AGEMA_signal_10198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5721 ( .C ( clk ), .D ( new_AGEMA_signal_10209 ), .Q ( new_AGEMA_signal_10210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5733 ( .C ( clk ), .D ( new_AGEMA_signal_10221 ), .Q ( new_AGEMA_signal_10222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5745 ( .C ( clk ), .D ( new_AGEMA_signal_10233 ), .Q ( new_AGEMA_signal_10234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5757 ( .C ( clk ), .D ( new_AGEMA_signal_10245 ), .Q ( new_AGEMA_signal_10246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5771 ( .C ( clk ), .D ( new_AGEMA_signal_10259 ), .Q ( new_AGEMA_signal_10260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5785 ( .C ( clk ), .D ( new_AGEMA_signal_10273 ), .Q ( new_AGEMA_signal_10274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5797 ( .C ( clk ), .D ( new_AGEMA_signal_10285 ), .Q ( new_AGEMA_signal_10286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5811 ( .C ( clk ), .D ( new_AGEMA_signal_10299 ), .Q ( new_AGEMA_signal_10300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5825 ( .C ( clk ), .D ( new_AGEMA_signal_10313 ), .Q ( new_AGEMA_signal_10314 ) ) ;

    /* cells in depth 24 */
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2130 ( .a ({new_AGEMA_signal_9669, new_AGEMA_signal_9665, new_AGEMA_signal_9661}), .b ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, n2001}), .clk ( clk ), .r ({Fresh[2531], Fresh[2530], Fresh[2529]}), .c ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, n2017}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2268 ( .a ({new_AGEMA_signal_9675, new_AGEMA_signal_9673, new_AGEMA_signal_9671}), .b ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, n2108}), .clk ( clk ), .r ({Fresh[2534], Fresh[2533], Fresh[2532]}), .c ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, n2110}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2319 ( .a ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, n2153}), .b ({new_AGEMA_signal_9723, new_AGEMA_signal_9707, new_AGEMA_signal_9691}), .clk ( clk ), .r ({Fresh[2537], Fresh[2536], Fresh[2535]}), .c ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, n2154}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2375 ( .a ({new_AGEMA_signal_9735, new_AGEMA_signal_9731, new_AGEMA_signal_9727}), .b ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, n2207}), .clk ( clk ), .r ({Fresh[2540], Fresh[2539], Fresh[2538]}), .c ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, n2209}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2478 ( .a ({new_AGEMA_signal_9741, new_AGEMA_signal_9739, new_AGEMA_signal_9737}), .b ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, n2309}), .clk ( clk ), .r ({Fresh[2543], Fresh[2542], Fresh[2541]}), .c ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, n2311}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2537 ( .a ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, n2373}), .b ({new_AGEMA_signal_9789, new_AGEMA_signal_9773, new_AGEMA_signal_9757}), .clk ( clk ), .r ({Fresh[2546], Fresh[2545], Fresh[2544]}), .c ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, n2374}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2672 ( .a ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, n2528}), .b ({new_AGEMA_signal_9819, new_AGEMA_signal_9809, new_AGEMA_signal_9799}), .clk ( clk ), .r ({Fresh[2549], Fresh[2548], Fresh[2547]}), .c ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, n2529}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2768 ( .a ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, n2669}), .b ({new_AGEMA_signal_9831, new_AGEMA_signal_9827, new_AGEMA_signal_9823}), .clk ( clk ), .r ({Fresh[2552], Fresh[2551], Fresh[2550]}), .c ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, n2670}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2854 ( .a ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, n2830}), .b ({new_AGEMA_signal_9855, new_AGEMA_signal_9847, new_AGEMA_signal_9839}), .clk ( clk ), .r ({Fresh[2555], Fresh[2554], Fresh[2553]}), .c ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, n2831}) ) ;
    buf_clk new_AGEMA_reg_buffer_5372 ( .C ( clk ), .D ( new_AGEMA_signal_9860 ), .Q ( new_AGEMA_signal_9861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5378 ( .C ( clk ), .D ( new_AGEMA_signal_9866 ), .Q ( new_AGEMA_signal_9867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5384 ( .C ( clk ), .D ( new_AGEMA_signal_9872 ), .Q ( new_AGEMA_signal_9873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5390 ( .C ( clk ), .D ( new_AGEMA_signal_9878 ), .Q ( new_AGEMA_signal_9879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5396 ( .C ( clk ), .D ( new_AGEMA_signal_9884 ), .Q ( new_AGEMA_signal_9885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5402 ( .C ( clk ), .D ( new_AGEMA_signal_9890 ), .Q ( new_AGEMA_signal_9891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5418 ( .C ( clk ), .D ( new_AGEMA_signal_9906 ), .Q ( new_AGEMA_signal_9907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5434 ( .C ( clk ), .D ( new_AGEMA_signal_9922 ), .Q ( new_AGEMA_signal_9923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5450 ( .C ( clk ), .D ( new_AGEMA_signal_9938 ), .Q ( new_AGEMA_signal_9939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5460 ( .C ( clk ), .D ( new_AGEMA_signal_9948 ), .Q ( new_AGEMA_signal_9949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5470 ( .C ( clk ), .D ( new_AGEMA_signal_9958 ), .Q ( new_AGEMA_signal_9959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5480 ( .C ( clk ), .D ( new_AGEMA_signal_9968 ), .Q ( new_AGEMA_signal_9969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5498 ( .C ( clk ), .D ( new_AGEMA_signal_9986 ), .Q ( new_AGEMA_signal_9987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5516 ( .C ( clk ), .D ( new_AGEMA_signal_10004 ), .Q ( new_AGEMA_signal_10005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5534 ( .C ( clk ), .D ( new_AGEMA_signal_10022 ), .Q ( new_AGEMA_signal_10023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5538 ( .C ( clk ), .D ( new_AGEMA_signal_10026 ), .Q ( new_AGEMA_signal_10027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5542 ( .C ( clk ), .D ( new_AGEMA_signal_10030 ), .Q ( new_AGEMA_signal_10031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5546 ( .C ( clk ), .D ( new_AGEMA_signal_10034 ), .Q ( new_AGEMA_signal_10035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5554 ( .C ( clk ), .D ( new_AGEMA_signal_10042 ), .Q ( new_AGEMA_signal_10043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5562 ( .C ( clk ), .D ( new_AGEMA_signal_10050 ), .Q ( new_AGEMA_signal_10051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5570 ( .C ( clk ), .D ( new_AGEMA_signal_10058 ), .Q ( new_AGEMA_signal_10059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5574 ( .C ( clk ), .D ( new_AGEMA_signal_10062 ), .Q ( new_AGEMA_signal_10063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5578 ( .C ( clk ), .D ( new_AGEMA_signal_10066 ), .Q ( new_AGEMA_signal_10067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5582 ( .C ( clk ), .D ( new_AGEMA_signal_10070 ), .Q ( new_AGEMA_signal_10071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5588 ( .C ( clk ), .D ( new_AGEMA_signal_10076 ), .Q ( new_AGEMA_signal_10077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5596 ( .C ( clk ), .D ( new_AGEMA_signal_10084 ), .Q ( new_AGEMA_signal_10085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5604 ( .C ( clk ), .D ( new_AGEMA_signal_10092 ), .Q ( new_AGEMA_signal_10093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5610 ( .C ( clk ), .D ( new_AGEMA_signal_10098 ), .Q ( new_AGEMA_signal_10099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5616 ( .C ( clk ), .D ( new_AGEMA_signal_10104 ), .Q ( new_AGEMA_signal_10105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5622 ( .C ( clk ), .D ( new_AGEMA_signal_10110 ), .Q ( new_AGEMA_signal_10111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5648 ( .C ( clk ), .D ( new_AGEMA_signal_10136 ), .Q ( new_AGEMA_signal_10137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5668 ( .C ( clk ), .D ( new_AGEMA_signal_10156 ), .Q ( new_AGEMA_signal_10157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5688 ( .C ( clk ), .D ( new_AGEMA_signal_10176 ), .Q ( new_AGEMA_signal_10177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5694 ( .C ( clk ), .D ( new_AGEMA_signal_10182 ), .Q ( new_AGEMA_signal_10183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5702 ( .C ( clk ), .D ( new_AGEMA_signal_10190 ), .Q ( new_AGEMA_signal_10191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5710 ( .C ( clk ), .D ( new_AGEMA_signal_10198 ), .Q ( new_AGEMA_signal_10199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5722 ( .C ( clk ), .D ( new_AGEMA_signal_10210 ), .Q ( new_AGEMA_signal_10211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5734 ( .C ( clk ), .D ( new_AGEMA_signal_10222 ), .Q ( new_AGEMA_signal_10223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5746 ( .C ( clk ), .D ( new_AGEMA_signal_10234 ), .Q ( new_AGEMA_signal_10235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5758 ( .C ( clk ), .D ( new_AGEMA_signal_10246 ), .Q ( new_AGEMA_signal_10247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5772 ( .C ( clk ), .D ( new_AGEMA_signal_10260 ), .Q ( new_AGEMA_signal_10261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5786 ( .C ( clk ), .D ( new_AGEMA_signal_10274 ), .Q ( new_AGEMA_signal_10275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5798 ( .C ( clk ), .D ( new_AGEMA_signal_10286 ), .Q ( new_AGEMA_signal_10287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5812 ( .C ( clk ), .D ( new_AGEMA_signal_10300 ), .Q ( new_AGEMA_signal_10301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5826 ( .C ( clk ), .D ( new_AGEMA_signal_10314 ), .Q ( new_AGEMA_signal_10315 ) ) ;

    /* cells in depth 25 */
    buf_clk new_AGEMA_reg_buffer_5589 ( .C ( clk ), .D ( new_AGEMA_signal_10077 ), .Q ( new_AGEMA_signal_10078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5597 ( .C ( clk ), .D ( new_AGEMA_signal_10085 ), .Q ( new_AGEMA_signal_10086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5605 ( .C ( clk ), .D ( new_AGEMA_signal_10093 ), .Q ( new_AGEMA_signal_10094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5611 ( .C ( clk ), .D ( new_AGEMA_signal_10099 ), .Q ( new_AGEMA_signal_10100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5617 ( .C ( clk ), .D ( new_AGEMA_signal_10105 ), .Q ( new_AGEMA_signal_10106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5623 ( .C ( clk ), .D ( new_AGEMA_signal_10111 ), .Q ( new_AGEMA_signal_10112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5625 ( .C ( clk ), .D ( n2209 ), .Q ( new_AGEMA_signal_10114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5627 ( .C ( clk ), .D ( new_AGEMA_signal_2754 ), .Q ( new_AGEMA_signal_10116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5629 ( .C ( clk ), .D ( new_AGEMA_signal_2755 ), .Q ( new_AGEMA_signal_10118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5649 ( .C ( clk ), .D ( new_AGEMA_signal_10137 ), .Q ( new_AGEMA_signal_10138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5669 ( .C ( clk ), .D ( new_AGEMA_signal_10157 ), .Q ( new_AGEMA_signal_10158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5689 ( .C ( clk ), .D ( new_AGEMA_signal_10177 ), .Q ( new_AGEMA_signal_10178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5695 ( .C ( clk ), .D ( new_AGEMA_signal_10183 ), .Q ( new_AGEMA_signal_10184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5703 ( .C ( clk ), .D ( new_AGEMA_signal_10191 ), .Q ( new_AGEMA_signal_10192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5711 ( .C ( clk ), .D ( new_AGEMA_signal_10199 ), .Q ( new_AGEMA_signal_10200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5723 ( .C ( clk ), .D ( new_AGEMA_signal_10211 ), .Q ( new_AGEMA_signal_10212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5735 ( .C ( clk ), .D ( new_AGEMA_signal_10223 ), .Q ( new_AGEMA_signal_10224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5747 ( .C ( clk ), .D ( new_AGEMA_signal_10235 ), .Q ( new_AGEMA_signal_10236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5759 ( .C ( clk ), .D ( new_AGEMA_signal_10247 ), .Q ( new_AGEMA_signal_10248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5773 ( .C ( clk ), .D ( new_AGEMA_signal_10261 ), .Q ( new_AGEMA_signal_10262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5787 ( .C ( clk ), .D ( new_AGEMA_signal_10275 ), .Q ( new_AGEMA_signal_10276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5799 ( .C ( clk ), .D ( new_AGEMA_signal_10287 ), .Q ( new_AGEMA_signal_10288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5813 ( .C ( clk ), .D ( new_AGEMA_signal_10301 ), .Q ( new_AGEMA_signal_10302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5827 ( .C ( clk ), .D ( new_AGEMA_signal_10315 ), .Q ( new_AGEMA_signal_10316 ) ) ;

    /* cells in depth 26 */
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2155 ( .a ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, n2017}), .b ({new_AGEMA_signal_9873, new_AGEMA_signal_9867, new_AGEMA_signal_9861}), .clk ( clk ), .r ({Fresh[2558], Fresh[2557], Fresh[2556]}), .c ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, n2018}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2269 ( .a ({new_AGEMA_signal_9891, new_AGEMA_signal_9885, new_AGEMA_signal_9879}), .b ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, n2110}), .clk ( clk ), .r ({Fresh[2561], Fresh[2560], Fresh[2559]}), .c ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, n2112}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2320 ( .a ({new_AGEMA_signal_9939, new_AGEMA_signal_9923, new_AGEMA_signal_9907}), .b ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, n2154}), .clk ( clk ), .r ({Fresh[2564], Fresh[2563], Fresh[2562]}), .c ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, n2210}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2479 ( .a ({new_AGEMA_signal_9969, new_AGEMA_signal_9959, new_AGEMA_signal_9949}), .b ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, n2311}), .clk ( clk ), .r ({Fresh[2567], Fresh[2566], Fresh[2565]}), .c ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, N470}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2538 ( .a ({new_AGEMA_signal_10023, new_AGEMA_signal_10005, new_AGEMA_signal_9987}), .b ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, n2374}), .clk ( clk ), .r ({Fresh[2570], Fresh[2569], Fresh[2568]}), .c ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, n2378}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2673 ( .a ({new_AGEMA_signal_10035, new_AGEMA_signal_10031, new_AGEMA_signal_10027}), .b ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, n2529}), .clk ( clk ), .r ({Fresh[2573], Fresh[2572], Fresh[2571]}), .c ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, N639}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2769 ( .a ({new_AGEMA_signal_10059, new_AGEMA_signal_10051, new_AGEMA_signal_10043}), .b ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, n2670}), .clk ( clk ), .r ({Fresh[2576], Fresh[2575], Fresh[2574]}), .c ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, N723}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2855 ( .a ({new_AGEMA_signal_10071, new_AGEMA_signal_10067, new_AGEMA_signal_10063}), .b ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, n2831}), .clk ( clk ), .r ({Fresh[2579], Fresh[2578], Fresh[2577]}), .c ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, N789}) ) ;
    buf_clk new_AGEMA_reg_buffer_5590 ( .C ( clk ), .D ( new_AGEMA_signal_10078 ), .Q ( new_AGEMA_signal_10079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5598 ( .C ( clk ), .D ( new_AGEMA_signal_10086 ), .Q ( new_AGEMA_signal_10087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5606 ( .C ( clk ), .D ( new_AGEMA_signal_10094 ), .Q ( new_AGEMA_signal_10095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5612 ( .C ( clk ), .D ( new_AGEMA_signal_10100 ), .Q ( new_AGEMA_signal_10101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5618 ( .C ( clk ), .D ( new_AGEMA_signal_10106 ), .Q ( new_AGEMA_signal_10107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5624 ( .C ( clk ), .D ( new_AGEMA_signal_10112 ), .Q ( new_AGEMA_signal_10113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5626 ( .C ( clk ), .D ( new_AGEMA_signal_10114 ), .Q ( new_AGEMA_signal_10115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5628 ( .C ( clk ), .D ( new_AGEMA_signal_10116 ), .Q ( new_AGEMA_signal_10117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5630 ( .C ( clk ), .D ( new_AGEMA_signal_10118 ), .Q ( new_AGEMA_signal_10119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5650 ( .C ( clk ), .D ( new_AGEMA_signal_10138 ), .Q ( new_AGEMA_signal_10139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5670 ( .C ( clk ), .D ( new_AGEMA_signal_10158 ), .Q ( new_AGEMA_signal_10159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5690 ( .C ( clk ), .D ( new_AGEMA_signal_10178 ), .Q ( new_AGEMA_signal_10179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5696 ( .C ( clk ), .D ( new_AGEMA_signal_10184 ), .Q ( new_AGEMA_signal_10185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5704 ( .C ( clk ), .D ( new_AGEMA_signal_10192 ), .Q ( new_AGEMA_signal_10193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5712 ( .C ( clk ), .D ( new_AGEMA_signal_10200 ), .Q ( new_AGEMA_signal_10201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5724 ( .C ( clk ), .D ( new_AGEMA_signal_10212 ), .Q ( new_AGEMA_signal_10213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5736 ( .C ( clk ), .D ( new_AGEMA_signal_10224 ), .Q ( new_AGEMA_signal_10225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5748 ( .C ( clk ), .D ( new_AGEMA_signal_10236 ), .Q ( new_AGEMA_signal_10237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5760 ( .C ( clk ), .D ( new_AGEMA_signal_10248 ), .Q ( new_AGEMA_signal_10249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5774 ( .C ( clk ), .D ( new_AGEMA_signal_10262 ), .Q ( new_AGEMA_signal_10263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5788 ( .C ( clk ), .D ( new_AGEMA_signal_10276 ), .Q ( new_AGEMA_signal_10277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5800 ( .C ( clk ), .D ( new_AGEMA_signal_10288 ), .Q ( new_AGEMA_signal_10289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5814 ( .C ( clk ), .D ( new_AGEMA_signal_10302 ), .Q ( new_AGEMA_signal_10303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5828 ( .C ( clk ), .D ( new_AGEMA_signal_10316 ), .Q ( new_AGEMA_signal_10317 ) ) ;

    /* cells in depth 27 */
    buf_clk new_AGEMA_reg_buffer_5697 ( .C ( clk ), .D ( new_AGEMA_signal_10185 ), .Q ( new_AGEMA_signal_10186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5705 ( .C ( clk ), .D ( new_AGEMA_signal_10193 ), .Q ( new_AGEMA_signal_10194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5713 ( .C ( clk ), .D ( new_AGEMA_signal_10201 ), .Q ( new_AGEMA_signal_10202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5725 ( .C ( clk ), .D ( new_AGEMA_signal_10213 ), .Q ( new_AGEMA_signal_10214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5737 ( .C ( clk ), .D ( new_AGEMA_signal_10225 ), .Q ( new_AGEMA_signal_10226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5749 ( .C ( clk ), .D ( new_AGEMA_signal_10237 ), .Q ( new_AGEMA_signal_10238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5761 ( .C ( clk ), .D ( new_AGEMA_signal_10249 ), .Q ( new_AGEMA_signal_10250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5775 ( .C ( clk ), .D ( new_AGEMA_signal_10263 ), .Q ( new_AGEMA_signal_10264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5789 ( .C ( clk ), .D ( new_AGEMA_signal_10277 ), .Q ( new_AGEMA_signal_10278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5801 ( .C ( clk ), .D ( new_AGEMA_signal_10289 ), .Q ( new_AGEMA_signal_10290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5815 ( .C ( clk ), .D ( new_AGEMA_signal_10303 ), .Q ( new_AGEMA_signal_10304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5829 ( .C ( clk ), .D ( new_AGEMA_signal_10317 ), .Q ( new_AGEMA_signal_10318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5883 ( .C ( clk ), .D ( N470 ), .Q ( new_AGEMA_signal_10372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5891 ( .C ( clk ), .D ( new_AGEMA_signal_2772 ), .Q ( new_AGEMA_signal_10380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5899 ( .C ( clk ), .D ( new_AGEMA_signal_2773 ), .Q ( new_AGEMA_signal_10388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5907 ( .C ( clk ), .D ( N639 ), .Q ( new_AGEMA_signal_10396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5915 ( .C ( clk ), .D ( new_AGEMA_signal_2776 ), .Q ( new_AGEMA_signal_10404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5923 ( .C ( clk ), .D ( new_AGEMA_signal_2777 ), .Q ( new_AGEMA_signal_10412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5931 ( .C ( clk ), .D ( N723 ), .Q ( new_AGEMA_signal_10420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5939 ( .C ( clk ), .D ( new_AGEMA_signal_2778 ), .Q ( new_AGEMA_signal_10428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5947 ( .C ( clk ), .D ( new_AGEMA_signal_2779 ), .Q ( new_AGEMA_signal_10436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5955 ( .C ( clk ), .D ( N789 ), .Q ( new_AGEMA_signal_10444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5963 ( .C ( clk ), .D ( new_AGEMA_signal_2764 ), .Q ( new_AGEMA_signal_10452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5971 ( .C ( clk ), .D ( new_AGEMA_signal_2765 ), .Q ( new_AGEMA_signal_10460 ) ) ;

    /* cells in depth 28 */
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2156 ( .a ({new_AGEMA_signal_10095, new_AGEMA_signal_10087, new_AGEMA_signal_10079}), .b ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, n2018}), .clk ( clk ), .r ({Fresh[2582], Fresh[2581], Fresh[2580]}), .c ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, N169}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2270 ( .a ({new_AGEMA_signal_10113, new_AGEMA_signal_10107, new_AGEMA_signal_10101}), .b ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, n2112}), .clk ( clk ), .r ({Fresh[2585], Fresh[2584], Fresh[2583]}), .c ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, N277}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2376 ( .a ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, n2210}), .b ({new_AGEMA_signal_10119, new_AGEMA_signal_10117, new_AGEMA_signal_10115}), .clk ( clk ), .r ({Fresh[2588], Fresh[2587], Fresh[2586]}), .c ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, n2211}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2540 ( .a ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, n2378}), .b ({new_AGEMA_signal_10179, new_AGEMA_signal_10159, new_AGEMA_signal_10139}), .clk ( clk ), .r ({Fresh[2591], Fresh[2590], Fresh[2589]}), .c ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, n2379}) ) ;
    buf_clk new_AGEMA_reg_buffer_5698 ( .C ( clk ), .D ( new_AGEMA_signal_10186 ), .Q ( new_AGEMA_signal_10187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5706 ( .C ( clk ), .D ( new_AGEMA_signal_10194 ), .Q ( new_AGEMA_signal_10195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5714 ( .C ( clk ), .D ( new_AGEMA_signal_10202 ), .Q ( new_AGEMA_signal_10203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5726 ( .C ( clk ), .D ( new_AGEMA_signal_10214 ), .Q ( new_AGEMA_signal_10215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5738 ( .C ( clk ), .D ( new_AGEMA_signal_10226 ), .Q ( new_AGEMA_signal_10227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5750 ( .C ( clk ), .D ( new_AGEMA_signal_10238 ), .Q ( new_AGEMA_signal_10239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5762 ( .C ( clk ), .D ( new_AGEMA_signal_10250 ), .Q ( new_AGEMA_signal_10251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5776 ( .C ( clk ), .D ( new_AGEMA_signal_10264 ), .Q ( new_AGEMA_signal_10265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5790 ( .C ( clk ), .D ( new_AGEMA_signal_10278 ), .Q ( new_AGEMA_signal_10279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5802 ( .C ( clk ), .D ( new_AGEMA_signal_10290 ), .Q ( new_AGEMA_signal_10291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5816 ( .C ( clk ), .D ( new_AGEMA_signal_10304 ), .Q ( new_AGEMA_signal_10305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5830 ( .C ( clk ), .D ( new_AGEMA_signal_10318 ), .Q ( new_AGEMA_signal_10319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5884 ( .C ( clk ), .D ( new_AGEMA_signal_10372 ), .Q ( new_AGEMA_signal_10373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5892 ( .C ( clk ), .D ( new_AGEMA_signal_10380 ), .Q ( new_AGEMA_signal_10381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5900 ( .C ( clk ), .D ( new_AGEMA_signal_10388 ), .Q ( new_AGEMA_signal_10389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5908 ( .C ( clk ), .D ( new_AGEMA_signal_10396 ), .Q ( new_AGEMA_signal_10397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5916 ( .C ( clk ), .D ( new_AGEMA_signal_10404 ), .Q ( new_AGEMA_signal_10405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5924 ( .C ( clk ), .D ( new_AGEMA_signal_10412 ), .Q ( new_AGEMA_signal_10413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5932 ( .C ( clk ), .D ( new_AGEMA_signal_10420 ), .Q ( new_AGEMA_signal_10421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5940 ( .C ( clk ), .D ( new_AGEMA_signal_10428 ), .Q ( new_AGEMA_signal_10429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5948 ( .C ( clk ), .D ( new_AGEMA_signal_10436 ), .Q ( new_AGEMA_signal_10437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5956 ( .C ( clk ), .D ( new_AGEMA_signal_10444 ), .Q ( new_AGEMA_signal_10445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5964 ( .C ( clk ), .D ( new_AGEMA_signal_10452 ), .Q ( new_AGEMA_signal_10453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5972 ( .C ( clk ), .D ( new_AGEMA_signal_10460 ), .Q ( new_AGEMA_signal_10461 ) ) ;

    /* cells in depth 29 */
    buf_clk new_AGEMA_reg_buffer_5763 ( .C ( clk ), .D ( new_AGEMA_signal_10251 ), .Q ( new_AGEMA_signal_10252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5777 ( .C ( clk ), .D ( new_AGEMA_signal_10265 ), .Q ( new_AGEMA_signal_10266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5791 ( .C ( clk ), .D ( new_AGEMA_signal_10279 ), .Q ( new_AGEMA_signal_10280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5803 ( .C ( clk ), .D ( new_AGEMA_signal_10291 ), .Q ( new_AGEMA_signal_10292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5817 ( .C ( clk ), .D ( new_AGEMA_signal_10305 ), .Q ( new_AGEMA_signal_10306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5831 ( .C ( clk ), .D ( new_AGEMA_signal_10319 ), .Q ( new_AGEMA_signal_10320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5835 ( .C ( clk ), .D ( N169 ), .Q ( new_AGEMA_signal_10324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5841 ( .C ( clk ), .D ( new_AGEMA_signal_2780 ), .Q ( new_AGEMA_signal_10330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5847 ( .C ( clk ), .D ( new_AGEMA_signal_2781 ), .Q ( new_AGEMA_signal_10336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5853 ( .C ( clk ), .D ( N277 ), .Q ( new_AGEMA_signal_10342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5859 ( .C ( clk ), .D ( new_AGEMA_signal_2782 ), .Q ( new_AGEMA_signal_10348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5865 ( .C ( clk ), .D ( new_AGEMA_signal_2783 ), .Q ( new_AGEMA_signal_10354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5885 ( .C ( clk ), .D ( new_AGEMA_signal_10373 ), .Q ( new_AGEMA_signal_10374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5893 ( .C ( clk ), .D ( new_AGEMA_signal_10381 ), .Q ( new_AGEMA_signal_10382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5901 ( .C ( clk ), .D ( new_AGEMA_signal_10389 ), .Q ( new_AGEMA_signal_10390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5909 ( .C ( clk ), .D ( new_AGEMA_signal_10397 ), .Q ( new_AGEMA_signal_10398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5917 ( .C ( clk ), .D ( new_AGEMA_signal_10405 ), .Q ( new_AGEMA_signal_10406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5925 ( .C ( clk ), .D ( new_AGEMA_signal_10413 ), .Q ( new_AGEMA_signal_10414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5933 ( .C ( clk ), .D ( new_AGEMA_signal_10421 ), .Q ( new_AGEMA_signal_10422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5941 ( .C ( clk ), .D ( new_AGEMA_signal_10429 ), .Q ( new_AGEMA_signal_10430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5949 ( .C ( clk ), .D ( new_AGEMA_signal_10437 ), .Q ( new_AGEMA_signal_10438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5957 ( .C ( clk ), .D ( new_AGEMA_signal_10445 ), .Q ( new_AGEMA_signal_10446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5965 ( .C ( clk ), .D ( new_AGEMA_signal_10453 ), .Q ( new_AGEMA_signal_10454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5973 ( .C ( clk ), .D ( new_AGEMA_signal_10461 ), .Q ( new_AGEMA_signal_10462 ) ) ;

    /* cells in depth 30 */
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2377 ( .a ({new_AGEMA_signal_10203, new_AGEMA_signal_10195, new_AGEMA_signal_10187}), .b ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, n2211}), .clk ( clk ), .r ({Fresh[2594], Fresh[2593], Fresh[2592]}), .c ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, N379}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2541 ( .a ({new_AGEMA_signal_10239, new_AGEMA_signal_10227, new_AGEMA_signal_10215}), .b ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, n2379}), .clk ( clk ), .r ({Fresh[2597], Fresh[2596], Fresh[2595]}), .c ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, n2381}) ) ;
    buf_clk new_AGEMA_reg_buffer_5764 ( .C ( clk ), .D ( new_AGEMA_signal_10252 ), .Q ( new_AGEMA_signal_10253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5778 ( .C ( clk ), .D ( new_AGEMA_signal_10266 ), .Q ( new_AGEMA_signal_10267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5792 ( .C ( clk ), .D ( new_AGEMA_signal_10280 ), .Q ( new_AGEMA_signal_10281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5804 ( .C ( clk ), .D ( new_AGEMA_signal_10292 ), .Q ( new_AGEMA_signal_10293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5818 ( .C ( clk ), .D ( new_AGEMA_signal_10306 ), .Q ( new_AGEMA_signal_10307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5832 ( .C ( clk ), .D ( new_AGEMA_signal_10320 ), .Q ( new_AGEMA_signal_10321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5836 ( .C ( clk ), .D ( new_AGEMA_signal_10324 ), .Q ( new_AGEMA_signal_10325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5842 ( .C ( clk ), .D ( new_AGEMA_signal_10330 ), .Q ( new_AGEMA_signal_10331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5848 ( .C ( clk ), .D ( new_AGEMA_signal_10336 ), .Q ( new_AGEMA_signal_10337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5854 ( .C ( clk ), .D ( new_AGEMA_signal_10342 ), .Q ( new_AGEMA_signal_10343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5860 ( .C ( clk ), .D ( new_AGEMA_signal_10348 ), .Q ( new_AGEMA_signal_10349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5866 ( .C ( clk ), .D ( new_AGEMA_signal_10354 ), .Q ( new_AGEMA_signal_10355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5886 ( .C ( clk ), .D ( new_AGEMA_signal_10374 ), .Q ( new_AGEMA_signal_10375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5894 ( .C ( clk ), .D ( new_AGEMA_signal_10382 ), .Q ( new_AGEMA_signal_10383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5902 ( .C ( clk ), .D ( new_AGEMA_signal_10390 ), .Q ( new_AGEMA_signal_10391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5910 ( .C ( clk ), .D ( new_AGEMA_signal_10398 ), .Q ( new_AGEMA_signal_10399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5918 ( .C ( clk ), .D ( new_AGEMA_signal_10406 ), .Q ( new_AGEMA_signal_10407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5926 ( .C ( clk ), .D ( new_AGEMA_signal_10414 ), .Q ( new_AGEMA_signal_10415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5934 ( .C ( clk ), .D ( new_AGEMA_signal_10422 ), .Q ( new_AGEMA_signal_10423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5942 ( .C ( clk ), .D ( new_AGEMA_signal_10430 ), .Q ( new_AGEMA_signal_10431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5950 ( .C ( clk ), .D ( new_AGEMA_signal_10438 ), .Q ( new_AGEMA_signal_10439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5958 ( .C ( clk ), .D ( new_AGEMA_signal_10446 ), .Q ( new_AGEMA_signal_10447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5966 ( .C ( clk ), .D ( new_AGEMA_signal_10454 ), .Q ( new_AGEMA_signal_10455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5974 ( .C ( clk ), .D ( new_AGEMA_signal_10462 ), .Q ( new_AGEMA_signal_10463 ) ) ;

    /* cells in depth 31 */
    buf_clk new_AGEMA_reg_buffer_5805 ( .C ( clk ), .D ( new_AGEMA_signal_10293 ), .Q ( new_AGEMA_signal_10294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5819 ( .C ( clk ), .D ( new_AGEMA_signal_10307 ), .Q ( new_AGEMA_signal_10308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5833 ( .C ( clk ), .D ( new_AGEMA_signal_10321 ), .Q ( new_AGEMA_signal_10322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5837 ( .C ( clk ), .D ( new_AGEMA_signal_10325 ), .Q ( new_AGEMA_signal_10326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5843 ( .C ( clk ), .D ( new_AGEMA_signal_10331 ), .Q ( new_AGEMA_signal_10332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5849 ( .C ( clk ), .D ( new_AGEMA_signal_10337 ), .Q ( new_AGEMA_signal_10338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5855 ( .C ( clk ), .D ( new_AGEMA_signal_10343 ), .Q ( new_AGEMA_signal_10344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5861 ( .C ( clk ), .D ( new_AGEMA_signal_10349 ), .Q ( new_AGEMA_signal_10350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5867 ( .C ( clk ), .D ( new_AGEMA_signal_10355 ), .Q ( new_AGEMA_signal_10356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5871 ( .C ( clk ), .D ( N379 ), .Q ( new_AGEMA_signal_10360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5875 ( .C ( clk ), .D ( new_AGEMA_signal_2788 ), .Q ( new_AGEMA_signal_10364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5879 ( .C ( clk ), .D ( new_AGEMA_signal_2789 ), .Q ( new_AGEMA_signal_10368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5887 ( .C ( clk ), .D ( new_AGEMA_signal_10375 ), .Q ( new_AGEMA_signal_10376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5895 ( .C ( clk ), .D ( new_AGEMA_signal_10383 ), .Q ( new_AGEMA_signal_10384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5903 ( .C ( clk ), .D ( new_AGEMA_signal_10391 ), .Q ( new_AGEMA_signal_10392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5911 ( .C ( clk ), .D ( new_AGEMA_signal_10399 ), .Q ( new_AGEMA_signal_10400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5919 ( .C ( clk ), .D ( new_AGEMA_signal_10407 ), .Q ( new_AGEMA_signal_10408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5927 ( .C ( clk ), .D ( new_AGEMA_signal_10415 ), .Q ( new_AGEMA_signal_10416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5935 ( .C ( clk ), .D ( new_AGEMA_signal_10423 ), .Q ( new_AGEMA_signal_10424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5943 ( .C ( clk ), .D ( new_AGEMA_signal_10431 ), .Q ( new_AGEMA_signal_10432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5951 ( .C ( clk ), .D ( new_AGEMA_signal_10439 ), .Q ( new_AGEMA_signal_10440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5959 ( .C ( clk ), .D ( new_AGEMA_signal_10447 ), .Q ( new_AGEMA_signal_10448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5967 ( .C ( clk ), .D ( new_AGEMA_signal_10455 ), .Q ( new_AGEMA_signal_10456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5975 ( .C ( clk ), .D ( new_AGEMA_signal_10463 ), .Q ( new_AGEMA_signal_10464 ) ) ;

    /* cells in depth 32 */
    nor_HPC2 #(.security_order(2), .pipeline(1)) U2542 ( .a ({new_AGEMA_signal_10281, new_AGEMA_signal_10267, new_AGEMA_signal_10253}), .b ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, n2381}), .clk ( clk ), .r ({Fresh[2600], Fresh[2599], Fresh[2598]}), .c ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, n2427}) ) ;
    buf_clk new_AGEMA_reg_buffer_5806 ( .C ( clk ), .D ( new_AGEMA_signal_10294 ), .Q ( new_AGEMA_signal_10295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5820 ( .C ( clk ), .D ( new_AGEMA_signal_10308 ), .Q ( new_AGEMA_signal_10309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5834 ( .C ( clk ), .D ( new_AGEMA_signal_10322 ), .Q ( new_AGEMA_signal_10323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5838 ( .C ( clk ), .D ( new_AGEMA_signal_10326 ), .Q ( new_AGEMA_signal_10327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5844 ( .C ( clk ), .D ( new_AGEMA_signal_10332 ), .Q ( new_AGEMA_signal_10333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5850 ( .C ( clk ), .D ( new_AGEMA_signal_10338 ), .Q ( new_AGEMA_signal_10339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5856 ( .C ( clk ), .D ( new_AGEMA_signal_10344 ), .Q ( new_AGEMA_signal_10345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5862 ( .C ( clk ), .D ( new_AGEMA_signal_10350 ), .Q ( new_AGEMA_signal_10351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5868 ( .C ( clk ), .D ( new_AGEMA_signal_10356 ), .Q ( new_AGEMA_signal_10357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5872 ( .C ( clk ), .D ( new_AGEMA_signal_10360 ), .Q ( new_AGEMA_signal_10361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5876 ( .C ( clk ), .D ( new_AGEMA_signal_10364 ), .Q ( new_AGEMA_signal_10365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5880 ( .C ( clk ), .D ( new_AGEMA_signal_10368 ), .Q ( new_AGEMA_signal_10369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5888 ( .C ( clk ), .D ( new_AGEMA_signal_10376 ), .Q ( new_AGEMA_signal_10377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5896 ( .C ( clk ), .D ( new_AGEMA_signal_10384 ), .Q ( new_AGEMA_signal_10385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5904 ( .C ( clk ), .D ( new_AGEMA_signal_10392 ), .Q ( new_AGEMA_signal_10393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5912 ( .C ( clk ), .D ( new_AGEMA_signal_10400 ), .Q ( new_AGEMA_signal_10401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5920 ( .C ( clk ), .D ( new_AGEMA_signal_10408 ), .Q ( new_AGEMA_signal_10409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5928 ( .C ( clk ), .D ( new_AGEMA_signal_10416 ), .Q ( new_AGEMA_signal_10417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5936 ( .C ( clk ), .D ( new_AGEMA_signal_10424 ), .Q ( new_AGEMA_signal_10425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5944 ( .C ( clk ), .D ( new_AGEMA_signal_10432 ), .Q ( new_AGEMA_signal_10433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5952 ( .C ( clk ), .D ( new_AGEMA_signal_10440 ), .Q ( new_AGEMA_signal_10441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5960 ( .C ( clk ), .D ( new_AGEMA_signal_10448 ), .Q ( new_AGEMA_signal_10449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5968 ( .C ( clk ), .D ( new_AGEMA_signal_10456 ), .Q ( new_AGEMA_signal_10457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5976 ( .C ( clk ), .D ( new_AGEMA_signal_10464 ), .Q ( new_AGEMA_signal_10465 ) ) ;

    /* cells in depth 33 */
    buf_clk new_AGEMA_reg_buffer_5839 ( .C ( clk ), .D ( new_AGEMA_signal_10327 ), .Q ( new_AGEMA_signal_10328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5845 ( .C ( clk ), .D ( new_AGEMA_signal_10333 ), .Q ( new_AGEMA_signal_10334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5851 ( .C ( clk ), .D ( new_AGEMA_signal_10339 ), .Q ( new_AGEMA_signal_10340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5857 ( .C ( clk ), .D ( new_AGEMA_signal_10345 ), .Q ( new_AGEMA_signal_10346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5863 ( .C ( clk ), .D ( new_AGEMA_signal_10351 ), .Q ( new_AGEMA_signal_10352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5869 ( .C ( clk ), .D ( new_AGEMA_signal_10357 ), .Q ( new_AGEMA_signal_10358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5873 ( .C ( clk ), .D ( new_AGEMA_signal_10361 ), .Q ( new_AGEMA_signal_10362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5877 ( .C ( clk ), .D ( new_AGEMA_signal_10365 ), .Q ( new_AGEMA_signal_10366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5881 ( .C ( clk ), .D ( new_AGEMA_signal_10369 ), .Q ( new_AGEMA_signal_10370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5889 ( .C ( clk ), .D ( new_AGEMA_signal_10377 ), .Q ( new_AGEMA_signal_10378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5897 ( .C ( clk ), .D ( new_AGEMA_signal_10385 ), .Q ( new_AGEMA_signal_10386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5905 ( .C ( clk ), .D ( new_AGEMA_signal_10393 ), .Q ( new_AGEMA_signal_10394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5913 ( .C ( clk ), .D ( new_AGEMA_signal_10401 ), .Q ( new_AGEMA_signal_10402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5921 ( .C ( clk ), .D ( new_AGEMA_signal_10409 ), .Q ( new_AGEMA_signal_10410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5929 ( .C ( clk ), .D ( new_AGEMA_signal_10417 ), .Q ( new_AGEMA_signal_10418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5937 ( .C ( clk ), .D ( new_AGEMA_signal_10425 ), .Q ( new_AGEMA_signal_10426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5945 ( .C ( clk ), .D ( new_AGEMA_signal_10433 ), .Q ( new_AGEMA_signal_10434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5953 ( .C ( clk ), .D ( new_AGEMA_signal_10441 ), .Q ( new_AGEMA_signal_10442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5961 ( .C ( clk ), .D ( new_AGEMA_signal_10449 ), .Q ( new_AGEMA_signal_10450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5969 ( .C ( clk ), .D ( new_AGEMA_signal_10457 ), .Q ( new_AGEMA_signal_10458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5977 ( .C ( clk ), .D ( new_AGEMA_signal_10465 ), .Q ( new_AGEMA_signal_10466 ) ) ;

    /* cells in depth 34 */
    nand_HPC2 #(.security_order(2), .pipeline(1)) U2584 ( .a ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, n2427}), .b ({new_AGEMA_signal_10323, new_AGEMA_signal_10309, new_AGEMA_signal_10295}), .clk ( clk ), .r ({Fresh[2603], Fresh[2602], Fresh[2601]}), .c ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, N563}) ) ;
    buf_clk new_AGEMA_reg_buffer_5840 ( .C ( clk ), .D ( new_AGEMA_signal_10328 ), .Q ( new_AGEMA_signal_10329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5846 ( .C ( clk ), .D ( new_AGEMA_signal_10334 ), .Q ( new_AGEMA_signal_10335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5852 ( .C ( clk ), .D ( new_AGEMA_signal_10340 ), .Q ( new_AGEMA_signal_10341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5858 ( .C ( clk ), .D ( new_AGEMA_signal_10346 ), .Q ( new_AGEMA_signal_10347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5864 ( .C ( clk ), .D ( new_AGEMA_signal_10352 ), .Q ( new_AGEMA_signal_10353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5870 ( .C ( clk ), .D ( new_AGEMA_signal_10358 ), .Q ( new_AGEMA_signal_10359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5874 ( .C ( clk ), .D ( new_AGEMA_signal_10362 ), .Q ( new_AGEMA_signal_10363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5878 ( .C ( clk ), .D ( new_AGEMA_signal_10366 ), .Q ( new_AGEMA_signal_10367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5882 ( .C ( clk ), .D ( new_AGEMA_signal_10370 ), .Q ( new_AGEMA_signal_10371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5890 ( .C ( clk ), .D ( new_AGEMA_signal_10378 ), .Q ( new_AGEMA_signal_10379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5898 ( .C ( clk ), .D ( new_AGEMA_signal_10386 ), .Q ( new_AGEMA_signal_10387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5906 ( .C ( clk ), .D ( new_AGEMA_signal_10394 ), .Q ( new_AGEMA_signal_10395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5914 ( .C ( clk ), .D ( new_AGEMA_signal_10402 ), .Q ( new_AGEMA_signal_10403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5922 ( .C ( clk ), .D ( new_AGEMA_signal_10410 ), .Q ( new_AGEMA_signal_10411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5930 ( .C ( clk ), .D ( new_AGEMA_signal_10418 ), .Q ( new_AGEMA_signal_10419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5938 ( .C ( clk ), .D ( new_AGEMA_signal_10426 ), .Q ( new_AGEMA_signal_10427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5946 ( .C ( clk ), .D ( new_AGEMA_signal_10434 ), .Q ( new_AGEMA_signal_10435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5954 ( .C ( clk ), .D ( new_AGEMA_signal_10442 ), .Q ( new_AGEMA_signal_10443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5962 ( .C ( clk ), .D ( new_AGEMA_signal_10450 ), .Q ( new_AGEMA_signal_10451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5970 ( .C ( clk ), .D ( new_AGEMA_signal_10458 ), .Q ( new_AGEMA_signal_10459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5978 ( .C ( clk ), .D ( new_AGEMA_signal_10466 ), .Q ( new_AGEMA_signal_10467 ) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(1)) SO_reg_7_ ( .clk ( clk ), .D ({new_AGEMA_signal_10341, new_AGEMA_signal_10335, new_AGEMA_signal_10329}), .Q ({SO_s2[7], SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) SO_reg_6_ ( .clk ( clk ), .D ({new_AGEMA_signal_10359, new_AGEMA_signal_10353, new_AGEMA_signal_10347}), .Q ({SO_s2[6], SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) SO_reg_5_ ( .clk ( clk ), .D ({new_AGEMA_signal_10371, new_AGEMA_signal_10367, new_AGEMA_signal_10363}), .Q ({SO_s2[5], SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) SO_reg_4_ ( .clk ( clk ), .D ({new_AGEMA_signal_10395, new_AGEMA_signal_10387, new_AGEMA_signal_10379}), .Q ({SO_s2[4], SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) SO_reg_3_ ( .clk ( clk ), .D ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, N563}), .Q ({SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) SO_reg_2_ ( .clk ( clk ), .D ({new_AGEMA_signal_10419, new_AGEMA_signal_10411, new_AGEMA_signal_10403}), .Q ({SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) SO_reg_1_ ( .clk ( clk ), .D ({new_AGEMA_signal_10443, new_AGEMA_signal_10435, new_AGEMA_signal_10427}), .Q ({SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) SO_reg_0_ ( .clk ( clk ), .D ({new_AGEMA_signal_10467, new_AGEMA_signal_10459, new_AGEMA_signal_10451}), .Q ({SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
