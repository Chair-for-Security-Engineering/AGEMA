/* modified netlist. Source: module AES in file AES.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module AES_HPC3_Pipeline_d3 (plaintext_s0, key_s0, clk, reset, plaintext_s1, plaintext_s2, plaintext_s3, key_s1, key_s2, key_s3, Fresh, ciphertext_s0, done, ciphertext_s1, ciphertext_s2, ciphertext_s3);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] plaintext_s1 ;
    input [127:0] plaintext_s2 ;
    input [127:0] plaintext_s3 ;
    input [127:0] key_s1 ;
    input [127:0] key_s2 ;
    input [127:0] key_s3 ;
    input [1631:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output [127:0] ciphertext_s2 ;
    output [127:0] ciphertext_s3 ;
    wire AKSRnotDone ;
    wire LastRoundorDone ;
    wire n44 ;
    wire n45 ;
    wire n46 ;
    wire n47 ;
    wire n48 ;
    wire n49 ;
    wire n50 ;
    wire n51 ;
    wire n52 ;
    wire n53 ;
    wire n54 ;
    wire n55 ;
    wire n56 ;
    wire n57 ;
    wire n58 ;
    wire n59 ;
    wire n60 ;
    wire n61 ;
    wire n62 ;
    wire RoundReg_Inst_ff_SDE_0_next_state ;
    wire RoundReg_Inst_ff_SDE_1_next_state ;
    wire RoundReg_Inst_ff_SDE_2_next_state ;
    wire RoundReg_Inst_ff_SDE_3_next_state ;
    wire RoundReg_Inst_ff_SDE_4_next_state ;
    wire RoundReg_Inst_ff_SDE_5_next_state ;
    wire RoundReg_Inst_ff_SDE_6_next_state ;
    wire RoundReg_Inst_ff_SDE_7_next_state ;
    wire RoundReg_Inst_ff_SDE_8_next_state ;
    wire RoundReg_Inst_ff_SDE_9_next_state ;
    wire RoundReg_Inst_ff_SDE_10_next_state ;
    wire RoundReg_Inst_ff_SDE_11_next_state ;
    wire RoundReg_Inst_ff_SDE_12_next_state ;
    wire RoundReg_Inst_ff_SDE_13_next_state ;
    wire RoundReg_Inst_ff_SDE_14_next_state ;
    wire RoundReg_Inst_ff_SDE_15_next_state ;
    wire RoundReg_Inst_ff_SDE_16_next_state ;
    wire RoundReg_Inst_ff_SDE_17_next_state ;
    wire RoundReg_Inst_ff_SDE_18_next_state ;
    wire RoundReg_Inst_ff_SDE_19_next_state ;
    wire RoundReg_Inst_ff_SDE_20_next_state ;
    wire RoundReg_Inst_ff_SDE_21_next_state ;
    wire RoundReg_Inst_ff_SDE_22_next_state ;
    wire RoundReg_Inst_ff_SDE_23_next_state ;
    wire RoundReg_Inst_ff_SDE_24_next_state ;
    wire RoundReg_Inst_ff_SDE_25_next_state ;
    wire RoundReg_Inst_ff_SDE_26_next_state ;
    wire RoundReg_Inst_ff_SDE_27_next_state ;
    wire RoundReg_Inst_ff_SDE_28_next_state ;
    wire RoundReg_Inst_ff_SDE_29_next_state ;
    wire RoundReg_Inst_ff_SDE_30_next_state ;
    wire RoundReg_Inst_ff_SDE_31_next_state ;
    wire RoundReg_Inst_ff_SDE_32_next_state ;
    wire RoundReg_Inst_ff_SDE_33_next_state ;
    wire RoundReg_Inst_ff_SDE_34_next_state ;
    wire RoundReg_Inst_ff_SDE_35_next_state ;
    wire RoundReg_Inst_ff_SDE_36_next_state ;
    wire RoundReg_Inst_ff_SDE_37_next_state ;
    wire RoundReg_Inst_ff_SDE_38_next_state ;
    wire RoundReg_Inst_ff_SDE_39_next_state ;
    wire RoundReg_Inst_ff_SDE_40_next_state ;
    wire RoundReg_Inst_ff_SDE_41_next_state ;
    wire RoundReg_Inst_ff_SDE_42_next_state ;
    wire RoundReg_Inst_ff_SDE_43_next_state ;
    wire RoundReg_Inst_ff_SDE_44_next_state ;
    wire RoundReg_Inst_ff_SDE_45_next_state ;
    wire RoundReg_Inst_ff_SDE_46_next_state ;
    wire RoundReg_Inst_ff_SDE_47_next_state ;
    wire RoundReg_Inst_ff_SDE_48_next_state ;
    wire RoundReg_Inst_ff_SDE_49_next_state ;
    wire RoundReg_Inst_ff_SDE_50_next_state ;
    wire RoundReg_Inst_ff_SDE_51_next_state ;
    wire RoundReg_Inst_ff_SDE_52_next_state ;
    wire RoundReg_Inst_ff_SDE_53_next_state ;
    wire RoundReg_Inst_ff_SDE_54_next_state ;
    wire RoundReg_Inst_ff_SDE_55_next_state ;
    wire RoundReg_Inst_ff_SDE_56_next_state ;
    wire RoundReg_Inst_ff_SDE_57_next_state ;
    wire RoundReg_Inst_ff_SDE_58_next_state ;
    wire RoundReg_Inst_ff_SDE_59_next_state ;
    wire RoundReg_Inst_ff_SDE_60_next_state ;
    wire RoundReg_Inst_ff_SDE_61_next_state ;
    wire RoundReg_Inst_ff_SDE_62_next_state ;
    wire RoundReg_Inst_ff_SDE_63_next_state ;
    wire RoundReg_Inst_ff_SDE_64_next_state ;
    wire RoundReg_Inst_ff_SDE_65_next_state ;
    wire RoundReg_Inst_ff_SDE_66_next_state ;
    wire RoundReg_Inst_ff_SDE_67_next_state ;
    wire RoundReg_Inst_ff_SDE_68_next_state ;
    wire RoundReg_Inst_ff_SDE_69_next_state ;
    wire RoundReg_Inst_ff_SDE_70_next_state ;
    wire RoundReg_Inst_ff_SDE_71_next_state ;
    wire RoundReg_Inst_ff_SDE_72_next_state ;
    wire RoundReg_Inst_ff_SDE_73_next_state ;
    wire RoundReg_Inst_ff_SDE_74_next_state ;
    wire RoundReg_Inst_ff_SDE_75_next_state ;
    wire RoundReg_Inst_ff_SDE_76_next_state ;
    wire RoundReg_Inst_ff_SDE_77_next_state ;
    wire RoundReg_Inst_ff_SDE_78_next_state ;
    wire RoundReg_Inst_ff_SDE_79_next_state ;
    wire RoundReg_Inst_ff_SDE_80_next_state ;
    wire RoundReg_Inst_ff_SDE_81_next_state ;
    wire RoundReg_Inst_ff_SDE_82_next_state ;
    wire RoundReg_Inst_ff_SDE_83_next_state ;
    wire RoundReg_Inst_ff_SDE_84_next_state ;
    wire RoundReg_Inst_ff_SDE_85_next_state ;
    wire RoundReg_Inst_ff_SDE_86_next_state ;
    wire RoundReg_Inst_ff_SDE_87_next_state ;
    wire RoundReg_Inst_ff_SDE_88_next_state ;
    wire RoundReg_Inst_ff_SDE_89_next_state ;
    wire RoundReg_Inst_ff_SDE_90_next_state ;
    wire RoundReg_Inst_ff_SDE_91_next_state ;
    wire RoundReg_Inst_ff_SDE_92_next_state ;
    wire RoundReg_Inst_ff_SDE_93_next_state ;
    wire RoundReg_Inst_ff_SDE_94_next_state ;
    wire RoundReg_Inst_ff_SDE_95_next_state ;
    wire RoundReg_Inst_ff_SDE_96_next_state ;
    wire RoundReg_Inst_ff_SDE_97_next_state ;
    wire RoundReg_Inst_ff_SDE_98_next_state ;
    wire RoundReg_Inst_ff_SDE_99_next_state ;
    wire RoundReg_Inst_ff_SDE_100_next_state ;
    wire RoundReg_Inst_ff_SDE_101_next_state ;
    wire RoundReg_Inst_ff_SDE_102_next_state ;
    wire RoundReg_Inst_ff_SDE_103_next_state ;
    wire RoundReg_Inst_ff_SDE_104_next_state ;
    wire RoundReg_Inst_ff_SDE_105_next_state ;
    wire RoundReg_Inst_ff_SDE_106_next_state ;
    wire RoundReg_Inst_ff_SDE_107_next_state ;
    wire RoundReg_Inst_ff_SDE_108_next_state ;
    wire RoundReg_Inst_ff_SDE_109_next_state ;
    wire RoundReg_Inst_ff_SDE_110_next_state ;
    wire RoundReg_Inst_ff_SDE_111_next_state ;
    wire RoundReg_Inst_ff_SDE_112_next_state ;
    wire RoundReg_Inst_ff_SDE_113_next_state ;
    wire RoundReg_Inst_ff_SDE_114_next_state ;
    wire RoundReg_Inst_ff_SDE_115_next_state ;
    wire RoundReg_Inst_ff_SDE_116_next_state ;
    wire RoundReg_Inst_ff_SDE_117_next_state ;
    wire RoundReg_Inst_ff_SDE_118_next_state ;
    wire RoundReg_Inst_ff_SDE_119_next_state ;
    wire RoundReg_Inst_ff_SDE_120_next_state ;
    wire RoundReg_Inst_ff_SDE_121_next_state ;
    wire RoundReg_Inst_ff_SDE_122_next_state ;
    wire RoundReg_Inst_ff_SDE_123_next_state ;
    wire RoundReg_Inst_ff_SDE_124_next_state ;
    wire RoundReg_Inst_ff_SDE_125_next_state ;
    wire RoundReg_Inst_ff_SDE_126_next_state ;
    wire RoundReg_Inst_ff_SDE_127_next_state ;
    wire MuxSboxIn_n7 ;
    wire MuxSboxIn_n6 ;
    wire MuxSboxIn_n5 ;
    wire SubBytesIns_Inst_Sbox_0_L29 ;
    wire SubBytesIns_Inst_Sbox_0_L28 ;
    wire SubBytesIns_Inst_Sbox_0_L27 ;
    wire SubBytesIns_Inst_Sbox_0_L26 ;
    wire SubBytesIns_Inst_Sbox_0_L25 ;
    wire SubBytesIns_Inst_Sbox_0_L24 ;
    wire SubBytesIns_Inst_Sbox_0_L23 ;
    wire SubBytesIns_Inst_Sbox_0_L22 ;
    wire SubBytesIns_Inst_Sbox_0_L21 ;
    wire SubBytesIns_Inst_Sbox_0_L20 ;
    wire SubBytesIns_Inst_Sbox_0_L19 ;
    wire SubBytesIns_Inst_Sbox_0_L18 ;
    wire SubBytesIns_Inst_Sbox_0_L17 ;
    wire SubBytesIns_Inst_Sbox_0_L16 ;
    wire SubBytesIns_Inst_Sbox_0_L15 ;
    wire SubBytesIns_Inst_Sbox_0_L14 ;
    wire SubBytesIns_Inst_Sbox_0_L13 ;
    wire SubBytesIns_Inst_Sbox_0_L12 ;
    wire SubBytesIns_Inst_Sbox_0_L11 ;
    wire SubBytesIns_Inst_Sbox_0_L10 ;
    wire SubBytesIns_Inst_Sbox_0_L9 ;
    wire SubBytesIns_Inst_Sbox_0_L8 ;
    wire SubBytesIns_Inst_Sbox_0_L7 ;
    wire SubBytesIns_Inst_Sbox_0_L6 ;
    wire SubBytesIns_Inst_Sbox_0_L5 ;
    wire SubBytesIns_Inst_Sbox_0_L4 ;
    wire SubBytesIns_Inst_Sbox_0_L3 ;
    wire SubBytesIns_Inst_Sbox_0_L2 ;
    wire SubBytesIns_Inst_Sbox_0_L1 ;
    wire SubBytesIns_Inst_Sbox_0_L0 ;
    wire SubBytesIns_Inst_Sbox_0_M63 ;
    wire SubBytesIns_Inst_Sbox_0_M62 ;
    wire SubBytesIns_Inst_Sbox_0_M61 ;
    wire SubBytesIns_Inst_Sbox_0_M60 ;
    wire SubBytesIns_Inst_Sbox_0_M59 ;
    wire SubBytesIns_Inst_Sbox_0_M58 ;
    wire SubBytesIns_Inst_Sbox_0_M57 ;
    wire SubBytesIns_Inst_Sbox_0_M56 ;
    wire SubBytesIns_Inst_Sbox_0_M55 ;
    wire SubBytesIns_Inst_Sbox_0_M54 ;
    wire SubBytesIns_Inst_Sbox_0_M53 ;
    wire SubBytesIns_Inst_Sbox_0_M52 ;
    wire SubBytesIns_Inst_Sbox_0_M51 ;
    wire SubBytesIns_Inst_Sbox_0_M50 ;
    wire SubBytesIns_Inst_Sbox_0_M49 ;
    wire SubBytesIns_Inst_Sbox_0_M48 ;
    wire SubBytesIns_Inst_Sbox_0_M47 ;
    wire SubBytesIns_Inst_Sbox_0_M46 ;
    wire SubBytesIns_Inst_Sbox_0_M45 ;
    wire SubBytesIns_Inst_Sbox_0_M44 ;
    wire SubBytesIns_Inst_Sbox_0_M43 ;
    wire SubBytesIns_Inst_Sbox_0_M42 ;
    wire SubBytesIns_Inst_Sbox_0_M41 ;
    wire SubBytesIns_Inst_Sbox_0_M40 ;
    wire SubBytesIns_Inst_Sbox_0_M39 ;
    wire SubBytesIns_Inst_Sbox_0_M38 ;
    wire SubBytesIns_Inst_Sbox_0_M37 ;
    wire SubBytesIns_Inst_Sbox_0_M36 ;
    wire SubBytesIns_Inst_Sbox_0_M35 ;
    wire SubBytesIns_Inst_Sbox_0_M34 ;
    wire SubBytesIns_Inst_Sbox_0_M33 ;
    wire SubBytesIns_Inst_Sbox_0_M32 ;
    wire SubBytesIns_Inst_Sbox_0_M31 ;
    wire SubBytesIns_Inst_Sbox_0_M30 ;
    wire SubBytesIns_Inst_Sbox_0_M29 ;
    wire SubBytesIns_Inst_Sbox_0_M28 ;
    wire SubBytesIns_Inst_Sbox_0_M27 ;
    wire SubBytesIns_Inst_Sbox_0_M26 ;
    wire SubBytesIns_Inst_Sbox_0_M25 ;
    wire SubBytesIns_Inst_Sbox_0_M24 ;
    wire SubBytesIns_Inst_Sbox_0_M23 ;
    wire SubBytesIns_Inst_Sbox_0_M22 ;
    wire SubBytesIns_Inst_Sbox_0_M21 ;
    wire SubBytesIns_Inst_Sbox_0_M20 ;
    wire SubBytesIns_Inst_Sbox_0_M19 ;
    wire SubBytesIns_Inst_Sbox_0_M18 ;
    wire SubBytesIns_Inst_Sbox_0_M17 ;
    wire SubBytesIns_Inst_Sbox_0_M16 ;
    wire SubBytesIns_Inst_Sbox_0_M15 ;
    wire SubBytesIns_Inst_Sbox_0_M14 ;
    wire SubBytesIns_Inst_Sbox_0_M13 ;
    wire SubBytesIns_Inst_Sbox_0_M12 ;
    wire SubBytesIns_Inst_Sbox_0_M11 ;
    wire SubBytesIns_Inst_Sbox_0_M10 ;
    wire SubBytesIns_Inst_Sbox_0_M9 ;
    wire SubBytesIns_Inst_Sbox_0_M8 ;
    wire SubBytesIns_Inst_Sbox_0_M7 ;
    wire SubBytesIns_Inst_Sbox_0_M6 ;
    wire SubBytesIns_Inst_Sbox_0_M5 ;
    wire SubBytesIns_Inst_Sbox_0_M4 ;
    wire SubBytesIns_Inst_Sbox_0_M3 ;
    wire SubBytesIns_Inst_Sbox_0_M2 ;
    wire SubBytesIns_Inst_Sbox_0_M1 ;
    wire SubBytesIns_Inst_Sbox_0_T27 ;
    wire SubBytesIns_Inst_Sbox_0_T26 ;
    wire SubBytesIns_Inst_Sbox_0_T25 ;
    wire SubBytesIns_Inst_Sbox_0_T24 ;
    wire SubBytesIns_Inst_Sbox_0_T23 ;
    wire SubBytesIns_Inst_Sbox_0_T22 ;
    wire SubBytesIns_Inst_Sbox_0_T21 ;
    wire SubBytesIns_Inst_Sbox_0_T20 ;
    wire SubBytesIns_Inst_Sbox_0_T19 ;
    wire SubBytesIns_Inst_Sbox_0_T18 ;
    wire SubBytesIns_Inst_Sbox_0_T17 ;
    wire SubBytesIns_Inst_Sbox_0_T16 ;
    wire SubBytesIns_Inst_Sbox_0_T15 ;
    wire SubBytesIns_Inst_Sbox_0_T14 ;
    wire SubBytesIns_Inst_Sbox_0_T13 ;
    wire SubBytesIns_Inst_Sbox_0_T12 ;
    wire SubBytesIns_Inst_Sbox_0_T11 ;
    wire SubBytesIns_Inst_Sbox_0_T10 ;
    wire SubBytesIns_Inst_Sbox_0_T9 ;
    wire SubBytesIns_Inst_Sbox_0_T8 ;
    wire SubBytesIns_Inst_Sbox_0_T7 ;
    wire SubBytesIns_Inst_Sbox_0_T6 ;
    wire SubBytesIns_Inst_Sbox_0_T5 ;
    wire SubBytesIns_Inst_Sbox_0_T4 ;
    wire SubBytesIns_Inst_Sbox_0_T3 ;
    wire SubBytesIns_Inst_Sbox_0_T2 ;
    wire SubBytesIns_Inst_Sbox_0_T1 ;
    wire SubBytesIns_Inst_Sbox_1_L29 ;
    wire SubBytesIns_Inst_Sbox_1_L28 ;
    wire SubBytesIns_Inst_Sbox_1_L27 ;
    wire SubBytesIns_Inst_Sbox_1_L26 ;
    wire SubBytesIns_Inst_Sbox_1_L25 ;
    wire SubBytesIns_Inst_Sbox_1_L24 ;
    wire SubBytesIns_Inst_Sbox_1_L23 ;
    wire SubBytesIns_Inst_Sbox_1_L22 ;
    wire SubBytesIns_Inst_Sbox_1_L21 ;
    wire SubBytesIns_Inst_Sbox_1_L20 ;
    wire SubBytesIns_Inst_Sbox_1_L19 ;
    wire SubBytesIns_Inst_Sbox_1_L18 ;
    wire SubBytesIns_Inst_Sbox_1_L17 ;
    wire SubBytesIns_Inst_Sbox_1_L16 ;
    wire SubBytesIns_Inst_Sbox_1_L15 ;
    wire SubBytesIns_Inst_Sbox_1_L14 ;
    wire SubBytesIns_Inst_Sbox_1_L13 ;
    wire SubBytesIns_Inst_Sbox_1_L12 ;
    wire SubBytesIns_Inst_Sbox_1_L11 ;
    wire SubBytesIns_Inst_Sbox_1_L10 ;
    wire SubBytesIns_Inst_Sbox_1_L9 ;
    wire SubBytesIns_Inst_Sbox_1_L8 ;
    wire SubBytesIns_Inst_Sbox_1_L7 ;
    wire SubBytesIns_Inst_Sbox_1_L6 ;
    wire SubBytesIns_Inst_Sbox_1_L5 ;
    wire SubBytesIns_Inst_Sbox_1_L4 ;
    wire SubBytesIns_Inst_Sbox_1_L3 ;
    wire SubBytesIns_Inst_Sbox_1_L2 ;
    wire SubBytesIns_Inst_Sbox_1_L1 ;
    wire SubBytesIns_Inst_Sbox_1_L0 ;
    wire SubBytesIns_Inst_Sbox_1_M63 ;
    wire SubBytesIns_Inst_Sbox_1_M62 ;
    wire SubBytesIns_Inst_Sbox_1_M61 ;
    wire SubBytesIns_Inst_Sbox_1_M60 ;
    wire SubBytesIns_Inst_Sbox_1_M59 ;
    wire SubBytesIns_Inst_Sbox_1_M58 ;
    wire SubBytesIns_Inst_Sbox_1_M57 ;
    wire SubBytesIns_Inst_Sbox_1_M56 ;
    wire SubBytesIns_Inst_Sbox_1_M55 ;
    wire SubBytesIns_Inst_Sbox_1_M54 ;
    wire SubBytesIns_Inst_Sbox_1_M53 ;
    wire SubBytesIns_Inst_Sbox_1_M52 ;
    wire SubBytesIns_Inst_Sbox_1_M51 ;
    wire SubBytesIns_Inst_Sbox_1_M50 ;
    wire SubBytesIns_Inst_Sbox_1_M49 ;
    wire SubBytesIns_Inst_Sbox_1_M48 ;
    wire SubBytesIns_Inst_Sbox_1_M47 ;
    wire SubBytesIns_Inst_Sbox_1_M46 ;
    wire SubBytesIns_Inst_Sbox_1_M45 ;
    wire SubBytesIns_Inst_Sbox_1_M44 ;
    wire SubBytesIns_Inst_Sbox_1_M43 ;
    wire SubBytesIns_Inst_Sbox_1_M42 ;
    wire SubBytesIns_Inst_Sbox_1_M41 ;
    wire SubBytesIns_Inst_Sbox_1_M40 ;
    wire SubBytesIns_Inst_Sbox_1_M39 ;
    wire SubBytesIns_Inst_Sbox_1_M38 ;
    wire SubBytesIns_Inst_Sbox_1_M37 ;
    wire SubBytesIns_Inst_Sbox_1_M36 ;
    wire SubBytesIns_Inst_Sbox_1_M35 ;
    wire SubBytesIns_Inst_Sbox_1_M34 ;
    wire SubBytesIns_Inst_Sbox_1_M33 ;
    wire SubBytesIns_Inst_Sbox_1_M32 ;
    wire SubBytesIns_Inst_Sbox_1_M31 ;
    wire SubBytesIns_Inst_Sbox_1_M30 ;
    wire SubBytesIns_Inst_Sbox_1_M29 ;
    wire SubBytesIns_Inst_Sbox_1_M28 ;
    wire SubBytesIns_Inst_Sbox_1_M27 ;
    wire SubBytesIns_Inst_Sbox_1_M26 ;
    wire SubBytesIns_Inst_Sbox_1_M25 ;
    wire SubBytesIns_Inst_Sbox_1_M24 ;
    wire SubBytesIns_Inst_Sbox_1_M23 ;
    wire SubBytesIns_Inst_Sbox_1_M22 ;
    wire SubBytesIns_Inst_Sbox_1_M21 ;
    wire SubBytesIns_Inst_Sbox_1_M20 ;
    wire SubBytesIns_Inst_Sbox_1_M19 ;
    wire SubBytesIns_Inst_Sbox_1_M18 ;
    wire SubBytesIns_Inst_Sbox_1_M17 ;
    wire SubBytesIns_Inst_Sbox_1_M16 ;
    wire SubBytesIns_Inst_Sbox_1_M15 ;
    wire SubBytesIns_Inst_Sbox_1_M14 ;
    wire SubBytesIns_Inst_Sbox_1_M13 ;
    wire SubBytesIns_Inst_Sbox_1_M12 ;
    wire SubBytesIns_Inst_Sbox_1_M11 ;
    wire SubBytesIns_Inst_Sbox_1_M10 ;
    wire SubBytesIns_Inst_Sbox_1_M9 ;
    wire SubBytesIns_Inst_Sbox_1_M8 ;
    wire SubBytesIns_Inst_Sbox_1_M7 ;
    wire SubBytesIns_Inst_Sbox_1_M6 ;
    wire SubBytesIns_Inst_Sbox_1_M5 ;
    wire SubBytesIns_Inst_Sbox_1_M4 ;
    wire SubBytesIns_Inst_Sbox_1_M3 ;
    wire SubBytesIns_Inst_Sbox_1_M2 ;
    wire SubBytesIns_Inst_Sbox_1_M1 ;
    wire SubBytesIns_Inst_Sbox_1_T27 ;
    wire SubBytesIns_Inst_Sbox_1_T26 ;
    wire SubBytesIns_Inst_Sbox_1_T25 ;
    wire SubBytesIns_Inst_Sbox_1_T24 ;
    wire SubBytesIns_Inst_Sbox_1_T23 ;
    wire SubBytesIns_Inst_Sbox_1_T22 ;
    wire SubBytesIns_Inst_Sbox_1_T21 ;
    wire SubBytesIns_Inst_Sbox_1_T20 ;
    wire SubBytesIns_Inst_Sbox_1_T19 ;
    wire SubBytesIns_Inst_Sbox_1_T18 ;
    wire SubBytesIns_Inst_Sbox_1_T17 ;
    wire SubBytesIns_Inst_Sbox_1_T16 ;
    wire SubBytesIns_Inst_Sbox_1_T15 ;
    wire SubBytesIns_Inst_Sbox_1_T14 ;
    wire SubBytesIns_Inst_Sbox_1_T13 ;
    wire SubBytesIns_Inst_Sbox_1_T12 ;
    wire SubBytesIns_Inst_Sbox_1_T11 ;
    wire SubBytesIns_Inst_Sbox_1_T10 ;
    wire SubBytesIns_Inst_Sbox_1_T9 ;
    wire SubBytesIns_Inst_Sbox_1_T8 ;
    wire SubBytesIns_Inst_Sbox_1_T7 ;
    wire SubBytesIns_Inst_Sbox_1_T6 ;
    wire SubBytesIns_Inst_Sbox_1_T5 ;
    wire SubBytesIns_Inst_Sbox_1_T4 ;
    wire SubBytesIns_Inst_Sbox_1_T3 ;
    wire SubBytesIns_Inst_Sbox_1_T2 ;
    wire SubBytesIns_Inst_Sbox_1_T1 ;
    wire SubBytesIns_Inst_Sbox_2_L29 ;
    wire SubBytesIns_Inst_Sbox_2_L28 ;
    wire SubBytesIns_Inst_Sbox_2_L27 ;
    wire SubBytesIns_Inst_Sbox_2_L26 ;
    wire SubBytesIns_Inst_Sbox_2_L25 ;
    wire SubBytesIns_Inst_Sbox_2_L24 ;
    wire SubBytesIns_Inst_Sbox_2_L23 ;
    wire SubBytesIns_Inst_Sbox_2_L22 ;
    wire SubBytesIns_Inst_Sbox_2_L21 ;
    wire SubBytesIns_Inst_Sbox_2_L20 ;
    wire SubBytesIns_Inst_Sbox_2_L19 ;
    wire SubBytesIns_Inst_Sbox_2_L18 ;
    wire SubBytesIns_Inst_Sbox_2_L17 ;
    wire SubBytesIns_Inst_Sbox_2_L16 ;
    wire SubBytesIns_Inst_Sbox_2_L15 ;
    wire SubBytesIns_Inst_Sbox_2_L14 ;
    wire SubBytesIns_Inst_Sbox_2_L13 ;
    wire SubBytesIns_Inst_Sbox_2_L12 ;
    wire SubBytesIns_Inst_Sbox_2_L11 ;
    wire SubBytesIns_Inst_Sbox_2_L10 ;
    wire SubBytesIns_Inst_Sbox_2_L9 ;
    wire SubBytesIns_Inst_Sbox_2_L8 ;
    wire SubBytesIns_Inst_Sbox_2_L7 ;
    wire SubBytesIns_Inst_Sbox_2_L6 ;
    wire SubBytesIns_Inst_Sbox_2_L5 ;
    wire SubBytesIns_Inst_Sbox_2_L4 ;
    wire SubBytesIns_Inst_Sbox_2_L3 ;
    wire SubBytesIns_Inst_Sbox_2_L2 ;
    wire SubBytesIns_Inst_Sbox_2_L1 ;
    wire SubBytesIns_Inst_Sbox_2_L0 ;
    wire SubBytesIns_Inst_Sbox_2_M63 ;
    wire SubBytesIns_Inst_Sbox_2_M62 ;
    wire SubBytesIns_Inst_Sbox_2_M61 ;
    wire SubBytesIns_Inst_Sbox_2_M60 ;
    wire SubBytesIns_Inst_Sbox_2_M59 ;
    wire SubBytesIns_Inst_Sbox_2_M58 ;
    wire SubBytesIns_Inst_Sbox_2_M57 ;
    wire SubBytesIns_Inst_Sbox_2_M56 ;
    wire SubBytesIns_Inst_Sbox_2_M55 ;
    wire SubBytesIns_Inst_Sbox_2_M54 ;
    wire SubBytesIns_Inst_Sbox_2_M53 ;
    wire SubBytesIns_Inst_Sbox_2_M52 ;
    wire SubBytesIns_Inst_Sbox_2_M51 ;
    wire SubBytesIns_Inst_Sbox_2_M50 ;
    wire SubBytesIns_Inst_Sbox_2_M49 ;
    wire SubBytesIns_Inst_Sbox_2_M48 ;
    wire SubBytesIns_Inst_Sbox_2_M47 ;
    wire SubBytesIns_Inst_Sbox_2_M46 ;
    wire SubBytesIns_Inst_Sbox_2_M45 ;
    wire SubBytesIns_Inst_Sbox_2_M44 ;
    wire SubBytesIns_Inst_Sbox_2_M43 ;
    wire SubBytesIns_Inst_Sbox_2_M42 ;
    wire SubBytesIns_Inst_Sbox_2_M41 ;
    wire SubBytesIns_Inst_Sbox_2_M40 ;
    wire SubBytesIns_Inst_Sbox_2_M39 ;
    wire SubBytesIns_Inst_Sbox_2_M38 ;
    wire SubBytesIns_Inst_Sbox_2_M37 ;
    wire SubBytesIns_Inst_Sbox_2_M36 ;
    wire SubBytesIns_Inst_Sbox_2_M35 ;
    wire SubBytesIns_Inst_Sbox_2_M34 ;
    wire SubBytesIns_Inst_Sbox_2_M33 ;
    wire SubBytesIns_Inst_Sbox_2_M32 ;
    wire SubBytesIns_Inst_Sbox_2_M31 ;
    wire SubBytesIns_Inst_Sbox_2_M30 ;
    wire SubBytesIns_Inst_Sbox_2_M29 ;
    wire SubBytesIns_Inst_Sbox_2_M28 ;
    wire SubBytesIns_Inst_Sbox_2_M27 ;
    wire SubBytesIns_Inst_Sbox_2_M26 ;
    wire SubBytesIns_Inst_Sbox_2_M25 ;
    wire SubBytesIns_Inst_Sbox_2_M24 ;
    wire SubBytesIns_Inst_Sbox_2_M23 ;
    wire SubBytesIns_Inst_Sbox_2_M22 ;
    wire SubBytesIns_Inst_Sbox_2_M21 ;
    wire SubBytesIns_Inst_Sbox_2_M20 ;
    wire SubBytesIns_Inst_Sbox_2_M19 ;
    wire SubBytesIns_Inst_Sbox_2_M18 ;
    wire SubBytesIns_Inst_Sbox_2_M17 ;
    wire SubBytesIns_Inst_Sbox_2_M16 ;
    wire SubBytesIns_Inst_Sbox_2_M15 ;
    wire SubBytesIns_Inst_Sbox_2_M14 ;
    wire SubBytesIns_Inst_Sbox_2_M13 ;
    wire SubBytesIns_Inst_Sbox_2_M12 ;
    wire SubBytesIns_Inst_Sbox_2_M11 ;
    wire SubBytesIns_Inst_Sbox_2_M10 ;
    wire SubBytesIns_Inst_Sbox_2_M9 ;
    wire SubBytesIns_Inst_Sbox_2_M8 ;
    wire SubBytesIns_Inst_Sbox_2_M7 ;
    wire SubBytesIns_Inst_Sbox_2_M6 ;
    wire SubBytesIns_Inst_Sbox_2_M5 ;
    wire SubBytesIns_Inst_Sbox_2_M4 ;
    wire SubBytesIns_Inst_Sbox_2_M3 ;
    wire SubBytesIns_Inst_Sbox_2_M2 ;
    wire SubBytesIns_Inst_Sbox_2_M1 ;
    wire SubBytesIns_Inst_Sbox_2_T27 ;
    wire SubBytesIns_Inst_Sbox_2_T26 ;
    wire SubBytesIns_Inst_Sbox_2_T25 ;
    wire SubBytesIns_Inst_Sbox_2_T24 ;
    wire SubBytesIns_Inst_Sbox_2_T23 ;
    wire SubBytesIns_Inst_Sbox_2_T22 ;
    wire SubBytesIns_Inst_Sbox_2_T21 ;
    wire SubBytesIns_Inst_Sbox_2_T20 ;
    wire SubBytesIns_Inst_Sbox_2_T19 ;
    wire SubBytesIns_Inst_Sbox_2_T18 ;
    wire SubBytesIns_Inst_Sbox_2_T17 ;
    wire SubBytesIns_Inst_Sbox_2_T16 ;
    wire SubBytesIns_Inst_Sbox_2_T15 ;
    wire SubBytesIns_Inst_Sbox_2_T14 ;
    wire SubBytesIns_Inst_Sbox_2_T13 ;
    wire SubBytesIns_Inst_Sbox_2_T12 ;
    wire SubBytesIns_Inst_Sbox_2_T11 ;
    wire SubBytesIns_Inst_Sbox_2_T10 ;
    wire SubBytesIns_Inst_Sbox_2_T9 ;
    wire SubBytesIns_Inst_Sbox_2_T8 ;
    wire SubBytesIns_Inst_Sbox_2_T7 ;
    wire SubBytesIns_Inst_Sbox_2_T6 ;
    wire SubBytesIns_Inst_Sbox_2_T5 ;
    wire SubBytesIns_Inst_Sbox_2_T4 ;
    wire SubBytesIns_Inst_Sbox_2_T3 ;
    wire SubBytesIns_Inst_Sbox_2_T2 ;
    wire SubBytesIns_Inst_Sbox_2_T1 ;
    wire SubBytesIns_Inst_Sbox_3_L29 ;
    wire SubBytesIns_Inst_Sbox_3_L28 ;
    wire SubBytesIns_Inst_Sbox_3_L27 ;
    wire SubBytesIns_Inst_Sbox_3_L26 ;
    wire SubBytesIns_Inst_Sbox_3_L25 ;
    wire SubBytesIns_Inst_Sbox_3_L24 ;
    wire SubBytesIns_Inst_Sbox_3_L23 ;
    wire SubBytesIns_Inst_Sbox_3_L22 ;
    wire SubBytesIns_Inst_Sbox_3_L21 ;
    wire SubBytesIns_Inst_Sbox_3_L20 ;
    wire SubBytesIns_Inst_Sbox_3_L19 ;
    wire SubBytesIns_Inst_Sbox_3_L18 ;
    wire SubBytesIns_Inst_Sbox_3_L17 ;
    wire SubBytesIns_Inst_Sbox_3_L16 ;
    wire SubBytesIns_Inst_Sbox_3_L15 ;
    wire SubBytesIns_Inst_Sbox_3_L14 ;
    wire SubBytesIns_Inst_Sbox_3_L13 ;
    wire SubBytesIns_Inst_Sbox_3_L12 ;
    wire SubBytesIns_Inst_Sbox_3_L11 ;
    wire SubBytesIns_Inst_Sbox_3_L10 ;
    wire SubBytesIns_Inst_Sbox_3_L9 ;
    wire SubBytesIns_Inst_Sbox_3_L8 ;
    wire SubBytesIns_Inst_Sbox_3_L7 ;
    wire SubBytesIns_Inst_Sbox_3_L6 ;
    wire SubBytesIns_Inst_Sbox_3_L5 ;
    wire SubBytesIns_Inst_Sbox_3_L4 ;
    wire SubBytesIns_Inst_Sbox_3_L3 ;
    wire SubBytesIns_Inst_Sbox_3_L2 ;
    wire SubBytesIns_Inst_Sbox_3_L1 ;
    wire SubBytesIns_Inst_Sbox_3_L0 ;
    wire SubBytesIns_Inst_Sbox_3_M63 ;
    wire SubBytesIns_Inst_Sbox_3_M62 ;
    wire SubBytesIns_Inst_Sbox_3_M61 ;
    wire SubBytesIns_Inst_Sbox_3_M60 ;
    wire SubBytesIns_Inst_Sbox_3_M59 ;
    wire SubBytesIns_Inst_Sbox_3_M58 ;
    wire SubBytesIns_Inst_Sbox_3_M57 ;
    wire SubBytesIns_Inst_Sbox_3_M56 ;
    wire SubBytesIns_Inst_Sbox_3_M55 ;
    wire SubBytesIns_Inst_Sbox_3_M54 ;
    wire SubBytesIns_Inst_Sbox_3_M53 ;
    wire SubBytesIns_Inst_Sbox_3_M52 ;
    wire SubBytesIns_Inst_Sbox_3_M51 ;
    wire SubBytesIns_Inst_Sbox_3_M50 ;
    wire SubBytesIns_Inst_Sbox_3_M49 ;
    wire SubBytesIns_Inst_Sbox_3_M48 ;
    wire SubBytesIns_Inst_Sbox_3_M47 ;
    wire SubBytesIns_Inst_Sbox_3_M46 ;
    wire SubBytesIns_Inst_Sbox_3_M45 ;
    wire SubBytesIns_Inst_Sbox_3_M44 ;
    wire SubBytesIns_Inst_Sbox_3_M43 ;
    wire SubBytesIns_Inst_Sbox_3_M42 ;
    wire SubBytesIns_Inst_Sbox_3_M41 ;
    wire SubBytesIns_Inst_Sbox_3_M40 ;
    wire SubBytesIns_Inst_Sbox_3_M39 ;
    wire SubBytesIns_Inst_Sbox_3_M38 ;
    wire SubBytesIns_Inst_Sbox_3_M37 ;
    wire SubBytesIns_Inst_Sbox_3_M36 ;
    wire SubBytesIns_Inst_Sbox_3_M35 ;
    wire SubBytesIns_Inst_Sbox_3_M34 ;
    wire SubBytesIns_Inst_Sbox_3_M33 ;
    wire SubBytesIns_Inst_Sbox_3_M32 ;
    wire SubBytesIns_Inst_Sbox_3_M31 ;
    wire SubBytesIns_Inst_Sbox_3_M30 ;
    wire SubBytesIns_Inst_Sbox_3_M29 ;
    wire SubBytesIns_Inst_Sbox_3_M28 ;
    wire SubBytesIns_Inst_Sbox_3_M27 ;
    wire SubBytesIns_Inst_Sbox_3_M26 ;
    wire SubBytesIns_Inst_Sbox_3_M25 ;
    wire SubBytesIns_Inst_Sbox_3_M24 ;
    wire SubBytesIns_Inst_Sbox_3_M23 ;
    wire SubBytesIns_Inst_Sbox_3_M22 ;
    wire SubBytesIns_Inst_Sbox_3_M21 ;
    wire SubBytesIns_Inst_Sbox_3_M20 ;
    wire SubBytesIns_Inst_Sbox_3_M19 ;
    wire SubBytesIns_Inst_Sbox_3_M18 ;
    wire SubBytesIns_Inst_Sbox_3_M17 ;
    wire SubBytesIns_Inst_Sbox_3_M16 ;
    wire SubBytesIns_Inst_Sbox_3_M15 ;
    wire SubBytesIns_Inst_Sbox_3_M14 ;
    wire SubBytesIns_Inst_Sbox_3_M13 ;
    wire SubBytesIns_Inst_Sbox_3_M12 ;
    wire SubBytesIns_Inst_Sbox_3_M11 ;
    wire SubBytesIns_Inst_Sbox_3_M10 ;
    wire SubBytesIns_Inst_Sbox_3_M9 ;
    wire SubBytesIns_Inst_Sbox_3_M8 ;
    wire SubBytesIns_Inst_Sbox_3_M7 ;
    wire SubBytesIns_Inst_Sbox_3_M6 ;
    wire SubBytesIns_Inst_Sbox_3_M5 ;
    wire SubBytesIns_Inst_Sbox_3_M4 ;
    wire SubBytesIns_Inst_Sbox_3_M3 ;
    wire SubBytesIns_Inst_Sbox_3_M2 ;
    wire SubBytesIns_Inst_Sbox_3_M1 ;
    wire SubBytesIns_Inst_Sbox_3_T27 ;
    wire SubBytesIns_Inst_Sbox_3_T26 ;
    wire SubBytesIns_Inst_Sbox_3_T25 ;
    wire SubBytesIns_Inst_Sbox_3_T24 ;
    wire SubBytesIns_Inst_Sbox_3_T23 ;
    wire SubBytesIns_Inst_Sbox_3_T22 ;
    wire SubBytesIns_Inst_Sbox_3_T21 ;
    wire SubBytesIns_Inst_Sbox_3_T20 ;
    wire SubBytesIns_Inst_Sbox_3_T19 ;
    wire SubBytesIns_Inst_Sbox_3_T18 ;
    wire SubBytesIns_Inst_Sbox_3_T17 ;
    wire SubBytesIns_Inst_Sbox_3_T16 ;
    wire SubBytesIns_Inst_Sbox_3_T15 ;
    wire SubBytesIns_Inst_Sbox_3_T14 ;
    wire SubBytesIns_Inst_Sbox_3_T13 ;
    wire SubBytesIns_Inst_Sbox_3_T12 ;
    wire SubBytesIns_Inst_Sbox_3_T11 ;
    wire SubBytesIns_Inst_Sbox_3_T10 ;
    wire SubBytesIns_Inst_Sbox_3_T9 ;
    wire SubBytesIns_Inst_Sbox_3_T8 ;
    wire SubBytesIns_Inst_Sbox_3_T7 ;
    wire SubBytesIns_Inst_Sbox_3_T6 ;
    wire SubBytesIns_Inst_Sbox_3_T5 ;
    wire SubBytesIns_Inst_Sbox_3_T4 ;
    wire SubBytesIns_Inst_Sbox_3_T3 ;
    wire SubBytesIns_Inst_Sbox_3_T2 ;
    wire SubBytesIns_Inst_Sbox_3_T1 ;
    wire MixColumnsIns_n64 ;
    wire MixColumnsIns_n63 ;
    wire MixColumnsIns_n62 ;
    wire MixColumnsIns_n61 ;
    wire MixColumnsIns_n60 ;
    wire MixColumnsIns_n59 ;
    wire MixColumnsIns_n58 ;
    wire MixColumnsIns_n57 ;
    wire MixColumnsIns_n56 ;
    wire MixColumnsIns_n55 ;
    wire MixColumnsIns_n54 ;
    wire MixColumnsIns_n53 ;
    wire MixColumnsIns_n52 ;
    wire MixColumnsIns_n51 ;
    wire MixColumnsIns_n50 ;
    wire MixColumnsIns_n49 ;
    wire MixColumnsIns_n48 ;
    wire MixColumnsIns_n47 ;
    wire MixColumnsIns_n46 ;
    wire MixColumnsIns_n45 ;
    wire MixColumnsIns_n44 ;
    wire MixColumnsIns_n43 ;
    wire MixColumnsIns_n42 ;
    wire MixColumnsIns_n41 ;
    wire MixColumnsIns_n40 ;
    wire MixColumnsIns_n39 ;
    wire MixColumnsIns_n38 ;
    wire MixColumnsIns_n37 ;
    wire MixColumnsIns_n36 ;
    wire MixColumnsIns_n35 ;
    wire MixColumnsIns_n34 ;
    wire MixColumnsIns_n33 ;
    wire MixColumnsIns_n32 ;
    wire MixColumnsIns_n31 ;
    wire MixColumnsIns_n30 ;
    wire MixColumnsIns_n29 ;
    wire MixColumnsIns_n28 ;
    wire MixColumnsIns_n27 ;
    wire MixColumnsIns_n26 ;
    wire MixColumnsIns_n25 ;
    wire MixColumnsIns_n24 ;
    wire MixColumnsIns_n23 ;
    wire MixColumnsIns_n22 ;
    wire MixColumnsIns_n21 ;
    wire MixColumnsIns_n20 ;
    wire MixColumnsIns_n19 ;
    wire MixColumnsIns_n18 ;
    wire MixColumnsIns_n17 ;
    wire MixColumnsIns_n16 ;
    wire MixColumnsIns_n15 ;
    wire MixColumnsIns_n14 ;
    wire MixColumnsIns_n13 ;
    wire MixColumnsIns_n12 ;
    wire MixColumnsIns_n11 ;
    wire MixColumnsIns_n10 ;
    wire MixColumnsIns_n9 ;
    wire MixColumnsIns_n8 ;
    wire MixColumnsIns_n7 ;
    wire MixColumnsIns_n6 ;
    wire MixColumnsIns_n5 ;
    wire MixColumnsIns_n4 ;
    wire MixColumnsIns_n3 ;
    wire MixColumnsIns_n2 ;
    wire MixColumnsIns_n1 ;
    wire MuxMCOut_n6 ;
    wire MuxMCOut_n5 ;
    wire MuxMCOut_n4 ;
    wire MuxRound_n19 ;
    wire MuxRound_n18 ;
    wire MuxRound_n17 ;
    wire MuxRound_n16 ;
    wire MuxRound_n15 ;
    wire MuxRound_n14 ;
    wire MuxRound_n13 ;
    wire KeyReg_Inst_ff_SDE_0_next_state ;
    wire KeyReg_Inst_ff_SDE_1_next_state ;
    wire KeyReg_Inst_ff_SDE_2_next_state ;
    wire KeyReg_Inst_ff_SDE_3_next_state ;
    wire KeyReg_Inst_ff_SDE_4_next_state ;
    wire KeyReg_Inst_ff_SDE_5_next_state ;
    wire KeyReg_Inst_ff_SDE_6_next_state ;
    wire KeyReg_Inst_ff_SDE_7_next_state ;
    wire KeyReg_Inst_ff_SDE_8_next_state ;
    wire KeyReg_Inst_ff_SDE_9_next_state ;
    wire KeyReg_Inst_ff_SDE_10_next_state ;
    wire KeyReg_Inst_ff_SDE_11_next_state ;
    wire KeyReg_Inst_ff_SDE_12_next_state ;
    wire KeyReg_Inst_ff_SDE_13_next_state ;
    wire KeyReg_Inst_ff_SDE_14_next_state ;
    wire KeyReg_Inst_ff_SDE_15_next_state ;
    wire KeyReg_Inst_ff_SDE_16_next_state ;
    wire KeyReg_Inst_ff_SDE_17_next_state ;
    wire KeyReg_Inst_ff_SDE_18_next_state ;
    wire KeyReg_Inst_ff_SDE_19_next_state ;
    wire KeyReg_Inst_ff_SDE_20_next_state ;
    wire KeyReg_Inst_ff_SDE_21_next_state ;
    wire KeyReg_Inst_ff_SDE_22_next_state ;
    wire KeyReg_Inst_ff_SDE_23_next_state ;
    wire KeyReg_Inst_ff_SDE_24_next_state ;
    wire KeyReg_Inst_ff_SDE_25_next_state ;
    wire KeyReg_Inst_ff_SDE_26_next_state ;
    wire KeyReg_Inst_ff_SDE_27_next_state ;
    wire KeyReg_Inst_ff_SDE_28_next_state ;
    wire KeyReg_Inst_ff_SDE_29_next_state ;
    wire KeyReg_Inst_ff_SDE_30_next_state ;
    wire KeyReg_Inst_ff_SDE_31_next_state ;
    wire KeyReg_Inst_ff_SDE_32_next_state ;
    wire KeyReg_Inst_ff_SDE_33_next_state ;
    wire KeyReg_Inst_ff_SDE_34_next_state ;
    wire KeyReg_Inst_ff_SDE_35_next_state ;
    wire KeyReg_Inst_ff_SDE_36_next_state ;
    wire KeyReg_Inst_ff_SDE_37_next_state ;
    wire KeyReg_Inst_ff_SDE_38_next_state ;
    wire KeyReg_Inst_ff_SDE_39_next_state ;
    wire KeyReg_Inst_ff_SDE_40_next_state ;
    wire KeyReg_Inst_ff_SDE_41_next_state ;
    wire KeyReg_Inst_ff_SDE_42_next_state ;
    wire KeyReg_Inst_ff_SDE_43_next_state ;
    wire KeyReg_Inst_ff_SDE_44_next_state ;
    wire KeyReg_Inst_ff_SDE_45_next_state ;
    wire KeyReg_Inst_ff_SDE_46_next_state ;
    wire KeyReg_Inst_ff_SDE_47_next_state ;
    wire KeyReg_Inst_ff_SDE_48_next_state ;
    wire KeyReg_Inst_ff_SDE_49_next_state ;
    wire KeyReg_Inst_ff_SDE_50_next_state ;
    wire KeyReg_Inst_ff_SDE_51_next_state ;
    wire KeyReg_Inst_ff_SDE_52_next_state ;
    wire KeyReg_Inst_ff_SDE_53_next_state ;
    wire KeyReg_Inst_ff_SDE_54_next_state ;
    wire KeyReg_Inst_ff_SDE_55_next_state ;
    wire KeyReg_Inst_ff_SDE_56_next_state ;
    wire KeyReg_Inst_ff_SDE_57_next_state ;
    wire KeyReg_Inst_ff_SDE_58_next_state ;
    wire KeyReg_Inst_ff_SDE_59_next_state ;
    wire KeyReg_Inst_ff_SDE_60_next_state ;
    wire KeyReg_Inst_ff_SDE_61_next_state ;
    wire KeyReg_Inst_ff_SDE_62_next_state ;
    wire KeyReg_Inst_ff_SDE_63_next_state ;
    wire KeyReg_Inst_ff_SDE_64_next_state ;
    wire KeyReg_Inst_ff_SDE_65_next_state ;
    wire KeyReg_Inst_ff_SDE_66_next_state ;
    wire KeyReg_Inst_ff_SDE_67_next_state ;
    wire KeyReg_Inst_ff_SDE_68_next_state ;
    wire KeyReg_Inst_ff_SDE_69_next_state ;
    wire KeyReg_Inst_ff_SDE_70_next_state ;
    wire KeyReg_Inst_ff_SDE_71_next_state ;
    wire KeyReg_Inst_ff_SDE_72_next_state ;
    wire KeyReg_Inst_ff_SDE_73_next_state ;
    wire KeyReg_Inst_ff_SDE_74_next_state ;
    wire KeyReg_Inst_ff_SDE_75_next_state ;
    wire KeyReg_Inst_ff_SDE_76_next_state ;
    wire KeyReg_Inst_ff_SDE_77_next_state ;
    wire KeyReg_Inst_ff_SDE_78_next_state ;
    wire KeyReg_Inst_ff_SDE_79_next_state ;
    wire KeyReg_Inst_ff_SDE_80_next_state ;
    wire KeyReg_Inst_ff_SDE_81_next_state ;
    wire KeyReg_Inst_ff_SDE_82_next_state ;
    wire KeyReg_Inst_ff_SDE_83_next_state ;
    wire KeyReg_Inst_ff_SDE_84_next_state ;
    wire KeyReg_Inst_ff_SDE_85_next_state ;
    wire KeyReg_Inst_ff_SDE_86_next_state ;
    wire KeyReg_Inst_ff_SDE_87_next_state ;
    wire KeyReg_Inst_ff_SDE_88_next_state ;
    wire KeyReg_Inst_ff_SDE_89_next_state ;
    wire KeyReg_Inst_ff_SDE_90_next_state ;
    wire KeyReg_Inst_ff_SDE_91_next_state ;
    wire KeyReg_Inst_ff_SDE_92_next_state ;
    wire KeyReg_Inst_ff_SDE_93_next_state ;
    wire KeyReg_Inst_ff_SDE_94_next_state ;
    wire KeyReg_Inst_ff_SDE_95_next_state ;
    wire KeyReg_Inst_ff_SDE_96_next_state ;
    wire KeyReg_Inst_ff_SDE_97_next_state ;
    wire KeyReg_Inst_ff_SDE_98_next_state ;
    wire KeyReg_Inst_ff_SDE_99_next_state ;
    wire KeyReg_Inst_ff_SDE_100_next_state ;
    wire KeyReg_Inst_ff_SDE_101_next_state ;
    wire KeyReg_Inst_ff_SDE_102_next_state ;
    wire KeyReg_Inst_ff_SDE_103_next_state ;
    wire KeyReg_Inst_ff_SDE_104_next_state ;
    wire KeyReg_Inst_ff_SDE_105_next_state ;
    wire KeyReg_Inst_ff_SDE_106_next_state ;
    wire KeyReg_Inst_ff_SDE_107_next_state ;
    wire KeyReg_Inst_ff_SDE_108_next_state ;
    wire KeyReg_Inst_ff_SDE_109_next_state ;
    wire KeyReg_Inst_ff_SDE_110_next_state ;
    wire KeyReg_Inst_ff_SDE_111_next_state ;
    wire KeyReg_Inst_ff_SDE_112_next_state ;
    wire KeyReg_Inst_ff_SDE_113_next_state ;
    wire KeyReg_Inst_ff_SDE_114_next_state ;
    wire KeyReg_Inst_ff_SDE_115_next_state ;
    wire KeyReg_Inst_ff_SDE_116_next_state ;
    wire KeyReg_Inst_ff_SDE_117_next_state ;
    wire KeyReg_Inst_ff_SDE_118_next_state ;
    wire KeyReg_Inst_ff_SDE_119_next_state ;
    wire KeyReg_Inst_ff_SDE_120_next_state ;
    wire KeyReg_Inst_ff_SDE_121_next_state ;
    wire KeyReg_Inst_ff_SDE_122_next_state ;
    wire KeyReg_Inst_ff_SDE_123_next_state ;
    wire KeyReg_Inst_ff_SDE_124_next_state ;
    wire KeyReg_Inst_ff_SDE_125_next_state ;
    wire KeyReg_Inst_ff_SDE_126_next_state ;
    wire KeyReg_Inst_ff_SDE_127_next_state ;
    wire MuxKeyExpansion_n21 ;
    wire MuxKeyExpansion_n20 ;
    wire MuxKeyExpansion_n19 ;
    wire MuxKeyExpansion_n18 ;
    wire MuxKeyExpansion_n17 ;
    wire MuxKeyExpansion_n16 ;
    wire MuxKeyExpansion_n15 ;
    wire MuxKeyExpansion_n14 ;
    wire RoundCounterIns_n10 ;
    wire RoundCounterIns_n9 ;
    wire RoundCounterIns_n8 ;
    wire RoundCounterIns_n7 ;
    wire RoundCounterIns_n6 ;
    wire RoundCounterIns_n5 ;
    wire RoundCounterIns_n4 ;
    wire RoundCounterIns_n42 ;
    wire RoundCounterIns_n1 ;
    wire RoundCounterIns_n2 ;
    wire RoundCounterIns_n44 ;
    wire RoundCounterIns_n45 ;
    wire InRoundCounterIns_n12 ;
    wire InRoundCounterIns_n11 ;
    wire InRoundCounterIns_n10 ;
    wire InRoundCounterIns_n9 ;
    wire InRoundCounterIns_n8 ;
    wire InRoundCounterIns_n7 ;
    wire InRoundCounterIns_n5 ;
    wire InRoundCounterIns_n4 ;
    wire InRoundCounterIns_n3 ;
    wire InRoundCounterIns_n2 ;
    wire InRoundCounterIns_n1 ;
    wire InRoundCounterIns_n6 ;
    wire InRoundCounterIns_n39 ;
    wire InRoundCounterIns_n40 ;
    wire InRoundCounterIns_n41 ;
    wire [127:0] RoundOutput ;
    wire [127:0] ShiftRowsOutput ;
    wire [31:0] KSSubBytesInput ;
    wire [31:0] SubBytesInput ;
    wire [3:0] SubBytesOutput ;
    wire [31:0] MixColumnsOutput ;
    wire [31:0] ColumnOutput ;
    wire [127:0] RoundKeyOutput ;
    wire [127:32] RoundKey ;
    wire [7:0] Rcon ;
    wire [127:0] KeyExpansionOutput ;
    wire [3:0] RoundCounter ;
    wire [2:0] InRoundCounter ;
    wire [28:0] MixColumnsIns_DoubleBytes ;
    wire [31:0] KeyExpansionIns_tmp ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8099 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8105 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8111 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8117 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8119 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8121 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8123 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8125 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8127 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8129 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8131 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8133 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8135 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8137 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8139 ;
    wire new_AGEMA_signal_8143 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8145 ;
    wire new_AGEMA_signal_8149 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8151 ;
    wire new_AGEMA_signal_8155 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8157 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8203 ;
    wire new_AGEMA_signal_8204 ;
    wire new_AGEMA_signal_8205 ;
    wire new_AGEMA_signal_8209 ;
    wire new_AGEMA_signal_8210 ;
    wire new_AGEMA_signal_8211 ;
    wire new_AGEMA_signal_8215 ;
    wire new_AGEMA_signal_8216 ;
    wire new_AGEMA_signal_8217 ;
    wire new_AGEMA_signal_8221 ;
    wire new_AGEMA_signal_8222 ;
    wire new_AGEMA_signal_8223 ;
    wire new_AGEMA_signal_8227 ;
    wire new_AGEMA_signal_8228 ;
    wire new_AGEMA_signal_8229 ;
    wire new_AGEMA_signal_8233 ;
    wire new_AGEMA_signal_8234 ;
    wire new_AGEMA_signal_8235 ;
    wire new_AGEMA_signal_8239 ;
    wire new_AGEMA_signal_8240 ;
    wire new_AGEMA_signal_8241 ;
    wire new_AGEMA_signal_8245 ;
    wire new_AGEMA_signal_8246 ;
    wire new_AGEMA_signal_8247 ;
    wire new_AGEMA_signal_8251 ;
    wire new_AGEMA_signal_8252 ;
    wire new_AGEMA_signal_8253 ;
    wire new_AGEMA_signal_9886 ;
    wire new_AGEMA_signal_9887 ;
    wire new_AGEMA_signal_9888 ;
    wire new_AGEMA_signal_9889 ;
    wire new_AGEMA_signal_9890 ;
    wire new_AGEMA_signal_9891 ;
    wire new_AGEMA_signal_9892 ;
    wire new_AGEMA_signal_9893 ;
    wire new_AGEMA_signal_9894 ;
    wire new_AGEMA_signal_9895 ;
    wire new_AGEMA_signal_9896 ;
    wire new_AGEMA_signal_9897 ;
    wire new_AGEMA_signal_9898 ;
    wire new_AGEMA_signal_9899 ;
    wire new_AGEMA_signal_9900 ;
    wire new_AGEMA_signal_9901 ;
    wire new_AGEMA_signal_9902 ;
    wire new_AGEMA_signal_9903 ;
    wire new_AGEMA_signal_9904 ;
    wire new_AGEMA_signal_9905 ;
    wire new_AGEMA_signal_9906 ;
    wire new_AGEMA_signal_9907 ;
    wire new_AGEMA_signal_9908 ;
    wire new_AGEMA_signal_9909 ;
    wire new_AGEMA_signal_9910 ;
    wire new_AGEMA_signal_9911 ;
    wire new_AGEMA_signal_9912 ;
    wire new_AGEMA_signal_9913 ;
    wire new_AGEMA_signal_9914 ;
    wire new_AGEMA_signal_9915 ;
    wire new_AGEMA_signal_9916 ;
    wire new_AGEMA_signal_9917 ;
    wire new_AGEMA_signal_9918 ;
    wire new_AGEMA_signal_9919 ;
    wire new_AGEMA_signal_9920 ;
    wire new_AGEMA_signal_9921 ;
    wire new_AGEMA_signal_9922 ;
    wire new_AGEMA_signal_9923 ;
    wire new_AGEMA_signal_9924 ;
    wire new_AGEMA_signal_9925 ;
    wire new_AGEMA_signal_9926 ;
    wire new_AGEMA_signal_9927 ;
    wire new_AGEMA_signal_9928 ;
    wire new_AGEMA_signal_9929 ;
    wire new_AGEMA_signal_9930 ;
    wire new_AGEMA_signal_9931 ;
    wire new_AGEMA_signal_9932 ;
    wire new_AGEMA_signal_9933 ;
    wire new_AGEMA_signal_9934 ;
    wire new_AGEMA_signal_9935 ;
    wire new_AGEMA_signal_9936 ;
    wire new_AGEMA_signal_9937 ;
    wire new_AGEMA_signal_9938 ;
    wire new_AGEMA_signal_9939 ;
    wire new_AGEMA_signal_9940 ;
    wire new_AGEMA_signal_9941 ;
    wire new_AGEMA_signal_9942 ;
    wire new_AGEMA_signal_9943 ;
    wire new_AGEMA_signal_9944 ;
    wire new_AGEMA_signal_9945 ;
    wire new_AGEMA_signal_9946 ;
    wire new_AGEMA_signal_9947 ;
    wire new_AGEMA_signal_9948 ;
    wire new_AGEMA_signal_9949 ;
    wire new_AGEMA_signal_9950 ;
    wire new_AGEMA_signal_9951 ;
    wire new_AGEMA_signal_9952 ;
    wire new_AGEMA_signal_9953 ;
    wire new_AGEMA_signal_9954 ;
    wire new_AGEMA_signal_9955 ;
    wire new_AGEMA_signal_9956 ;
    wire new_AGEMA_signal_9957 ;
    wire new_AGEMA_signal_9958 ;
    wire new_AGEMA_signal_9959 ;
    wire new_AGEMA_signal_9960 ;
    wire new_AGEMA_signal_9961 ;
    wire new_AGEMA_signal_9962 ;
    wire new_AGEMA_signal_9963 ;
    wire new_AGEMA_signal_9964 ;
    wire new_AGEMA_signal_9965 ;
    wire new_AGEMA_signal_9966 ;
    wire new_AGEMA_signal_9967 ;
    wire new_AGEMA_signal_9968 ;
    wire new_AGEMA_signal_9969 ;
    wire new_AGEMA_signal_9970 ;
    wire new_AGEMA_signal_9971 ;
    wire new_AGEMA_signal_9972 ;
    wire new_AGEMA_signal_9973 ;
    wire new_AGEMA_signal_9974 ;
    wire new_AGEMA_signal_9975 ;
    wire new_AGEMA_signal_9976 ;
    wire new_AGEMA_signal_9977 ;
    wire new_AGEMA_signal_9978 ;
    wire new_AGEMA_signal_9979 ;
    wire new_AGEMA_signal_9980 ;
    wire new_AGEMA_signal_9981 ;
    wire new_AGEMA_signal_9982 ;
    wire new_AGEMA_signal_9983 ;
    wire new_AGEMA_signal_9984 ;
    wire new_AGEMA_signal_9985 ;
    wire new_AGEMA_signal_9986 ;
    wire new_AGEMA_signal_9987 ;
    wire new_AGEMA_signal_9988 ;
    wire new_AGEMA_signal_9989 ;
    wire new_AGEMA_signal_9990 ;
    wire new_AGEMA_signal_9991 ;
    wire new_AGEMA_signal_9992 ;
    wire new_AGEMA_signal_9993 ;
    wire new_AGEMA_signal_9994 ;
    wire new_AGEMA_signal_9995 ;
    wire new_AGEMA_signal_9996 ;
    wire new_AGEMA_signal_9997 ;
    wire new_AGEMA_signal_9998 ;
    wire new_AGEMA_signal_9999 ;
    wire new_AGEMA_signal_10000 ;
    wire new_AGEMA_signal_10001 ;
    wire new_AGEMA_signal_10002 ;
    wire new_AGEMA_signal_10003 ;
    wire new_AGEMA_signal_10004 ;
    wire new_AGEMA_signal_10005 ;
    wire new_AGEMA_signal_10006 ;
    wire new_AGEMA_signal_10007 ;
    wire new_AGEMA_signal_10008 ;
    wire new_AGEMA_signal_10009 ;
    wire new_AGEMA_signal_10010 ;
    wire new_AGEMA_signal_10011 ;
    wire new_AGEMA_signal_10012 ;
    wire new_AGEMA_signal_10013 ;
    wire new_AGEMA_signal_10014 ;
    wire new_AGEMA_signal_10015 ;
    wire new_AGEMA_signal_10016 ;
    wire new_AGEMA_signal_10017 ;
    wire new_AGEMA_signal_10018 ;
    wire new_AGEMA_signal_10019 ;
    wire new_AGEMA_signal_10020 ;
    wire new_AGEMA_signal_10021 ;
    wire new_AGEMA_signal_10022 ;
    wire new_AGEMA_signal_10023 ;
    wire new_AGEMA_signal_10024 ;
    wire new_AGEMA_signal_10025 ;
    wire new_AGEMA_signal_10026 ;
    wire new_AGEMA_signal_10027 ;
    wire new_AGEMA_signal_10028 ;
    wire new_AGEMA_signal_10029 ;
    wire new_AGEMA_signal_10030 ;
    wire new_AGEMA_signal_10031 ;
    wire new_AGEMA_signal_10032 ;
    wire new_AGEMA_signal_10033 ;
    wire new_AGEMA_signal_10034 ;
    wire new_AGEMA_signal_10035 ;
    wire new_AGEMA_signal_10036 ;
    wire new_AGEMA_signal_10037 ;
    wire new_AGEMA_signal_10038 ;
    wire new_AGEMA_signal_10039 ;
    wire new_AGEMA_signal_10040 ;
    wire new_AGEMA_signal_10041 ;
    wire new_AGEMA_signal_10042 ;
    wire new_AGEMA_signal_10043 ;
    wire new_AGEMA_signal_10044 ;
    wire new_AGEMA_signal_10045 ;
    wire new_AGEMA_signal_10046 ;
    wire new_AGEMA_signal_10047 ;
    wire new_AGEMA_signal_10048 ;
    wire new_AGEMA_signal_10049 ;
    wire new_AGEMA_signal_10050 ;
    wire new_AGEMA_signal_10051 ;
    wire new_AGEMA_signal_10052 ;
    wire new_AGEMA_signal_10053 ;
    wire new_AGEMA_signal_10054 ;
    wire new_AGEMA_signal_10055 ;
    wire new_AGEMA_signal_10056 ;
    wire new_AGEMA_signal_10057 ;
    wire new_AGEMA_signal_10058 ;
    wire new_AGEMA_signal_10059 ;
    wire new_AGEMA_signal_10060 ;
    wire new_AGEMA_signal_10061 ;
    wire new_AGEMA_signal_10062 ;
    wire new_AGEMA_signal_10063 ;
    wire new_AGEMA_signal_10064 ;
    wire new_AGEMA_signal_10065 ;
    wire new_AGEMA_signal_10066 ;
    wire new_AGEMA_signal_10067 ;
    wire new_AGEMA_signal_10068 ;
    wire new_AGEMA_signal_10069 ;
    wire new_AGEMA_signal_10070 ;
    wire new_AGEMA_signal_10071 ;
    wire new_AGEMA_signal_10072 ;
    wire new_AGEMA_signal_10073 ;
    wire new_AGEMA_signal_10074 ;
    wire new_AGEMA_signal_10075 ;
    wire new_AGEMA_signal_10076 ;
    wire new_AGEMA_signal_10077 ;
    wire new_AGEMA_signal_10078 ;
    wire new_AGEMA_signal_10079 ;
    wire new_AGEMA_signal_10080 ;
    wire new_AGEMA_signal_10081 ;
    wire new_AGEMA_signal_10082 ;
    wire new_AGEMA_signal_10083 ;
    wire new_AGEMA_signal_10084 ;
    wire new_AGEMA_signal_10085 ;
    wire new_AGEMA_signal_10086 ;
    wire new_AGEMA_signal_10087 ;
    wire new_AGEMA_signal_10088 ;
    wire new_AGEMA_signal_10089 ;
    wire new_AGEMA_signal_10090 ;
    wire new_AGEMA_signal_10091 ;
    wire new_AGEMA_signal_10092 ;
    wire new_AGEMA_signal_10093 ;
    wire new_AGEMA_signal_10094 ;
    wire new_AGEMA_signal_10095 ;
    wire new_AGEMA_signal_10096 ;
    wire new_AGEMA_signal_10097 ;
    wire new_AGEMA_signal_10098 ;
    wire new_AGEMA_signal_10099 ;
    wire new_AGEMA_signal_10100 ;
    wire new_AGEMA_signal_10101 ;
    wire new_AGEMA_signal_10102 ;
    wire new_AGEMA_signal_10103 ;
    wire new_AGEMA_signal_10104 ;
    wire new_AGEMA_signal_10105 ;
    wire new_AGEMA_signal_10106 ;
    wire new_AGEMA_signal_10107 ;
    wire new_AGEMA_signal_10108 ;
    wire new_AGEMA_signal_10109 ;
    wire new_AGEMA_signal_10110 ;
    wire new_AGEMA_signal_10111 ;
    wire new_AGEMA_signal_10112 ;
    wire new_AGEMA_signal_10113 ;
    wire new_AGEMA_signal_10114 ;
    wire new_AGEMA_signal_10115 ;
    wire new_AGEMA_signal_10116 ;
    wire new_AGEMA_signal_10117 ;
    wire new_AGEMA_signal_10118 ;
    wire new_AGEMA_signal_10119 ;
    wire new_AGEMA_signal_10120 ;
    wire new_AGEMA_signal_10121 ;
    wire new_AGEMA_signal_10122 ;
    wire new_AGEMA_signal_10123 ;
    wire new_AGEMA_signal_10124 ;
    wire new_AGEMA_signal_10125 ;
    wire new_AGEMA_signal_10126 ;
    wire new_AGEMA_signal_10127 ;
    wire new_AGEMA_signal_10128 ;
    wire new_AGEMA_signal_10129 ;
    wire new_AGEMA_signal_10130 ;
    wire new_AGEMA_signal_10131 ;
    wire new_AGEMA_signal_10132 ;
    wire new_AGEMA_signal_10133 ;
    wire new_AGEMA_signal_10134 ;
    wire new_AGEMA_signal_10135 ;
    wire new_AGEMA_signal_10136 ;
    wire new_AGEMA_signal_10137 ;
    wire new_AGEMA_signal_10138 ;
    wire new_AGEMA_signal_10139 ;
    wire new_AGEMA_signal_10140 ;
    wire new_AGEMA_signal_10141 ;
    wire new_AGEMA_signal_10142 ;
    wire new_AGEMA_signal_10143 ;
    wire new_AGEMA_signal_10144 ;
    wire new_AGEMA_signal_10145 ;
    wire new_AGEMA_signal_10146 ;
    wire new_AGEMA_signal_10147 ;
    wire new_AGEMA_signal_10148 ;
    wire new_AGEMA_signal_10149 ;
    wire new_AGEMA_signal_10150 ;
    wire new_AGEMA_signal_10151 ;
    wire new_AGEMA_signal_10152 ;
    wire new_AGEMA_signal_10153 ;
    wire new_AGEMA_signal_10154 ;
    wire new_AGEMA_signal_10155 ;
    wire new_AGEMA_signal_10156 ;
    wire new_AGEMA_signal_10157 ;
    wire new_AGEMA_signal_10158 ;
    wire new_AGEMA_signal_10159 ;
    wire new_AGEMA_signal_10160 ;
    wire new_AGEMA_signal_10161 ;
    wire new_AGEMA_signal_10162 ;
    wire new_AGEMA_signal_10163 ;
    wire new_AGEMA_signal_10164 ;
    wire new_AGEMA_signal_10165 ;
    wire new_AGEMA_signal_10166 ;
    wire new_AGEMA_signal_10167 ;
    wire new_AGEMA_signal_10168 ;
    wire new_AGEMA_signal_10169 ;
    wire new_AGEMA_signal_10170 ;
    wire new_AGEMA_signal_10171 ;
    wire new_AGEMA_signal_10172 ;
    wire new_AGEMA_signal_10173 ;
    wire new_AGEMA_signal_10174 ;
    wire new_AGEMA_signal_10175 ;
    wire new_AGEMA_signal_10176 ;
    wire new_AGEMA_signal_10177 ;
    wire new_AGEMA_signal_10178 ;
    wire new_AGEMA_signal_10179 ;
    wire new_AGEMA_signal_10180 ;
    wire new_AGEMA_signal_10181 ;
    wire new_AGEMA_signal_10182 ;
    wire new_AGEMA_signal_10183 ;
    wire new_AGEMA_signal_10184 ;
    wire new_AGEMA_signal_10185 ;
    wire new_AGEMA_signal_10186 ;
    wire new_AGEMA_signal_10187 ;
    wire new_AGEMA_signal_10188 ;
    wire new_AGEMA_signal_10189 ;
    wire new_AGEMA_signal_10190 ;
    wire new_AGEMA_signal_10191 ;
    wire new_AGEMA_signal_10192 ;
    wire new_AGEMA_signal_10193 ;
    wire new_AGEMA_signal_10194 ;
    wire new_AGEMA_signal_10195 ;
    wire new_AGEMA_signal_10196 ;
    wire new_AGEMA_signal_10197 ;
    wire new_AGEMA_signal_10198 ;
    wire new_AGEMA_signal_10199 ;
    wire new_AGEMA_signal_10200 ;
    wire new_AGEMA_signal_10201 ;
    wire new_AGEMA_signal_10202 ;
    wire new_AGEMA_signal_10203 ;
    wire new_AGEMA_signal_10204 ;
    wire new_AGEMA_signal_10205 ;
    wire new_AGEMA_signal_10206 ;
    wire new_AGEMA_signal_10207 ;
    wire new_AGEMA_signal_10208 ;
    wire new_AGEMA_signal_10209 ;
    wire new_AGEMA_signal_10210 ;
    wire new_AGEMA_signal_10211 ;
    wire new_AGEMA_signal_10212 ;
    wire new_AGEMA_signal_10213 ;
    wire new_AGEMA_signal_10214 ;
    wire new_AGEMA_signal_10215 ;
    wire new_AGEMA_signal_10216 ;
    wire new_AGEMA_signal_10217 ;
    wire new_AGEMA_signal_10218 ;
    wire new_AGEMA_signal_10219 ;
    wire new_AGEMA_signal_10220 ;
    wire new_AGEMA_signal_10221 ;
    wire new_AGEMA_signal_10222 ;
    wire new_AGEMA_signal_10223 ;
    wire new_AGEMA_signal_10224 ;
    wire new_AGEMA_signal_10225 ;
    wire new_AGEMA_signal_10226 ;
    wire new_AGEMA_signal_10227 ;
    wire new_AGEMA_signal_10228 ;
    wire new_AGEMA_signal_10229 ;
    wire new_AGEMA_signal_10230 ;
    wire new_AGEMA_signal_10231 ;
    wire new_AGEMA_signal_10232 ;
    wire new_AGEMA_signal_10233 ;
    wire new_AGEMA_signal_10234 ;
    wire new_AGEMA_signal_10235 ;
    wire new_AGEMA_signal_10236 ;
    wire new_AGEMA_signal_10237 ;
    wire new_AGEMA_signal_10238 ;
    wire new_AGEMA_signal_10239 ;
    wire new_AGEMA_signal_10240 ;
    wire new_AGEMA_signal_10241 ;
    wire new_AGEMA_signal_10242 ;
    wire new_AGEMA_signal_10243 ;
    wire new_AGEMA_signal_10244 ;
    wire new_AGEMA_signal_10245 ;
    wire new_AGEMA_signal_10246 ;
    wire new_AGEMA_signal_10247 ;
    wire new_AGEMA_signal_10248 ;
    wire new_AGEMA_signal_10249 ;
    wire new_AGEMA_signal_10250 ;
    wire new_AGEMA_signal_10251 ;
    wire new_AGEMA_signal_10252 ;
    wire new_AGEMA_signal_10253 ;
    wire new_AGEMA_signal_10254 ;
    wire new_AGEMA_signal_10255 ;
    wire new_AGEMA_signal_10256 ;
    wire new_AGEMA_signal_10257 ;
    wire new_AGEMA_signal_10258 ;
    wire new_AGEMA_signal_10259 ;
    wire new_AGEMA_signal_10260 ;
    wire new_AGEMA_signal_10261 ;
    wire new_AGEMA_signal_10262 ;
    wire new_AGEMA_signal_10263 ;
    wire new_AGEMA_signal_10264 ;
    wire new_AGEMA_signal_10265 ;
    wire new_AGEMA_signal_10266 ;
    wire new_AGEMA_signal_10267 ;
    wire new_AGEMA_signal_10268 ;
    wire new_AGEMA_signal_10269 ;
    wire new_AGEMA_signal_10270 ;
    wire new_AGEMA_signal_10271 ;
    wire new_AGEMA_signal_10272 ;
    wire new_AGEMA_signal_10273 ;
    wire new_AGEMA_signal_10274 ;
    wire new_AGEMA_signal_10275 ;
    wire new_AGEMA_signal_10276 ;
    wire new_AGEMA_signal_10277 ;
    wire new_AGEMA_signal_10278 ;
    wire new_AGEMA_signal_10279 ;
    wire new_AGEMA_signal_10280 ;
    wire new_AGEMA_signal_10281 ;
    wire new_AGEMA_signal_10282 ;
    wire new_AGEMA_signal_10283 ;
    wire new_AGEMA_signal_10284 ;
    wire new_AGEMA_signal_10285 ;
    wire new_AGEMA_signal_10286 ;
    wire new_AGEMA_signal_10287 ;
    wire new_AGEMA_signal_10288 ;
    wire new_AGEMA_signal_10289 ;
    wire new_AGEMA_signal_10290 ;
    wire new_AGEMA_signal_10291 ;
    wire new_AGEMA_signal_10292 ;
    wire new_AGEMA_signal_10293 ;
    wire new_AGEMA_signal_10294 ;
    wire new_AGEMA_signal_10295 ;
    wire new_AGEMA_signal_10296 ;
    wire new_AGEMA_signal_10297 ;
    wire new_AGEMA_signal_10298 ;
    wire new_AGEMA_signal_10299 ;
    wire new_AGEMA_signal_10300 ;
    wire new_AGEMA_signal_10301 ;
    wire new_AGEMA_signal_10302 ;
    wire new_AGEMA_signal_10303 ;
    wire new_AGEMA_signal_10304 ;
    wire new_AGEMA_signal_10305 ;
    wire new_AGEMA_signal_10306 ;
    wire new_AGEMA_signal_10307 ;
    wire new_AGEMA_signal_10308 ;
    wire new_AGEMA_signal_10309 ;
    wire new_AGEMA_signal_10310 ;
    wire new_AGEMA_signal_10311 ;
    wire new_AGEMA_signal_10312 ;
    wire new_AGEMA_signal_10313 ;
    wire new_AGEMA_signal_10314 ;
    wire new_AGEMA_signal_10315 ;
    wire new_AGEMA_signal_10316 ;
    wire new_AGEMA_signal_10317 ;
    wire new_AGEMA_signal_10318 ;
    wire new_AGEMA_signal_10319 ;
    wire new_AGEMA_signal_10320 ;
    wire new_AGEMA_signal_10321 ;
    wire new_AGEMA_signal_10322 ;
    wire new_AGEMA_signal_10323 ;
    wire new_AGEMA_signal_10324 ;
    wire new_AGEMA_signal_10325 ;
    wire new_AGEMA_signal_10326 ;
    wire new_AGEMA_signal_10327 ;
    wire new_AGEMA_signal_10328 ;
    wire new_AGEMA_signal_10329 ;
    wire new_AGEMA_signal_10330 ;
    wire new_AGEMA_signal_10331 ;
    wire new_AGEMA_signal_10332 ;
    wire new_AGEMA_signal_10333 ;
    wire new_AGEMA_signal_10334 ;
    wire new_AGEMA_signal_10335 ;
    wire new_AGEMA_signal_10336 ;
    wire new_AGEMA_signal_10337 ;
    wire new_AGEMA_signal_10338 ;
    wire new_AGEMA_signal_10339 ;
    wire new_AGEMA_signal_10340 ;
    wire new_AGEMA_signal_10341 ;
    wire new_AGEMA_signal_10342 ;
    wire new_AGEMA_signal_10343 ;
    wire new_AGEMA_signal_10344 ;
    wire new_AGEMA_signal_10345 ;
    wire new_AGEMA_signal_10346 ;
    wire new_AGEMA_signal_10347 ;
    wire new_AGEMA_signal_10348 ;
    wire new_AGEMA_signal_10349 ;
    wire new_AGEMA_signal_10350 ;
    wire new_AGEMA_signal_10351 ;
    wire new_AGEMA_signal_10352 ;
    wire new_AGEMA_signal_10353 ;
    wire new_AGEMA_signal_10354 ;
    wire new_AGEMA_signal_10355 ;
    wire new_AGEMA_signal_10356 ;
    wire new_AGEMA_signal_10357 ;
    wire new_AGEMA_signal_10358 ;
    wire new_AGEMA_signal_10359 ;
    wire new_AGEMA_signal_10360 ;
    wire new_AGEMA_signal_10361 ;
    wire new_AGEMA_signal_10362 ;
    wire new_AGEMA_signal_10363 ;
    wire new_AGEMA_signal_10364 ;
    wire new_AGEMA_signal_10365 ;
    wire new_AGEMA_signal_10366 ;
    wire new_AGEMA_signal_10367 ;
    wire new_AGEMA_signal_10368 ;
    wire new_AGEMA_signal_10369 ;
    wire new_AGEMA_signal_10370 ;
    wire new_AGEMA_signal_10371 ;
    wire new_AGEMA_signal_10372 ;
    wire new_AGEMA_signal_10373 ;
    wire new_AGEMA_signal_10374 ;
    wire new_AGEMA_signal_10375 ;
    wire new_AGEMA_signal_10376 ;
    wire new_AGEMA_signal_10377 ;
    wire new_AGEMA_signal_10378 ;
    wire new_AGEMA_signal_10379 ;
    wire new_AGEMA_signal_10380 ;
    wire new_AGEMA_signal_10381 ;
    wire new_AGEMA_signal_10382 ;
    wire new_AGEMA_signal_10383 ;
    wire new_AGEMA_signal_10384 ;
    wire new_AGEMA_signal_10385 ;
    wire new_AGEMA_signal_10386 ;
    wire new_AGEMA_signal_10387 ;
    wire new_AGEMA_signal_10388 ;
    wire new_AGEMA_signal_10389 ;
    wire new_AGEMA_signal_10390 ;
    wire new_AGEMA_signal_10391 ;
    wire new_AGEMA_signal_10392 ;
    wire new_AGEMA_signal_10393 ;
    wire new_AGEMA_signal_10394 ;
    wire new_AGEMA_signal_10395 ;
    wire new_AGEMA_signal_10396 ;
    wire new_AGEMA_signal_10397 ;
    wire new_AGEMA_signal_10398 ;
    wire new_AGEMA_signal_10399 ;
    wire new_AGEMA_signal_10400 ;
    wire new_AGEMA_signal_10401 ;
    wire new_AGEMA_signal_10402 ;
    wire new_AGEMA_signal_10403 ;
    wire new_AGEMA_signal_10404 ;
    wire new_AGEMA_signal_10405 ;
    wire new_AGEMA_signal_10406 ;
    wire new_AGEMA_signal_10407 ;
    wire new_AGEMA_signal_10408 ;
    wire new_AGEMA_signal_10409 ;
    wire new_AGEMA_signal_10410 ;
    wire new_AGEMA_signal_10411 ;
    wire new_AGEMA_signal_10412 ;
    wire new_AGEMA_signal_10413 ;
    wire new_AGEMA_signal_10414 ;
    wire new_AGEMA_signal_10415 ;
    wire new_AGEMA_signal_10416 ;
    wire new_AGEMA_signal_10417 ;
    wire new_AGEMA_signal_10418 ;
    wire new_AGEMA_signal_10419 ;
    wire new_AGEMA_signal_10420 ;
    wire new_AGEMA_signal_10421 ;
    wire new_AGEMA_signal_10422 ;
    wire new_AGEMA_signal_10423 ;
    wire new_AGEMA_signal_10424 ;
    wire new_AGEMA_signal_10425 ;
    wire new_AGEMA_signal_10426 ;
    wire new_AGEMA_signal_10427 ;
    wire new_AGEMA_signal_10428 ;
    wire new_AGEMA_signal_10429 ;
    wire new_AGEMA_signal_10430 ;
    wire new_AGEMA_signal_10431 ;
    wire new_AGEMA_signal_10432 ;
    wire new_AGEMA_signal_10433 ;
    wire new_AGEMA_signal_10434 ;
    wire new_AGEMA_signal_10435 ;
    wire new_AGEMA_signal_10436 ;
    wire new_AGEMA_signal_10437 ;
    wire new_AGEMA_signal_10438 ;
    wire new_AGEMA_signal_10439 ;
    wire new_AGEMA_signal_10440 ;
    wire new_AGEMA_signal_10441 ;
    wire new_AGEMA_signal_10442 ;
    wire new_AGEMA_signal_10443 ;
    wire new_AGEMA_signal_10444 ;
    wire new_AGEMA_signal_10445 ;
    wire new_AGEMA_signal_10446 ;
    wire new_AGEMA_signal_10447 ;
    wire new_AGEMA_signal_10448 ;
    wire new_AGEMA_signal_10449 ;
    wire new_AGEMA_signal_10450 ;
    wire new_AGEMA_signal_10451 ;
    wire new_AGEMA_signal_10452 ;
    wire new_AGEMA_signal_10453 ;
    wire new_AGEMA_signal_10454 ;
    wire new_AGEMA_signal_10455 ;
    wire new_AGEMA_signal_10456 ;
    wire new_AGEMA_signal_10457 ;
    wire new_AGEMA_signal_10458 ;
    wire new_AGEMA_signal_10459 ;
    wire new_AGEMA_signal_10460 ;
    wire new_AGEMA_signal_10461 ;
    wire new_AGEMA_signal_10462 ;
    wire new_AGEMA_signal_10463 ;
    wire new_AGEMA_signal_10464 ;
    wire new_AGEMA_signal_10465 ;
    wire new_AGEMA_signal_10466 ;
    wire new_AGEMA_signal_10467 ;
    wire new_AGEMA_signal_10468 ;
    wire new_AGEMA_signal_10469 ;
    wire new_AGEMA_signal_10470 ;
    wire new_AGEMA_signal_10471 ;
    wire new_AGEMA_signal_10472 ;
    wire new_AGEMA_signal_10473 ;
    wire new_AGEMA_signal_10474 ;
    wire new_AGEMA_signal_10475 ;
    wire new_AGEMA_signal_10476 ;
    wire new_AGEMA_signal_10477 ;
    wire new_AGEMA_signal_10478 ;
    wire new_AGEMA_signal_10479 ;
    wire new_AGEMA_signal_10480 ;
    wire new_AGEMA_signal_10481 ;
    wire new_AGEMA_signal_10482 ;
    wire new_AGEMA_signal_10483 ;
    wire new_AGEMA_signal_10484 ;
    wire new_AGEMA_signal_10485 ;
    wire new_AGEMA_signal_10486 ;
    wire new_AGEMA_signal_10487 ;
    wire new_AGEMA_signal_10488 ;
    wire new_AGEMA_signal_10489 ;
    wire new_AGEMA_signal_10490 ;
    wire new_AGEMA_signal_10491 ;
    wire new_AGEMA_signal_10492 ;
    wire new_AGEMA_signal_10493 ;
    wire new_AGEMA_signal_10494 ;
    wire new_AGEMA_signal_10495 ;
    wire new_AGEMA_signal_10496 ;
    wire new_AGEMA_signal_10497 ;
    wire new_AGEMA_signal_10498 ;
    wire new_AGEMA_signal_10499 ;
    wire new_AGEMA_signal_10500 ;
    wire new_AGEMA_signal_10501 ;
    wire new_AGEMA_signal_10502 ;
    wire new_AGEMA_signal_10503 ;
    wire new_AGEMA_signal_10504 ;
    wire new_AGEMA_signal_10505 ;
    wire new_AGEMA_signal_10506 ;
    wire new_AGEMA_signal_10507 ;
    wire new_AGEMA_signal_10508 ;
    wire new_AGEMA_signal_10509 ;
    wire new_AGEMA_signal_10510 ;
    wire new_AGEMA_signal_10511 ;
    wire new_AGEMA_signal_10512 ;
    wire new_AGEMA_signal_10513 ;
    wire new_AGEMA_signal_10514 ;
    wire new_AGEMA_signal_10515 ;
    wire new_AGEMA_signal_10516 ;
    wire new_AGEMA_signal_10517 ;
    wire new_AGEMA_signal_10518 ;
    wire new_AGEMA_signal_10519 ;
    wire new_AGEMA_signal_10520 ;
    wire new_AGEMA_signal_10521 ;
    wire new_AGEMA_signal_10522 ;
    wire new_AGEMA_signal_10523 ;
    wire new_AGEMA_signal_10524 ;
    wire new_AGEMA_signal_10525 ;
    wire new_AGEMA_signal_10526 ;
    wire new_AGEMA_signal_10527 ;
    wire new_AGEMA_signal_10528 ;
    wire new_AGEMA_signal_10529 ;
    wire new_AGEMA_signal_10530 ;
    wire new_AGEMA_signal_10531 ;
    wire new_AGEMA_signal_10532 ;
    wire new_AGEMA_signal_10533 ;
    wire new_AGEMA_signal_10534 ;
    wire new_AGEMA_signal_10535 ;
    wire new_AGEMA_signal_10536 ;
    wire new_AGEMA_signal_10537 ;
    wire new_AGEMA_signal_10538 ;
    wire new_AGEMA_signal_10539 ;
    wire new_AGEMA_signal_10540 ;
    wire new_AGEMA_signal_10541 ;
    wire new_AGEMA_signal_10542 ;
    wire new_AGEMA_signal_10543 ;
    wire new_AGEMA_signal_10544 ;
    wire new_AGEMA_signal_10545 ;
    wire new_AGEMA_signal_10546 ;
    wire new_AGEMA_signal_10547 ;
    wire new_AGEMA_signal_10548 ;
    wire new_AGEMA_signal_10549 ;
    wire new_AGEMA_signal_10550 ;
    wire new_AGEMA_signal_10551 ;
    wire new_AGEMA_signal_10552 ;
    wire new_AGEMA_signal_10553 ;
    wire new_AGEMA_signal_10554 ;
    wire new_AGEMA_signal_10555 ;
    wire new_AGEMA_signal_10556 ;
    wire new_AGEMA_signal_10557 ;
    wire new_AGEMA_signal_10558 ;
    wire new_AGEMA_signal_10559 ;
    wire new_AGEMA_signal_10560 ;
    wire new_AGEMA_signal_10561 ;
    wire new_AGEMA_signal_10562 ;
    wire new_AGEMA_signal_10563 ;
    wire new_AGEMA_signal_10564 ;
    wire new_AGEMA_signal_10565 ;
    wire new_AGEMA_signal_10566 ;
    wire new_AGEMA_signal_10567 ;
    wire new_AGEMA_signal_10568 ;
    wire new_AGEMA_signal_10569 ;
    wire new_AGEMA_signal_10570 ;
    wire new_AGEMA_signal_10571 ;
    wire new_AGEMA_signal_10572 ;
    wire new_AGEMA_signal_10573 ;
    wire new_AGEMA_signal_10574 ;
    wire new_AGEMA_signal_10575 ;
    wire new_AGEMA_signal_10576 ;
    wire new_AGEMA_signal_10577 ;
    wire new_AGEMA_signal_10578 ;
    wire new_AGEMA_signal_10579 ;
    wire new_AGEMA_signal_10580 ;
    wire new_AGEMA_signal_10581 ;
    wire new_AGEMA_signal_10582 ;
    wire new_AGEMA_signal_10583 ;
    wire new_AGEMA_signal_10584 ;
    wire new_AGEMA_signal_10585 ;
    wire new_AGEMA_signal_10586 ;
    wire new_AGEMA_signal_10587 ;
    wire new_AGEMA_signal_10588 ;
    wire new_AGEMA_signal_10589 ;
    wire new_AGEMA_signal_10590 ;
    wire new_AGEMA_signal_10591 ;
    wire new_AGEMA_signal_10592 ;
    wire new_AGEMA_signal_10593 ;
    wire new_AGEMA_signal_10594 ;
    wire new_AGEMA_signal_10595 ;
    wire new_AGEMA_signal_10596 ;
    wire new_AGEMA_signal_10597 ;
    wire new_AGEMA_signal_10598 ;
    wire new_AGEMA_signal_10599 ;
    wire new_AGEMA_signal_10600 ;
    wire new_AGEMA_signal_10601 ;
    wire new_AGEMA_signal_10602 ;
    wire new_AGEMA_signal_10603 ;
    wire new_AGEMA_signal_10604 ;
    wire new_AGEMA_signal_10605 ;
    wire new_AGEMA_signal_10606 ;
    wire new_AGEMA_signal_10607 ;
    wire new_AGEMA_signal_10608 ;
    wire new_AGEMA_signal_10609 ;
    wire new_AGEMA_signal_10610 ;
    wire new_AGEMA_signal_10611 ;
    wire new_AGEMA_signal_10612 ;
    wire new_AGEMA_signal_10613 ;
    wire new_AGEMA_signal_10614 ;
    wire new_AGEMA_signal_10615 ;
    wire new_AGEMA_signal_10616 ;
    wire new_AGEMA_signal_10617 ;
    wire new_AGEMA_signal_10618 ;
    wire new_AGEMA_signal_10619 ;
    wire new_AGEMA_signal_10620 ;
    wire new_AGEMA_signal_10621 ;
    wire new_AGEMA_signal_10622 ;
    wire new_AGEMA_signal_10623 ;
    wire new_AGEMA_signal_10624 ;
    wire new_AGEMA_signal_10625 ;
    wire new_AGEMA_signal_10626 ;
    wire new_AGEMA_signal_10627 ;
    wire new_AGEMA_signal_10628 ;
    wire new_AGEMA_signal_10629 ;
    wire new_AGEMA_signal_10630 ;
    wire new_AGEMA_signal_10631 ;
    wire new_AGEMA_signal_10632 ;
    wire new_AGEMA_signal_10633 ;
    wire new_AGEMA_signal_10634 ;
    wire new_AGEMA_signal_10635 ;
    wire new_AGEMA_signal_10636 ;
    wire new_AGEMA_signal_10637 ;
    wire new_AGEMA_signal_10638 ;
    wire new_AGEMA_signal_10639 ;
    wire new_AGEMA_signal_10640 ;
    wire new_AGEMA_signal_10641 ;
    wire new_AGEMA_signal_10642 ;
    wire new_AGEMA_signal_10643 ;
    wire new_AGEMA_signal_10644 ;
    wire new_AGEMA_signal_10645 ;
    wire new_AGEMA_signal_10646 ;
    wire new_AGEMA_signal_10647 ;
    wire new_AGEMA_signal_10648 ;
    wire new_AGEMA_signal_10649 ;
    wire new_AGEMA_signal_10650 ;
    wire new_AGEMA_signal_10651 ;
    wire new_AGEMA_signal_10652 ;
    wire new_AGEMA_signal_10653 ;
    wire new_AGEMA_signal_10654 ;
    wire new_AGEMA_signal_10655 ;
    wire new_AGEMA_signal_10656 ;
    wire new_AGEMA_signal_10657 ;
    wire new_AGEMA_signal_10658 ;
    wire new_AGEMA_signal_10659 ;
    wire new_AGEMA_signal_10660 ;
    wire new_AGEMA_signal_10661 ;
    wire new_AGEMA_signal_10662 ;
    wire new_AGEMA_signal_10663 ;
    wire new_AGEMA_signal_10664 ;
    wire new_AGEMA_signal_10665 ;
    wire new_AGEMA_signal_10666 ;
    wire new_AGEMA_signal_10667 ;
    wire new_AGEMA_signal_10668 ;
    wire new_AGEMA_signal_10669 ;
    wire new_AGEMA_signal_10670 ;
    wire new_AGEMA_signal_10671 ;
    wire new_AGEMA_signal_10672 ;
    wire new_AGEMA_signal_10673 ;
    wire new_AGEMA_signal_10674 ;
    wire new_AGEMA_signal_10675 ;
    wire new_AGEMA_signal_10676 ;
    wire new_AGEMA_signal_10677 ;
    wire new_AGEMA_signal_10678 ;
    wire new_AGEMA_signal_10679 ;
    wire new_AGEMA_signal_10680 ;
    wire new_AGEMA_signal_10681 ;
    wire new_AGEMA_signal_10682 ;
    wire new_AGEMA_signal_10683 ;
    wire new_AGEMA_signal_10684 ;
    wire new_AGEMA_signal_10685 ;
    wire new_AGEMA_signal_10686 ;
    wire new_AGEMA_signal_10687 ;
    wire new_AGEMA_signal_10688 ;
    wire new_AGEMA_signal_10689 ;
    wire new_AGEMA_signal_10690 ;
    wire new_AGEMA_signal_10691 ;
    wire new_AGEMA_signal_10692 ;
    wire new_AGEMA_signal_10693 ;
    wire new_AGEMA_signal_10694 ;
    wire new_AGEMA_signal_10695 ;
    wire new_AGEMA_signal_10696 ;
    wire new_AGEMA_signal_10697 ;
    wire new_AGEMA_signal_10698 ;
    wire new_AGEMA_signal_10699 ;
    wire new_AGEMA_signal_10700 ;
    wire new_AGEMA_signal_10701 ;
    wire new_AGEMA_signal_10702 ;
    wire new_AGEMA_signal_10703 ;
    wire new_AGEMA_signal_10704 ;
    wire new_AGEMA_signal_10705 ;
    wire new_AGEMA_signal_10706 ;
    wire new_AGEMA_signal_10707 ;
    wire new_AGEMA_signal_10708 ;
    wire new_AGEMA_signal_10709 ;
    wire new_AGEMA_signal_10710 ;
    wire new_AGEMA_signal_10711 ;
    wire new_AGEMA_signal_10712 ;
    wire new_AGEMA_signal_10713 ;
    wire new_AGEMA_signal_10714 ;
    wire new_AGEMA_signal_10715 ;
    wire new_AGEMA_signal_10716 ;
    wire new_AGEMA_signal_10717 ;
    wire new_AGEMA_signal_10718 ;
    wire new_AGEMA_signal_10719 ;
    wire new_AGEMA_signal_10720 ;
    wire new_AGEMA_signal_10721 ;
    wire new_AGEMA_signal_10722 ;
    wire new_AGEMA_signal_10723 ;
    wire new_AGEMA_signal_10724 ;
    wire new_AGEMA_signal_10725 ;
    wire new_AGEMA_signal_10726 ;
    wire new_AGEMA_signal_10727 ;
    wire new_AGEMA_signal_10728 ;
    wire new_AGEMA_signal_10729 ;
    wire new_AGEMA_signal_10730 ;
    wire new_AGEMA_signal_10731 ;
    wire new_AGEMA_signal_10732 ;
    wire new_AGEMA_signal_10733 ;
    wire new_AGEMA_signal_10734 ;
    wire new_AGEMA_signal_10735 ;
    wire new_AGEMA_signal_10736 ;
    wire new_AGEMA_signal_10737 ;
    wire new_AGEMA_signal_10738 ;
    wire new_AGEMA_signal_10739 ;
    wire new_AGEMA_signal_10740 ;
    wire new_AGEMA_signal_10741 ;
    wire new_AGEMA_signal_10742 ;
    wire new_AGEMA_signal_10743 ;
    wire new_AGEMA_signal_10744 ;
    wire new_AGEMA_signal_10745 ;
    wire new_AGEMA_signal_10746 ;
    wire new_AGEMA_signal_10747 ;
    wire new_AGEMA_signal_10748 ;
    wire new_AGEMA_signal_10749 ;
    wire new_AGEMA_signal_10750 ;
    wire new_AGEMA_signal_10751 ;
    wire new_AGEMA_signal_10752 ;
    wire new_AGEMA_signal_10753 ;
    wire new_AGEMA_signal_10754 ;
    wire new_AGEMA_signal_10755 ;
    wire new_AGEMA_signal_10756 ;
    wire new_AGEMA_signal_10757 ;
    wire new_AGEMA_signal_10758 ;
    wire new_AGEMA_signal_10759 ;
    wire new_AGEMA_signal_10760 ;
    wire new_AGEMA_signal_10761 ;
    wire new_AGEMA_signal_10762 ;
    wire new_AGEMA_signal_10763 ;
    wire new_AGEMA_signal_10764 ;
    wire new_AGEMA_signal_10765 ;
    wire new_AGEMA_signal_10766 ;
    wire new_AGEMA_signal_10767 ;
    wire new_AGEMA_signal_10768 ;
    wire new_AGEMA_signal_10769 ;
    wire new_AGEMA_signal_10770 ;
    wire new_AGEMA_signal_10771 ;
    wire new_AGEMA_signal_10772 ;
    wire new_AGEMA_signal_10773 ;
    wire new_AGEMA_signal_10774 ;
    wire new_AGEMA_signal_10775 ;
    wire new_AGEMA_signal_10776 ;
    wire new_AGEMA_signal_10777 ;
    wire new_AGEMA_signal_10778 ;
    wire new_AGEMA_signal_10779 ;
    wire new_AGEMA_signal_10780 ;
    wire new_AGEMA_signal_10781 ;
    wire new_AGEMA_signal_10782 ;
    wire new_AGEMA_signal_10783 ;
    wire new_AGEMA_signal_10784 ;
    wire new_AGEMA_signal_10785 ;
    wire new_AGEMA_signal_10786 ;
    wire new_AGEMA_signal_10787 ;
    wire new_AGEMA_signal_10788 ;
    wire new_AGEMA_signal_10789 ;
    wire new_AGEMA_signal_10790 ;
    wire new_AGEMA_signal_10791 ;
    wire new_AGEMA_signal_10792 ;
    wire new_AGEMA_signal_10793 ;
    wire new_AGEMA_signal_10794 ;
    wire new_AGEMA_signal_10795 ;
    wire new_AGEMA_signal_10796 ;
    wire new_AGEMA_signal_10797 ;
    wire new_AGEMA_signal_10798 ;
    wire new_AGEMA_signal_10799 ;
    wire new_AGEMA_signal_10800 ;
    wire new_AGEMA_signal_10801 ;
    wire new_AGEMA_signal_10802 ;
    wire new_AGEMA_signal_10803 ;
    wire new_AGEMA_signal_10804 ;
    wire new_AGEMA_signal_10805 ;
    wire new_AGEMA_signal_10806 ;
    wire new_AGEMA_signal_10807 ;
    wire new_AGEMA_signal_10808 ;
    wire new_AGEMA_signal_10809 ;
    wire new_AGEMA_signal_10810 ;
    wire new_AGEMA_signal_10811 ;
    wire new_AGEMA_signal_10812 ;
    wire new_AGEMA_signal_10813 ;
    wire new_AGEMA_signal_10814 ;
    wire new_AGEMA_signal_10815 ;
    wire new_AGEMA_signal_10816 ;
    wire new_AGEMA_signal_10817 ;
    wire new_AGEMA_signal_10818 ;
    wire new_AGEMA_signal_10819 ;
    wire new_AGEMA_signal_10820 ;
    wire new_AGEMA_signal_10821 ;
    wire new_AGEMA_signal_10822 ;
    wire new_AGEMA_signal_10823 ;
    wire new_AGEMA_signal_10824 ;
    wire new_AGEMA_signal_10825 ;
    wire new_AGEMA_signal_10826 ;
    wire new_AGEMA_signal_10827 ;
    wire new_AGEMA_signal_10828 ;
    wire new_AGEMA_signal_10829 ;
    wire new_AGEMA_signal_10830 ;
    wire new_AGEMA_signal_10831 ;
    wire new_AGEMA_signal_10832 ;
    wire new_AGEMA_signal_10833 ;
    wire new_AGEMA_signal_10834 ;
    wire new_AGEMA_signal_10835 ;
    wire new_AGEMA_signal_10836 ;
    wire new_AGEMA_signal_10837 ;
    wire new_AGEMA_signal_10838 ;
    wire new_AGEMA_signal_10839 ;
    wire new_AGEMA_signal_10840 ;
    wire new_AGEMA_signal_10841 ;
    wire new_AGEMA_signal_10842 ;
    wire new_AGEMA_signal_10843 ;
    wire new_AGEMA_signal_10844 ;
    wire new_AGEMA_signal_10845 ;
    wire new_AGEMA_signal_10846 ;
    wire new_AGEMA_signal_10847 ;
    wire new_AGEMA_signal_10848 ;
    wire new_AGEMA_signal_10849 ;
    wire new_AGEMA_signal_10850 ;
    wire new_AGEMA_signal_10851 ;
    wire new_AGEMA_signal_10852 ;
    wire new_AGEMA_signal_10853 ;
    wire new_AGEMA_signal_10854 ;
    wire new_AGEMA_signal_10855 ;
    wire new_AGEMA_signal_10856 ;
    wire new_AGEMA_signal_10857 ;
    wire new_AGEMA_signal_10858 ;
    wire new_AGEMA_signal_10859 ;
    wire new_AGEMA_signal_10860 ;
    wire new_AGEMA_signal_10861 ;
    wire new_AGEMA_signal_10862 ;
    wire new_AGEMA_signal_10863 ;
    wire new_AGEMA_signal_10864 ;
    wire new_AGEMA_signal_10865 ;
    wire new_AGEMA_signal_10866 ;
    wire new_AGEMA_signal_10867 ;
    wire new_AGEMA_signal_10868 ;
    wire new_AGEMA_signal_10869 ;
    wire new_AGEMA_signal_10870 ;
    wire new_AGEMA_signal_10871 ;
    wire new_AGEMA_signal_10872 ;
    wire new_AGEMA_signal_10873 ;
    wire new_AGEMA_signal_10874 ;
    wire new_AGEMA_signal_10875 ;
    wire new_AGEMA_signal_10876 ;
    wire new_AGEMA_signal_10877 ;
    wire new_AGEMA_signal_10878 ;
    wire new_AGEMA_signal_10879 ;
    wire new_AGEMA_signal_10880 ;
    wire new_AGEMA_signal_10881 ;
    wire new_AGEMA_signal_10882 ;
    wire new_AGEMA_signal_10883 ;
    wire new_AGEMA_signal_10884 ;
    wire new_AGEMA_signal_10885 ;
    wire new_AGEMA_signal_10886 ;
    wire new_AGEMA_signal_10887 ;
    wire new_AGEMA_signal_10888 ;
    wire new_AGEMA_signal_10889 ;
    wire new_AGEMA_signal_10890 ;
    wire new_AGEMA_signal_10891 ;
    wire new_AGEMA_signal_10892 ;
    wire new_AGEMA_signal_10893 ;
    wire new_AGEMA_signal_10894 ;
    wire new_AGEMA_signal_10895 ;
    wire new_AGEMA_signal_10896 ;
    wire new_AGEMA_signal_10897 ;
    wire new_AGEMA_signal_10898 ;
    wire new_AGEMA_signal_10899 ;
    wire new_AGEMA_signal_10900 ;
    wire new_AGEMA_signal_10901 ;
    wire new_AGEMA_signal_10902 ;
    wire new_AGEMA_signal_10903 ;
    wire new_AGEMA_signal_10904 ;
    wire new_AGEMA_signal_10905 ;
    wire new_AGEMA_signal_10906 ;
    wire new_AGEMA_signal_10907 ;
    wire new_AGEMA_signal_10908 ;
    wire new_AGEMA_signal_10909 ;
    wire new_AGEMA_signal_10910 ;
    wire new_AGEMA_signal_10911 ;
    wire new_AGEMA_signal_10912 ;
    wire new_AGEMA_signal_10913 ;
    wire new_AGEMA_signal_10914 ;
    wire new_AGEMA_signal_10915 ;
    wire new_AGEMA_signal_10916 ;
    wire new_AGEMA_signal_10917 ;
    wire new_AGEMA_signal_10918 ;
    wire new_AGEMA_signal_10919 ;
    wire new_AGEMA_signal_10920 ;
    wire new_AGEMA_signal_10921 ;
    wire new_AGEMA_signal_10922 ;
    wire new_AGEMA_signal_10923 ;
    wire new_AGEMA_signal_10924 ;
    wire new_AGEMA_signal_10925 ;
    wire new_AGEMA_signal_10926 ;
    wire new_AGEMA_signal_10927 ;
    wire new_AGEMA_signal_10928 ;
    wire new_AGEMA_signal_10929 ;
    wire new_AGEMA_signal_10930 ;
    wire new_AGEMA_signal_10931 ;
    wire new_AGEMA_signal_10932 ;
    wire new_AGEMA_signal_10933 ;
    wire new_AGEMA_signal_10934 ;
    wire new_AGEMA_signal_10935 ;
    wire new_AGEMA_signal_10936 ;
    wire new_AGEMA_signal_10937 ;
    wire new_AGEMA_signal_10938 ;
    wire new_AGEMA_signal_10939 ;
    wire new_AGEMA_signal_10940 ;
    wire new_AGEMA_signal_10941 ;
    wire new_AGEMA_signal_10942 ;
    wire new_AGEMA_signal_10943 ;
    wire new_AGEMA_signal_10944 ;
    wire new_AGEMA_signal_10945 ;
    wire new_AGEMA_signal_10946 ;
    wire new_AGEMA_signal_10947 ;
    wire new_AGEMA_signal_10948 ;
    wire new_AGEMA_signal_10949 ;
    wire new_AGEMA_signal_10950 ;
    wire new_AGEMA_signal_10951 ;
    wire new_AGEMA_signal_10952 ;
    wire new_AGEMA_signal_10953 ;
    wire new_AGEMA_signal_10954 ;
    wire new_AGEMA_signal_10955 ;
    wire new_AGEMA_signal_10956 ;
    wire new_AGEMA_signal_10957 ;
    wire new_AGEMA_signal_10958 ;
    wire new_AGEMA_signal_10959 ;
    wire new_AGEMA_signal_10960 ;
    wire new_AGEMA_signal_10961 ;
    wire new_AGEMA_signal_10962 ;
    wire new_AGEMA_signal_10963 ;
    wire new_AGEMA_signal_10964 ;
    wire new_AGEMA_signal_10965 ;
    wire new_AGEMA_signal_10966 ;
    wire new_AGEMA_signal_10967 ;
    wire new_AGEMA_signal_10968 ;
    wire new_AGEMA_signal_10969 ;
    wire new_AGEMA_signal_10970 ;
    wire new_AGEMA_signal_10971 ;
    wire new_AGEMA_signal_10972 ;
    wire new_AGEMA_signal_10973 ;
    wire new_AGEMA_signal_10974 ;
    wire new_AGEMA_signal_10975 ;
    wire new_AGEMA_signal_10976 ;
    wire new_AGEMA_signal_10977 ;
    wire new_AGEMA_signal_10978 ;
    wire new_AGEMA_signal_10979 ;
    wire new_AGEMA_signal_10980 ;
    wire new_AGEMA_signal_10981 ;
    wire new_AGEMA_signal_10982 ;
    wire new_AGEMA_signal_10983 ;
    wire new_AGEMA_signal_10984 ;
    wire new_AGEMA_signal_10985 ;
    wire new_AGEMA_signal_10986 ;
    wire new_AGEMA_signal_10987 ;
    wire new_AGEMA_signal_10988 ;
    wire new_AGEMA_signal_10989 ;
    wire new_AGEMA_signal_10990 ;
    wire new_AGEMA_signal_10991 ;
    wire new_AGEMA_signal_10992 ;
    wire new_AGEMA_signal_10993 ;
    wire new_AGEMA_signal_10994 ;
    wire new_AGEMA_signal_10995 ;
    wire new_AGEMA_signal_10996 ;
    wire new_AGEMA_signal_10997 ;
    wire new_AGEMA_signal_10998 ;
    wire new_AGEMA_signal_10999 ;
    wire new_AGEMA_signal_11000 ;
    wire new_AGEMA_signal_11001 ;
    wire new_AGEMA_signal_11002 ;
    wire new_AGEMA_signal_11003 ;
    wire new_AGEMA_signal_11004 ;
    wire new_AGEMA_signal_11005 ;
    wire new_AGEMA_signal_11006 ;
    wire new_AGEMA_signal_11007 ;
    wire new_AGEMA_signal_11008 ;
    wire new_AGEMA_signal_11009 ;
    wire new_AGEMA_signal_11010 ;
    wire new_AGEMA_signal_11011 ;
    wire new_AGEMA_signal_11012 ;
    wire new_AGEMA_signal_11013 ;
    wire new_AGEMA_signal_11014 ;
    wire new_AGEMA_signal_11015 ;
    wire new_AGEMA_signal_11016 ;
    wire new_AGEMA_signal_11017 ;
    wire new_AGEMA_signal_11018 ;
    wire new_AGEMA_signal_11019 ;
    wire new_AGEMA_signal_11020 ;
    wire new_AGEMA_signal_11021 ;
    wire new_AGEMA_signal_11022 ;
    wire new_AGEMA_signal_11023 ;
    wire new_AGEMA_signal_11024 ;
    wire new_AGEMA_signal_11025 ;
    wire new_AGEMA_signal_11026 ;
    wire new_AGEMA_signal_11027 ;
    wire new_AGEMA_signal_11028 ;
    wire new_AGEMA_signal_11029 ;
    wire new_AGEMA_signal_11030 ;
    wire new_AGEMA_signal_11031 ;
    wire new_AGEMA_signal_11032 ;
    wire new_AGEMA_signal_11033 ;
    wire new_AGEMA_signal_11034 ;
    wire new_AGEMA_signal_11035 ;
    wire new_AGEMA_signal_11036 ;
    wire new_AGEMA_signal_11037 ;
    wire new_AGEMA_signal_11038 ;
    wire new_AGEMA_signal_11039 ;
    wire new_AGEMA_signal_11040 ;
    wire new_AGEMA_signal_11041 ;
    wire new_AGEMA_signal_11042 ;
    wire new_AGEMA_signal_11043 ;
    wire new_AGEMA_signal_11044 ;
    wire new_AGEMA_signal_11045 ;
    wire new_AGEMA_signal_11046 ;
    wire new_AGEMA_signal_11047 ;
    wire new_AGEMA_signal_11048 ;
    wire new_AGEMA_signal_11049 ;
    wire new_AGEMA_signal_11050 ;
    wire new_AGEMA_signal_11051 ;
    wire new_AGEMA_signal_11052 ;
    wire new_AGEMA_signal_11053 ;
    wire new_AGEMA_signal_11054 ;
    wire new_AGEMA_signal_11055 ;
    wire new_AGEMA_signal_11056 ;
    wire new_AGEMA_signal_11057 ;
    wire new_AGEMA_signal_11058 ;
    wire new_AGEMA_signal_11059 ;
    wire new_AGEMA_signal_11060 ;
    wire new_AGEMA_signal_11061 ;
    wire new_AGEMA_signal_11062 ;
    wire new_AGEMA_signal_11063 ;
    wire new_AGEMA_signal_11064 ;
    wire new_AGEMA_signal_11065 ;
    wire new_AGEMA_signal_11066 ;
    wire new_AGEMA_signal_11067 ;
    wire new_AGEMA_signal_11068 ;
    wire new_AGEMA_signal_11069 ;
    wire new_AGEMA_signal_11070 ;
    wire new_AGEMA_signal_11071 ;
    wire new_AGEMA_signal_11072 ;
    wire new_AGEMA_signal_11073 ;
    wire new_AGEMA_signal_11074 ;
    wire new_AGEMA_signal_11075 ;
    wire new_AGEMA_signal_11076 ;
    wire new_AGEMA_signal_11077 ;
    wire new_AGEMA_signal_11078 ;
    wire new_AGEMA_signal_11079 ;
    wire new_AGEMA_signal_11080 ;
    wire new_AGEMA_signal_11081 ;
    wire new_AGEMA_signal_11082 ;
    wire new_AGEMA_signal_11083 ;
    wire new_AGEMA_signal_11084 ;
    wire new_AGEMA_signal_11085 ;
    wire new_AGEMA_signal_11086 ;
    wire new_AGEMA_signal_11087 ;
    wire new_AGEMA_signal_11088 ;
    wire new_AGEMA_signal_11089 ;
    wire new_AGEMA_signal_11090 ;
    wire new_AGEMA_signal_11091 ;
    wire new_AGEMA_signal_11092 ;
    wire new_AGEMA_signal_11093 ;
    wire new_AGEMA_signal_11094 ;
    wire new_AGEMA_signal_11095 ;
    wire new_AGEMA_signal_11096 ;
    wire new_AGEMA_signal_11097 ;
    wire new_AGEMA_signal_11098 ;
    wire new_AGEMA_signal_11099 ;
    wire new_AGEMA_signal_11100 ;
    wire new_AGEMA_signal_11101 ;
    wire new_AGEMA_signal_11102 ;
    wire new_AGEMA_signal_11103 ;
    wire new_AGEMA_signal_11104 ;
    wire new_AGEMA_signal_11105 ;
    wire new_AGEMA_signal_11106 ;
    wire new_AGEMA_signal_11107 ;
    wire new_AGEMA_signal_11108 ;
    wire new_AGEMA_signal_11109 ;
    wire new_AGEMA_signal_11110 ;
    wire new_AGEMA_signal_11111 ;
    wire new_AGEMA_signal_11112 ;
    wire new_AGEMA_signal_11113 ;
    wire new_AGEMA_signal_11114 ;
    wire new_AGEMA_signal_11115 ;
    wire new_AGEMA_signal_11116 ;
    wire new_AGEMA_signal_11117 ;
    wire new_AGEMA_signal_11118 ;
    wire new_AGEMA_signal_11119 ;
    wire new_AGEMA_signal_11120 ;
    wire new_AGEMA_signal_11121 ;
    wire new_AGEMA_signal_11122 ;
    wire new_AGEMA_signal_11123 ;
    wire new_AGEMA_signal_11124 ;
    wire new_AGEMA_signal_11125 ;
    wire new_AGEMA_signal_11126 ;
    wire new_AGEMA_signal_11127 ;
    wire new_AGEMA_signal_11128 ;
    wire new_AGEMA_signal_11129 ;
    wire new_AGEMA_signal_11130 ;
    wire new_AGEMA_signal_11131 ;
    wire new_AGEMA_signal_11132 ;
    wire new_AGEMA_signal_11133 ;
    wire new_AGEMA_signal_11134 ;
    wire new_AGEMA_signal_11135 ;
    wire new_AGEMA_signal_11136 ;
    wire new_AGEMA_signal_11137 ;
    wire new_AGEMA_signal_11138 ;
    wire new_AGEMA_signal_11139 ;
    wire new_AGEMA_signal_11140 ;
    wire new_AGEMA_signal_11141 ;
    wire new_AGEMA_signal_11142 ;
    wire new_AGEMA_signal_11143 ;
    wire new_AGEMA_signal_11144 ;
    wire new_AGEMA_signal_11145 ;
    wire new_AGEMA_signal_11146 ;
    wire new_AGEMA_signal_11147 ;
    wire new_AGEMA_signal_11148 ;
    wire new_AGEMA_signal_11149 ;
    wire new_AGEMA_signal_11150 ;
    wire new_AGEMA_signal_11151 ;
    wire new_AGEMA_signal_11152 ;
    wire new_AGEMA_signal_11153 ;
    wire new_AGEMA_signal_11154 ;
    wire new_AGEMA_signal_11155 ;
    wire new_AGEMA_signal_11156 ;
    wire new_AGEMA_signal_11157 ;
    wire new_AGEMA_signal_11158 ;
    wire new_AGEMA_signal_11159 ;
    wire new_AGEMA_signal_11160 ;
    wire new_AGEMA_signal_11161 ;
    wire new_AGEMA_signal_11162 ;
    wire new_AGEMA_signal_11163 ;
    wire new_AGEMA_signal_11164 ;
    wire new_AGEMA_signal_11165 ;
    wire new_AGEMA_signal_11166 ;
    wire new_AGEMA_signal_11167 ;
    wire new_AGEMA_signal_11168 ;
    wire new_AGEMA_signal_11169 ;
    wire new_AGEMA_signal_11170 ;
    wire new_AGEMA_signal_11171 ;
    wire new_AGEMA_signal_11172 ;
    wire new_AGEMA_signal_11173 ;
    wire new_AGEMA_signal_11174 ;
    wire new_AGEMA_signal_11175 ;
    wire new_AGEMA_signal_11176 ;
    wire new_AGEMA_signal_11177 ;
    wire new_AGEMA_signal_11178 ;
    wire new_AGEMA_signal_11179 ;
    wire new_AGEMA_signal_11180 ;
    wire new_AGEMA_signal_11181 ;
    wire new_AGEMA_signal_11182 ;
    wire new_AGEMA_signal_11183 ;
    wire new_AGEMA_signal_11184 ;
    wire new_AGEMA_signal_11185 ;
    wire new_AGEMA_signal_11186 ;
    wire new_AGEMA_signal_11187 ;
    wire new_AGEMA_signal_11188 ;
    wire new_AGEMA_signal_11189 ;
    wire new_AGEMA_signal_11190 ;
    wire new_AGEMA_signal_11191 ;
    wire new_AGEMA_signal_11192 ;
    wire new_AGEMA_signal_11193 ;
    wire new_AGEMA_signal_11194 ;
    wire new_AGEMA_signal_11195 ;
    wire new_AGEMA_signal_11196 ;
    wire new_AGEMA_signal_11197 ;
    wire new_AGEMA_signal_11198 ;
    wire new_AGEMA_signal_11199 ;
    wire new_AGEMA_signal_11200 ;
    wire new_AGEMA_signal_11201 ;
    wire new_AGEMA_signal_11202 ;
    wire new_AGEMA_signal_11203 ;
    wire new_AGEMA_signal_11204 ;
    wire new_AGEMA_signal_11205 ;
    wire new_AGEMA_signal_11206 ;
    wire new_AGEMA_signal_11207 ;
    wire new_AGEMA_signal_11208 ;
    wire new_AGEMA_signal_11209 ;
    wire new_AGEMA_signal_11210 ;
    wire new_AGEMA_signal_11211 ;
    wire new_AGEMA_signal_11212 ;
    wire new_AGEMA_signal_11213 ;
    wire new_AGEMA_signal_11214 ;
    wire new_AGEMA_signal_11215 ;
    wire new_AGEMA_signal_11216 ;
    wire new_AGEMA_signal_11217 ;
    wire new_AGEMA_signal_11218 ;
    wire new_AGEMA_signal_11219 ;
    wire new_AGEMA_signal_11220 ;
    wire new_AGEMA_signal_11221 ;
    wire new_AGEMA_signal_11222 ;
    wire new_AGEMA_signal_11223 ;
    wire new_AGEMA_signal_11224 ;
    wire new_AGEMA_signal_11225 ;
    wire new_AGEMA_signal_11226 ;
    wire new_AGEMA_signal_11227 ;
    wire new_AGEMA_signal_11228 ;
    wire new_AGEMA_signal_11229 ;
    wire new_AGEMA_signal_11230 ;
    wire new_AGEMA_signal_11231 ;
    wire new_AGEMA_signal_11232 ;
    wire new_AGEMA_signal_11233 ;
    wire new_AGEMA_signal_11234 ;
    wire new_AGEMA_signal_11235 ;
    wire new_AGEMA_signal_11236 ;
    wire new_AGEMA_signal_11237 ;
    wire new_AGEMA_signal_11238 ;
    wire new_AGEMA_signal_11239 ;
    wire new_AGEMA_signal_11240 ;
    wire new_AGEMA_signal_11241 ;
    wire new_AGEMA_signal_11242 ;
    wire new_AGEMA_signal_11243 ;
    wire new_AGEMA_signal_11244 ;
    wire new_AGEMA_signal_11245 ;
    wire new_AGEMA_signal_11246 ;
    wire new_AGEMA_signal_11247 ;
    wire new_AGEMA_signal_11248 ;
    wire new_AGEMA_signal_11249 ;
    wire new_AGEMA_signal_11250 ;
    wire new_AGEMA_signal_11251 ;
    wire new_AGEMA_signal_11252 ;
    wire new_AGEMA_signal_11253 ;
    wire new_AGEMA_signal_11254 ;
    wire new_AGEMA_signal_11255 ;
    wire new_AGEMA_signal_11256 ;
    wire new_AGEMA_signal_11257 ;
    wire new_AGEMA_signal_11258 ;
    wire new_AGEMA_signal_11259 ;
    wire new_AGEMA_signal_11260 ;
    wire new_AGEMA_signal_11261 ;
    wire new_AGEMA_signal_11262 ;
    wire new_AGEMA_signal_11263 ;
    wire new_AGEMA_signal_11264 ;
    wire new_AGEMA_signal_11265 ;
    wire new_AGEMA_signal_11266 ;
    wire new_AGEMA_signal_11267 ;
    wire new_AGEMA_signal_11268 ;
    wire new_AGEMA_signal_11269 ;
    wire new_AGEMA_signal_11270 ;
    wire new_AGEMA_signal_11271 ;
    wire new_AGEMA_signal_11272 ;
    wire new_AGEMA_signal_11273 ;
    wire new_AGEMA_signal_11274 ;
    wire new_AGEMA_signal_11275 ;
    wire new_AGEMA_signal_11276 ;
    wire new_AGEMA_signal_11277 ;
    wire new_AGEMA_signal_11278 ;
    wire new_AGEMA_signal_11279 ;
    wire new_AGEMA_signal_11280 ;
    wire new_AGEMA_signal_11281 ;
    wire new_AGEMA_signal_11282 ;
    wire new_AGEMA_signal_11283 ;
    wire new_AGEMA_signal_11284 ;
    wire new_AGEMA_signal_11285 ;
    wire new_AGEMA_signal_11286 ;
    wire new_AGEMA_signal_11287 ;
    wire new_AGEMA_signal_11288 ;
    wire new_AGEMA_signal_11289 ;
    wire new_AGEMA_signal_11290 ;
    wire new_AGEMA_signal_11291 ;
    wire new_AGEMA_signal_11292 ;
    wire new_AGEMA_signal_11293 ;
    wire new_AGEMA_signal_11294 ;
    wire new_AGEMA_signal_11295 ;
    wire new_AGEMA_signal_11296 ;
    wire new_AGEMA_signal_11297 ;
    wire new_AGEMA_signal_11298 ;
    wire new_AGEMA_signal_11299 ;
    wire new_AGEMA_signal_11300 ;
    wire new_AGEMA_signal_11301 ;
    wire new_AGEMA_signal_11302 ;
    wire new_AGEMA_signal_11303 ;
    wire new_AGEMA_signal_11304 ;
    wire new_AGEMA_signal_11305 ;
    wire new_AGEMA_signal_11306 ;
    wire new_AGEMA_signal_11307 ;
    wire new_AGEMA_signal_11308 ;
    wire new_AGEMA_signal_11309 ;
    wire new_AGEMA_signal_11310 ;
    wire new_AGEMA_signal_11311 ;
    wire new_AGEMA_signal_11312 ;
    wire new_AGEMA_signal_11313 ;
    wire new_AGEMA_signal_11314 ;
    wire new_AGEMA_signal_11315 ;
    wire new_AGEMA_signal_11316 ;
    wire new_AGEMA_signal_11317 ;
    wire new_AGEMA_signal_11318 ;
    wire new_AGEMA_signal_11319 ;
    wire new_AGEMA_signal_11320 ;
    wire new_AGEMA_signal_11321 ;
    wire new_AGEMA_signal_11322 ;
    wire new_AGEMA_signal_11323 ;
    wire new_AGEMA_signal_11324 ;
    wire new_AGEMA_signal_11325 ;
    wire new_AGEMA_signal_11326 ;
    wire new_AGEMA_signal_11327 ;
    wire new_AGEMA_signal_11328 ;
    wire new_AGEMA_signal_11329 ;
    wire new_AGEMA_signal_11330 ;
    wire new_AGEMA_signal_11331 ;
    wire new_AGEMA_signal_11332 ;
    wire new_AGEMA_signal_11333 ;
    wire new_AGEMA_signal_11334 ;
    wire new_AGEMA_signal_11335 ;
    wire new_AGEMA_signal_11336 ;
    wire new_AGEMA_signal_11337 ;
    wire new_AGEMA_signal_11338 ;
    wire new_AGEMA_signal_11339 ;
    wire new_AGEMA_signal_11340 ;
    wire new_AGEMA_signal_11341 ;
    wire new_AGEMA_signal_11342 ;
    wire new_AGEMA_signal_11343 ;
    wire new_AGEMA_signal_11344 ;
    wire new_AGEMA_signal_11345 ;
    wire new_AGEMA_signal_11346 ;
    wire new_AGEMA_signal_11347 ;
    wire new_AGEMA_signal_11348 ;
    wire new_AGEMA_signal_11349 ;
    wire new_AGEMA_signal_11350 ;
    wire new_AGEMA_signal_11351 ;
    wire new_AGEMA_signal_11352 ;
    wire new_AGEMA_signal_11353 ;
    wire new_AGEMA_signal_11354 ;
    wire new_AGEMA_signal_11355 ;
    wire new_AGEMA_signal_11356 ;
    wire new_AGEMA_signal_11357 ;
    wire new_AGEMA_signal_11358 ;
    wire new_AGEMA_signal_11359 ;
    wire new_AGEMA_signal_11360 ;
    wire new_AGEMA_signal_11361 ;
    wire new_AGEMA_signal_11362 ;
    wire new_AGEMA_signal_11363 ;
    wire new_AGEMA_signal_11364 ;
    wire new_AGEMA_signal_11365 ;
    wire new_AGEMA_signal_11366 ;
    wire new_AGEMA_signal_11367 ;
    wire new_AGEMA_signal_11368 ;
    wire new_AGEMA_signal_11369 ;
    wire new_AGEMA_signal_11370 ;
    wire new_AGEMA_signal_11371 ;
    wire new_AGEMA_signal_11372 ;
    wire new_AGEMA_signal_11373 ;
    wire new_AGEMA_signal_11374 ;
    wire new_AGEMA_signal_11375 ;
    wire new_AGEMA_signal_11376 ;
    wire new_AGEMA_signal_11377 ;
    wire new_AGEMA_signal_11378 ;
    wire new_AGEMA_signal_11379 ;
    wire new_AGEMA_signal_11380 ;
    wire new_AGEMA_signal_11381 ;
    wire new_AGEMA_signal_11382 ;
    wire new_AGEMA_signal_11383 ;
    wire new_AGEMA_signal_11384 ;
    wire new_AGEMA_signal_11385 ;
    wire new_AGEMA_signal_11386 ;
    wire new_AGEMA_signal_11387 ;
    wire new_AGEMA_signal_11388 ;
    wire new_AGEMA_signal_11389 ;
    wire new_AGEMA_signal_11390 ;
    wire new_AGEMA_signal_11391 ;
    wire new_AGEMA_signal_11392 ;
    wire new_AGEMA_signal_11393 ;
    wire new_AGEMA_signal_11394 ;
    wire new_AGEMA_signal_11395 ;
    wire new_AGEMA_signal_11396 ;
    wire new_AGEMA_signal_11397 ;
    wire new_AGEMA_signal_11398 ;
    wire new_AGEMA_signal_11399 ;
    wire new_AGEMA_signal_11400 ;
    wire new_AGEMA_signal_11401 ;
    wire new_AGEMA_signal_11402 ;
    wire new_AGEMA_signal_11403 ;
    wire new_AGEMA_signal_11404 ;
    wire new_AGEMA_signal_11405 ;
    wire new_AGEMA_signal_11406 ;
    wire new_AGEMA_signal_11407 ;
    wire new_AGEMA_signal_11408 ;
    wire new_AGEMA_signal_11409 ;
    wire new_AGEMA_signal_11410 ;
    wire new_AGEMA_signal_11411 ;
    wire new_AGEMA_signal_11412 ;
    wire new_AGEMA_signal_11413 ;
    wire new_AGEMA_signal_11414 ;
    wire new_AGEMA_signal_11415 ;
    wire new_AGEMA_signal_11416 ;
    wire new_AGEMA_signal_11417 ;
    wire new_AGEMA_signal_11418 ;
    wire new_AGEMA_signal_11419 ;
    wire new_AGEMA_signal_11420 ;
    wire new_AGEMA_signal_11421 ;
    wire new_AGEMA_signal_11422 ;
    wire new_AGEMA_signal_11423 ;
    wire new_AGEMA_signal_11424 ;
    wire new_AGEMA_signal_11425 ;
    wire new_AGEMA_signal_11426 ;
    wire new_AGEMA_signal_11427 ;
    wire new_AGEMA_signal_11428 ;
    wire new_AGEMA_signal_11429 ;
    wire new_AGEMA_signal_11430 ;
    wire new_AGEMA_signal_11431 ;
    wire new_AGEMA_signal_11432 ;
    wire new_AGEMA_signal_11433 ;
    wire new_AGEMA_signal_11434 ;
    wire new_AGEMA_signal_11435 ;
    wire new_AGEMA_signal_11436 ;
    wire new_AGEMA_signal_11437 ;
    wire new_AGEMA_signal_11438 ;
    wire new_AGEMA_signal_11439 ;
    wire new_AGEMA_signal_11440 ;
    wire new_AGEMA_signal_11441 ;
    wire new_AGEMA_signal_11442 ;
    wire new_AGEMA_signal_11443 ;
    wire new_AGEMA_signal_11444 ;
    wire new_AGEMA_signal_11445 ;
    wire new_AGEMA_signal_11446 ;
    wire new_AGEMA_signal_11447 ;
    wire new_AGEMA_signal_11448 ;
    wire new_AGEMA_signal_11449 ;
    wire new_AGEMA_signal_11450 ;
    wire new_AGEMA_signal_11451 ;
    wire new_AGEMA_signal_11452 ;
    wire new_AGEMA_signal_11453 ;
    wire new_AGEMA_signal_11454 ;
    wire new_AGEMA_signal_11455 ;
    wire new_AGEMA_signal_11456 ;
    wire new_AGEMA_signal_11457 ;
    wire new_AGEMA_signal_11458 ;
    wire new_AGEMA_signal_11459 ;
    wire new_AGEMA_signal_11460 ;
    wire new_AGEMA_signal_11461 ;
    wire new_AGEMA_signal_11462 ;
    wire new_AGEMA_signal_11463 ;
    wire new_AGEMA_signal_11464 ;
    wire new_AGEMA_signal_11465 ;
    wire new_AGEMA_signal_11466 ;
    wire new_AGEMA_signal_11467 ;
    wire new_AGEMA_signal_11468 ;
    wire new_AGEMA_signal_11469 ;
    wire new_AGEMA_signal_11470 ;
    wire new_AGEMA_signal_11471 ;
    wire new_AGEMA_signal_11472 ;
    wire new_AGEMA_signal_11473 ;
    wire new_AGEMA_signal_11474 ;
    wire new_AGEMA_signal_11475 ;
    wire new_AGEMA_signal_11476 ;
    wire new_AGEMA_signal_11477 ;
    wire new_AGEMA_signal_11478 ;
    wire new_AGEMA_signal_11479 ;
    wire new_AGEMA_signal_11480 ;
    wire new_AGEMA_signal_11481 ;
    wire new_AGEMA_signal_11482 ;
    wire new_AGEMA_signal_11483 ;
    wire new_AGEMA_signal_11484 ;
    wire new_AGEMA_signal_11485 ;
    wire new_AGEMA_signal_11486 ;
    wire new_AGEMA_signal_11487 ;
    wire new_AGEMA_signal_11488 ;
    wire new_AGEMA_signal_11489 ;
    wire new_AGEMA_signal_11490 ;
    wire new_AGEMA_signal_11491 ;
    wire new_AGEMA_signal_11492 ;
    wire new_AGEMA_signal_11493 ;
    wire new_AGEMA_signal_11494 ;
    wire new_AGEMA_signal_11495 ;
    wire new_AGEMA_signal_11496 ;
    wire new_AGEMA_signal_11497 ;
    wire new_AGEMA_signal_11498 ;
    wire new_AGEMA_signal_11499 ;
    wire new_AGEMA_signal_11500 ;
    wire new_AGEMA_signal_11501 ;
    wire new_AGEMA_signal_11502 ;
    wire new_AGEMA_signal_11503 ;
    wire new_AGEMA_signal_11504 ;
    wire new_AGEMA_signal_11505 ;
    wire new_AGEMA_signal_11506 ;
    wire new_AGEMA_signal_11507 ;
    wire new_AGEMA_signal_11508 ;
    wire new_AGEMA_signal_11509 ;
    wire new_AGEMA_signal_11510 ;
    wire new_AGEMA_signal_11511 ;
    wire new_AGEMA_signal_11512 ;
    wire new_AGEMA_signal_11513 ;
    wire new_AGEMA_signal_11514 ;
    wire new_AGEMA_signal_11515 ;
    wire new_AGEMA_signal_11516 ;
    wire new_AGEMA_signal_11517 ;
    wire new_AGEMA_signal_11518 ;
    wire new_AGEMA_signal_11519 ;
    wire new_AGEMA_signal_11520 ;
    wire new_AGEMA_signal_11521 ;
    wire new_AGEMA_signal_11522 ;
    wire new_AGEMA_signal_11523 ;
    wire new_AGEMA_signal_11524 ;
    wire new_AGEMA_signal_11525 ;
    wire new_AGEMA_signal_11526 ;
    wire new_AGEMA_signal_11527 ;
    wire new_AGEMA_signal_11528 ;
    wire new_AGEMA_signal_11529 ;
    wire new_AGEMA_signal_11530 ;
    wire new_AGEMA_signal_11531 ;
    wire new_AGEMA_signal_11532 ;
    wire new_AGEMA_signal_11533 ;
    wire new_AGEMA_signal_11534 ;
    wire new_AGEMA_signal_11535 ;
    wire new_AGEMA_signal_11536 ;
    wire new_AGEMA_signal_11537 ;
    wire new_AGEMA_signal_11538 ;
    wire new_AGEMA_signal_11539 ;
    wire new_AGEMA_signal_11540 ;
    wire new_AGEMA_signal_11541 ;
    wire new_AGEMA_signal_11542 ;
    wire new_AGEMA_signal_11543 ;
    wire new_AGEMA_signal_11544 ;
    wire new_AGEMA_signal_11545 ;
    wire new_AGEMA_signal_11546 ;
    wire new_AGEMA_signal_11547 ;
    wire new_AGEMA_signal_11548 ;
    wire new_AGEMA_signal_11549 ;
    wire new_AGEMA_signal_11550 ;
    wire new_AGEMA_signal_11551 ;
    wire new_AGEMA_signal_11552 ;
    wire new_AGEMA_signal_11553 ;
    wire new_AGEMA_signal_11554 ;
    wire new_AGEMA_signal_11555 ;
    wire new_AGEMA_signal_11556 ;
    wire new_AGEMA_signal_11557 ;
    wire new_AGEMA_signal_11558 ;
    wire new_AGEMA_signal_11559 ;
    wire new_AGEMA_signal_11560 ;
    wire new_AGEMA_signal_11561 ;
    wire new_AGEMA_signal_11562 ;
    wire new_AGEMA_signal_11563 ;
    wire new_AGEMA_signal_11564 ;
    wire new_AGEMA_signal_11565 ;
    wire new_AGEMA_signal_11566 ;
    wire new_AGEMA_signal_11567 ;
    wire new_AGEMA_signal_11568 ;
    wire new_AGEMA_signal_11569 ;
    wire new_AGEMA_signal_11570 ;
    wire new_AGEMA_signal_11571 ;
    wire new_AGEMA_signal_11572 ;
    wire new_AGEMA_signal_11573 ;
    wire new_AGEMA_signal_11574 ;
    wire new_AGEMA_signal_11575 ;
    wire new_AGEMA_signal_11576 ;
    wire new_AGEMA_signal_11577 ;
    wire new_AGEMA_signal_11578 ;
    wire new_AGEMA_signal_11579 ;
    wire new_AGEMA_signal_11580 ;
    wire new_AGEMA_signal_11581 ;
    wire new_AGEMA_signal_11582 ;
    wire new_AGEMA_signal_11583 ;
    wire new_AGEMA_signal_11584 ;
    wire new_AGEMA_signal_11585 ;
    wire new_AGEMA_signal_11586 ;
    wire new_AGEMA_signal_11587 ;
    wire new_AGEMA_signal_11588 ;
    wire new_AGEMA_signal_11589 ;
    wire new_AGEMA_signal_11590 ;
    wire new_AGEMA_signal_11591 ;
    wire new_AGEMA_signal_11592 ;
    wire new_AGEMA_signal_11593 ;
    wire new_AGEMA_signal_11594 ;
    wire new_AGEMA_signal_11595 ;
    wire new_AGEMA_signal_11596 ;
    wire new_AGEMA_signal_11597 ;
    wire new_AGEMA_signal_11598 ;
    wire new_AGEMA_signal_11599 ;
    wire new_AGEMA_signal_11600 ;
    wire new_AGEMA_signal_11601 ;
    wire new_AGEMA_signal_11602 ;
    wire new_AGEMA_signal_11603 ;
    wire new_AGEMA_signal_11604 ;
    wire new_AGEMA_signal_11605 ;
    wire new_AGEMA_signal_11606 ;
    wire new_AGEMA_signal_11607 ;
    wire new_AGEMA_signal_11608 ;
    wire new_AGEMA_signal_11609 ;
    wire new_AGEMA_signal_11610 ;
    wire new_AGEMA_signal_11611 ;
    wire new_AGEMA_signal_11612 ;
    wire new_AGEMA_signal_11613 ;
    wire new_AGEMA_signal_11614 ;
    wire new_AGEMA_signal_11615 ;
    wire new_AGEMA_signal_11616 ;
    wire new_AGEMA_signal_11617 ;
    wire new_AGEMA_signal_11618 ;
    wire new_AGEMA_signal_11619 ;
    wire new_AGEMA_signal_11620 ;
    wire new_AGEMA_signal_11621 ;
    wire new_AGEMA_signal_11622 ;
    wire new_AGEMA_signal_11623 ;
    wire new_AGEMA_signal_11624 ;
    wire new_AGEMA_signal_11625 ;
    wire new_AGEMA_signal_11626 ;
    wire new_AGEMA_signal_11627 ;
    wire new_AGEMA_signal_11628 ;
    wire new_AGEMA_signal_11629 ;
    wire new_AGEMA_signal_11630 ;
    wire new_AGEMA_signal_11631 ;
    wire new_AGEMA_signal_11632 ;
    wire new_AGEMA_signal_11633 ;
    wire new_AGEMA_signal_11634 ;
    wire new_AGEMA_signal_11635 ;
    wire new_AGEMA_signal_11636 ;
    wire new_AGEMA_signal_11637 ;
    wire new_AGEMA_signal_11638 ;
    wire new_AGEMA_signal_11639 ;
    wire new_AGEMA_signal_11640 ;
    wire new_AGEMA_signal_11641 ;
    wire new_AGEMA_signal_11642 ;
    wire new_AGEMA_signal_11643 ;
    wire new_AGEMA_signal_11644 ;
    wire new_AGEMA_signal_11645 ;
    wire new_AGEMA_signal_11646 ;
    wire new_AGEMA_signal_11647 ;
    wire new_AGEMA_signal_11648 ;
    wire new_AGEMA_signal_11649 ;
    wire new_AGEMA_signal_11650 ;
    wire new_AGEMA_signal_11651 ;
    wire new_AGEMA_signal_11652 ;
    wire new_AGEMA_signal_11653 ;
    wire new_AGEMA_signal_11654 ;
    wire new_AGEMA_signal_11655 ;
    wire new_AGEMA_signal_11656 ;
    wire new_AGEMA_signal_11657 ;
    wire new_AGEMA_signal_11658 ;
    wire new_AGEMA_signal_11659 ;
    wire new_AGEMA_signal_11660 ;
    wire new_AGEMA_signal_11661 ;
    wire new_AGEMA_signal_11662 ;
    wire new_AGEMA_signal_11663 ;
    wire new_AGEMA_signal_11664 ;
    wire new_AGEMA_signal_11665 ;
    wire new_AGEMA_signal_11666 ;
    wire new_AGEMA_signal_11667 ;
    wire new_AGEMA_signal_11668 ;
    wire new_AGEMA_signal_11669 ;
    wire new_AGEMA_signal_11670 ;
    wire new_AGEMA_signal_11671 ;
    wire new_AGEMA_signal_11672 ;
    wire new_AGEMA_signal_11673 ;
    wire new_AGEMA_signal_11674 ;
    wire new_AGEMA_signal_11675 ;
    wire new_AGEMA_signal_11676 ;
    wire new_AGEMA_signal_11677 ;
    wire new_AGEMA_signal_11678 ;
    wire new_AGEMA_signal_11679 ;
    wire new_AGEMA_signal_11680 ;
    wire new_AGEMA_signal_11681 ;
    wire new_AGEMA_signal_11682 ;
    wire new_AGEMA_signal_11683 ;
    wire new_AGEMA_signal_11684 ;
    wire new_AGEMA_signal_11685 ;
    wire new_AGEMA_signal_11686 ;
    wire new_AGEMA_signal_11687 ;
    wire new_AGEMA_signal_11688 ;
    wire new_AGEMA_signal_11689 ;
    wire new_AGEMA_signal_11690 ;
    wire new_AGEMA_signal_11691 ;
    wire new_AGEMA_signal_11692 ;
    wire new_AGEMA_signal_11693 ;
    wire new_AGEMA_signal_11694 ;
    wire new_AGEMA_signal_11695 ;
    wire new_AGEMA_signal_11696 ;
    wire new_AGEMA_signal_11697 ;
    wire new_AGEMA_signal_11698 ;
    wire new_AGEMA_signal_11699 ;
    wire new_AGEMA_signal_11700 ;
    wire new_AGEMA_signal_11701 ;
    wire new_AGEMA_signal_11702 ;
    wire new_AGEMA_signal_11703 ;
    wire new_AGEMA_signal_11704 ;
    wire new_AGEMA_signal_11705 ;
    wire new_AGEMA_signal_11706 ;
    wire new_AGEMA_signal_11707 ;
    wire new_AGEMA_signal_11708 ;
    wire new_AGEMA_signal_11709 ;
    wire new_AGEMA_signal_11710 ;
    wire new_AGEMA_signal_11711 ;
    wire new_AGEMA_signal_11712 ;
    wire new_AGEMA_signal_11713 ;
    wire new_AGEMA_signal_11714 ;
    wire new_AGEMA_signal_11715 ;
    wire new_AGEMA_signal_11716 ;
    wire new_AGEMA_signal_11717 ;
    wire new_AGEMA_signal_11718 ;
    wire new_AGEMA_signal_11719 ;
    wire new_AGEMA_signal_11720 ;
    wire new_AGEMA_signal_11721 ;
    wire new_AGEMA_signal_11722 ;
    wire new_AGEMA_signal_11723 ;
    wire new_AGEMA_signal_11724 ;
    wire new_AGEMA_signal_11725 ;
    wire new_AGEMA_signal_11726 ;
    wire new_AGEMA_signal_11727 ;
    wire new_AGEMA_signal_11728 ;
    wire new_AGEMA_signal_11729 ;
    wire new_AGEMA_signal_11730 ;
    wire new_AGEMA_signal_11731 ;
    wire new_AGEMA_signal_11732 ;
    wire new_AGEMA_signal_11733 ;
    wire new_AGEMA_signal_11734 ;
    wire new_AGEMA_signal_11735 ;
    wire new_AGEMA_signal_11736 ;
    wire new_AGEMA_signal_11737 ;
    wire new_AGEMA_signal_11738 ;
    wire new_AGEMA_signal_11739 ;
    wire new_AGEMA_signal_11740 ;
    wire new_AGEMA_signal_11741 ;
    wire new_AGEMA_signal_11742 ;
    wire new_AGEMA_signal_11743 ;
    wire new_AGEMA_signal_11744 ;
    wire new_AGEMA_signal_11745 ;
    wire new_AGEMA_signal_11746 ;
    wire new_AGEMA_signal_11747 ;
    wire new_AGEMA_signal_11748 ;
    wire new_AGEMA_signal_11749 ;
    wire new_AGEMA_signal_11750 ;
    wire new_AGEMA_signal_11751 ;
    wire new_AGEMA_signal_11752 ;
    wire new_AGEMA_signal_11753 ;
    wire new_AGEMA_signal_11754 ;
    wire new_AGEMA_signal_11755 ;
    wire new_AGEMA_signal_11756 ;
    wire new_AGEMA_signal_11757 ;
    wire new_AGEMA_signal_11758 ;
    wire new_AGEMA_signal_11759 ;
    wire new_AGEMA_signal_11760 ;
    wire new_AGEMA_signal_11761 ;
    wire new_AGEMA_signal_11762 ;
    wire new_AGEMA_signal_11763 ;
    wire new_AGEMA_signal_11764 ;
    wire new_AGEMA_signal_11765 ;
    wire new_AGEMA_signal_11766 ;
    wire new_AGEMA_signal_11767 ;
    wire new_AGEMA_signal_11768 ;
    wire new_AGEMA_signal_11769 ;
    wire new_AGEMA_signal_11770 ;
    wire new_AGEMA_signal_11771 ;
    wire new_AGEMA_signal_11772 ;
    wire new_AGEMA_signal_11773 ;
    wire new_AGEMA_signal_11774 ;
    wire new_AGEMA_signal_11775 ;
    wire new_AGEMA_signal_11776 ;
    wire new_AGEMA_signal_11777 ;
    wire new_AGEMA_signal_11778 ;
    wire new_AGEMA_signal_11779 ;
    wire new_AGEMA_signal_11780 ;
    wire new_AGEMA_signal_11781 ;
    wire new_AGEMA_signal_11782 ;
    wire new_AGEMA_signal_11783 ;
    wire new_AGEMA_signal_11784 ;
    wire new_AGEMA_signal_11785 ;
    wire new_AGEMA_signal_11786 ;
    wire new_AGEMA_signal_11787 ;
    wire new_AGEMA_signal_11788 ;
    wire new_AGEMA_signal_11789 ;
    wire new_AGEMA_signal_11790 ;
    wire new_AGEMA_signal_11791 ;
    wire new_AGEMA_signal_11792 ;
    wire new_AGEMA_signal_11793 ;
    wire new_AGEMA_signal_11794 ;
    wire new_AGEMA_signal_11795 ;
    wire new_AGEMA_signal_11796 ;
    wire new_AGEMA_signal_11797 ;
    wire new_AGEMA_signal_11798 ;
    wire new_AGEMA_signal_11799 ;
    wire new_AGEMA_signal_11800 ;
    wire new_AGEMA_signal_11801 ;
    wire new_AGEMA_signal_11802 ;
    wire new_AGEMA_signal_11803 ;
    wire new_AGEMA_signal_11804 ;
    wire new_AGEMA_signal_11805 ;
    wire new_AGEMA_signal_11806 ;
    wire new_AGEMA_signal_11807 ;
    wire new_AGEMA_signal_11808 ;
    wire new_AGEMA_signal_11809 ;
    wire new_AGEMA_signal_11810 ;
    wire new_AGEMA_signal_11811 ;
    wire new_AGEMA_signal_11812 ;
    wire new_AGEMA_signal_11813 ;
    wire new_AGEMA_signal_11814 ;
    wire new_AGEMA_signal_11815 ;
    wire new_AGEMA_signal_11816 ;
    wire new_AGEMA_signal_11817 ;
    wire new_AGEMA_signal_11818 ;
    wire new_AGEMA_signal_11819 ;
    wire new_AGEMA_signal_11820 ;
    wire new_AGEMA_signal_11821 ;
    wire new_AGEMA_signal_11822 ;
    wire new_AGEMA_signal_11823 ;
    wire new_AGEMA_signal_11824 ;
    wire new_AGEMA_signal_11825 ;
    wire new_AGEMA_signal_11826 ;
    wire new_AGEMA_signal_11827 ;
    wire new_AGEMA_signal_11828 ;
    wire new_AGEMA_signal_11829 ;
    wire new_AGEMA_signal_11830 ;
    wire new_AGEMA_signal_11831 ;
    wire new_AGEMA_signal_11832 ;
    wire new_AGEMA_signal_11833 ;
    wire new_AGEMA_signal_11834 ;
    wire new_AGEMA_signal_11835 ;
    wire new_AGEMA_signal_11836 ;
    wire new_AGEMA_signal_11837 ;
    wire new_AGEMA_signal_11838 ;
    wire new_AGEMA_signal_11839 ;
    wire new_AGEMA_signal_11840 ;
    wire new_AGEMA_signal_11841 ;
    wire new_AGEMA_signal_11842 ;
    wire new_AGEMA_signal_11843 ;
    wire new_AGEMA_signal_11844 ;
    wire new_AGEMA_signal_11845 ;
    wire new_AGEMA_signal_11846 ;
    wire new_AGEMA_signal_11847 ;
    wire new_AGEMA_signal_11848 ;
    wire new_AGEMA_signal_11849 ;
    wire new_AGEMA_signal_11850 ;
    wire new_AGEMA_signal_11851 ;
    wire new_AGEMA_signal_11852 ;
    wire new_AGEMA_signal_11853 ;
    wire new_AGEMA_signal_11854 ;
    wire new_AGEMA_signal_11855 ;
    wire new_AGEMA_signal_11856 ;
    wire new_AGEMA_signal_11857 ;
    wire new_AGEMA_signal_11858 ;
    wire new_AGEMA_signal_11859 ;
    wire new_AGEMA_signal_11860 ;
    wire new_AGEMA_signal_11861 ;
    wire new_AGEMA_signal_11862 ;
    wire new_AGEMA_signal_11863 ;
    wire new_AGEMA_signal_11864 ;
    wire new_AGEMA_signal_11865 ;
    wire new_AGEMA_signal_11866 ;
    wire new_AGEMA_signal_11867 ;
    wire new_AGEMA_signal_11868 ;
    wire new_AGEMA_signal_11869 ;
    wire new_AGEMA_signal_11870 ;
    wire new_AGEMA_signal_11871 ;
    wire new_AGEMA_signal_11872 ;
    wire new_AGEMA_signal_11873 ;
    wire new_AGEMA_signal_11874 ;
    wire new_AGEMA_signal_11875 ;
    wire new_AGEMA_signal_11876 ;
    wire new_AGEMA_signal_11877 ;
    wire new_AGEMA_signal_11878 ;
    wire new_AGEMA_signal_11879 ;
    wire new_AGEMA_signal_11880 ;
    wire new_AGEMA_signal_11881 ;
    wire new_AGEMA_signal_11882 ;
    wire new_AGEMA_signal_11883 ;
    wire new_AGEMA_signal_11884 ;
    wire new_AGEMA_signal_11885 ;
    wire new_AGEMA_signal_11886 ;
    wire new_AGEMA_signal_11887 ;
    wire new_AGEMA_signal_11888 ;
    wire new_AGEMA_signal_11889 ;
    wire new_AGEMA_signal_11890 ;
    wire new_AGEMA_signal_11891 ;
    wire new_AGEMA_signal_11892 ;
    wire new_AGEMA_signal_11893 ;
    wire new_AGEMA_signal_11894 ;
    wire new_AGEMA_signal_11895 ;
    wire new_AGEMA_signal_11896 ;
    wire new_AGEMA_signal_11897 ;
    wire new_AGEMA_signal_11898 ;
    wire new_AGEMA_signal_11899 ;
    wire new_AGEMA_signal_11900 ;
    wire new_AGEMA_signal_11901 ;
    wire new_AGEMA_signal_11902 ;
    wire new_AGEMA_signal_11903 ;
    wire new_AGEMA_signal_11904 ;
    wire new_AGEMA_signal_11905 ;
    wire new_AGEMA_signal_11906 ;
    wire new_AGEMA_signal_11907 ;
    wire new_AGEMA_signal_11908 ;
    wire new_AGEMA_signal_11909 ;
    wire new_AGEMA_signal_11910 ;
    wire new_AGEMA_signal_11911 ;
    wire new_AGEMA_signal_11912 ;
    wire new_AGEMA_signal_11913 ;
    wire new_AGEMA_signal_11914 ;
    wire new_AGEMA_signal_11915 ;
    wire new_AGEMA_signal_11916 ;
    wire new_AGEMA_signal_11917 ;
    wire new_AGEMA_signal_11918 ;
    wire new_AGEMA_signal_11919 ;
    wire new_AGEMA_signal_11920 ;
    wire new_AGEMA_signal_11921 ;
    wire new_AGEMA_signal_11922 ;
    wire new_AGEMA_signal_11923 ;
    wire new_AGEMA_signal_11924 ;
    wire new_AGEMA_signal_11925 ;
    wire new_AGEMA_signal_11926 ;
    wire new_AGEMA_signal_11927 ;
    wire new_AGEMA_signal_11928 ;
    wire new_AGEMA_signal_11929 ;
    wire new_AGEMA_signal_11930 ;
    wire new_AGEMA_signal_11931 ;
    wire new_AGEMA_signal_11932 ;
    wire new_AGEMA_signal_11933 ;
    wire new_AGEMA_signal_11934 ;
    wire new_AGEMA_signal_11935 ;
    wire new_AGEMA_signal_11936 ;
    wire new_AGEMA_signal_11937 ;
    wire new_AGEMA_signal_11938 ;
    wire new_AGEMA_signal_11939 ;
    wire new_AGEMA_signal_11940 ;
    wire new_AGEMA_signal_11941 ;
    wire new_AGEMA_signal_11942 ;
    wire new_AGEMA_signal_11943 ;
    wire new_AGEMA_signal_11944 ;
    wire new_AGEMA_signal_11945 ;
    wire new_AGEMA_signal_11946 ;
    wire new_AGEMA_signal_11947 ;
    wire new_AGEMA_signal_11948 ;
    wire new_AGEMA_signal_11949 ;
    wire new_AGEMA_signal_11950 ;
    wire new_AGEMA_signal_11951 ;
    wire new_AGEMA_signal_11952 ;
    wire new_AGEMA_signal_11953 ;
    wire new_AGEMA_signal_11954 ;
    wire new_AGEMA_signal_11955 ;
    wire new_AGEMA_signal_11956 ;
    wire new_AGEMA_signal_11957 ;
    wire new_AGEMA_signal_11958 ;
    wire new_AGEMA_signal_11959 ;
    wire new_AGEMA_signal_11960 ;
    wire new_AGEMA_signal_11961 ;
    wire new_AGEMA_signal_11962 ;
    wire new_AGEMA_signal_11963 ;
    wire new_AGEMA_signal_11964 ;
    wire new_AGEMA_signal_11965 ;
    wire new_AGEMA_signal_11966 ;
    wire new_AGEMA_signal_11967 ;
    wire new_AGEMA_signal_11968 ;
    wire new_AGEMA_signal_11969 ;
    wire new_AGEMA_signal_11970 ;
    wire new_AGEMA_signal_11971 ;
    wire new_AGEMA_signal_11972 ;
    wire new_AGEMA_signal_11973 ;
    wire new_AGEMA_signal_11974 ;
    wire new_AGEMA_signal_11975 ;
    wire new_AGEMA_signal_11976 ;
    wire new_AGEMA_signal_11977 ;
    wire new_AGEMA_signal_11978 ;
    wire new_AGEMA_signal_11979 ;
    wire new_AGEMA_signal_11980 ;
    wire new_AGEMA_signal_11981 ;
    wire new_AGEMA_signal_11982 ;
    wire new_AGEMA_signal_11983 ;
    wire new_AGEMA_signal_11984 ;
    wire new_AGEMA_signal_11985 ;
    wire new_AGEMA_signal_11986 ;
    wire new_AGEMA_signal_11987 ;
    wire new_AGEMA_signal_11988 ;
    wire new_AGEMA_signal_11989 ;
    wire new_AGEMA_signal_11990 ;
    wire new_AGEMA_signal_11991 ;
    wire new_AGEMA_signal_11992 ;
    wire new_AGEMA_signal_11993 ;
    wire new_AGEMA_signal_11994 ;
    wire new_AGEMA_signal_11995 ;
    wire new_AGEMA_signal_11996 ;
    wire new_AGEMA_signal_11997 ;
    wire new_AGEMA_signal_11998 ;
    wire new_AGEMA_signal_11999 ;
    wire new_AGEMA_signal_12000 ;
    wire new_AGEMA_signal_12001 ;
    wire new_AGEMA_signal_12002 ;
    wire new_AGEMA_signal_12003 ;
    wire new_AGEMA_signal_12004 ;
    wire new_AGEMA_signal_12005 ;
    wire new_AGEMA_signal_12006 ;
    wire new_AGEMA_signal_12007 ;
    wire new_AGEMA_signal_12008 ;
    wire new_AGEMA_signal_12009 ;
    wire new_AGEMA_signal_12010 ;
    wire new_AGEMA_signal_12011 ;
    wire new_AGEMA_signal_12012 ;
    wire new_AGEMA_signal_12013 ;
    wire new_AGEMA_signal_12014 ;
    wire new_AGEMA_signal_12015 ;
    wire new_AGEMA_signal_12016 ;
    wire new_AGEMA_signal_12017 ;
    wire new_AGEMA_signal_12018 ;
    wire new_AGEMA_signal_12019 ;
    wire new_AGEMA_signal_12020 ;
    wire new_AGEMA_signal_12021 ;
    wire new_AGEMA_signal_12022 ;
    wire new_AGEMA_signal_12023 ;
    wire new_AGEMA_signal_12024 ;
    wire new_AGEMA_signal_12025 ;
    wire new_AGEMA_signal_12026 ;
    wire new_AGEMA_signal_12027 ;
    wire new_AGEMA_signal_12028 ;
    wire new_AGEMA_signal_12029 ;
    wire new_AGEMA_signal_12030 ;
    wire new_AGEMA_signal_12031 ;
    wire new_AGEMA_signal_12032 ;
    wire new_AGEMA_signal_12033 ;
    wire new_AGEMA_signal_12034 ;
    wire new_AGEMA_signal_12035 ;
    wire new_AGEMA_signal_12036 ;
    wire new_AGEMA_signal_12037 ;
    wire new_AGEMA_signal_12038 ;
    wire new_AGEMA_signal_12039 ;
    wire new_AGEMA_signal_12040 ;
    wire new_AGEMA_signal_12041 ;
    wire new_AGEMA_signal_12042 ;
    wire new_AGEMA_signal_12043 ;
    wire new_AGEMA_signal_12044 ;
    wire new_AGEMA_signal_12045 ;
    wire new_AGEMA_signal_12046 ;
    wire new_AGEMA_signal_12047 ;
    wire new_AGEMA_signal_12048 ;
    wire new_AGEMA_signal_12049 ;
    wire new_AGEMA_signal_12050 ;
    wire new_AGEMA_signal_12051 ;
    wire new_AGEMA_signal_12052 ;
    wire new_AGEMA_signal_12053 ;
    wire new_AGEMA_signal_12054 ;
    wire new_AGEMA_signal_12055 ;
    wire new_AGEMA_signal_12056 ;
    wire new_AGEMA_signal_12057 ;
    wire new_AGEMA_signal_12058 ;
    wire new_AGEMA_signal_12059 ;
    wire new_AGEMA_signal_12060 ;
    wire new_AGEMA_signal_12061 ;
    wire new_AGEMA_signal_12062 ;
    wire new_AGEMA_signal_12063 ;
    wire new_AGEMA_signal_12064 ;
    wire new_AGEMA_signal_12065 ;
    wire new_AGEMA_signal_12066 ;
    wire new_AGEMA_signal_12067 ;
    wire new_AGEMA_signal_12068 ;
    wire new_AGEMA_signal_12069 ;
    wire new_AGEMA_signal_12070 ;
    wire new_AGEMA_signal_12071 ;
    wire new_AGEMA_signal_12072 ;
    wire new_AGEMA_signal_12073 ;
    wire new_AGEMA_signal_12074 ;
    wire new_AGEMA_signal_12075 ;
    wire new_AGEMA_signal_12076 ;
    wire new_AGEMA_signal_12077 ;
    wire new_AGEMA_signal_12078 ;
    wire new_AGEMA_signal_12079 ;
    wire new_AGEMA_signal_12080 ;
    wire new_AGEMA_signal_12081 ;
    wire new_AGEMA_signal_12082 ;
    wire new_AGEMA_signal_12083 ;
    wire new_AGEMA_signal_12084 ;
    wire new_AGEMA_signal_12085 ;
    wire new_AGEMA_signal_12086 ;
    wire new_AGEMA_signal_12087 ;
    wire new_AGEMA_signal_12088 ;
    wire new_AGEMA_signal_12089 ;
    wire new_AGEMA_signal_12090 ;
    wire new_AGEMA_signal_12091 ;
    wire new_AGEMA_signal_12092 ;
    wire new_AGEMA_signal_12093 ;
    wire new_AGEMA_signal_12094 ;
    wire new_AGEMA_signal_12095 ;
    wire new_AGEMA_signal_12096 ;
    wire new_AGEMA_signal_12097 ;
    wire new_AGEMA_signal_12098 ;
    wire new_AGEMA_signal_12099 ;
    wire new_AGEMA_signal_12100 ;
    wire new_AGEMA_signal_12101 ;
    wire new_AGEMA_signal_12102 ;
    wire new_AGEMA_signal_12103 ;
    wire new_AGEMA_signal_12104 ;
    wire new_AGEMA_signal_12105 ;
    wire new_AGEMA_signal_12106 ;
    wire new_AGEMA_signal_12107 ;
    wire new_AGEMA_signal_12108 ;
    wire new_AGEMA_signal_12109 ;
    wire new_AGEMA_signal_12110 ;
    wire new_AGEMA_signal_12111 ;
    wire new_AGEMA_signal_12112 ;
    wire new_AGEMA_signal_12113 ;
    wire new_AGEMA_signal_12114 ;
    wire new_AGEMA_signal_12115 ;
    wire new_AGEMA_signal_12116 ;
    wire new_AGEMA_signal_12117 ;
    wire new_AGEMA_signal_12118 ;
    wire new_AGEMA_signal_12119 ;
    wire new_AGEMA_signal_12120 ;
    wire new_AGEMA_signal_12121 ;
    wire new_AGEMA_signal_12122 ;
    wire new_AGEMA_signal_12123 ;
    wire new_AGEMA_signal_12124 ;
    wire new_AGEMA_signal_12125 ;
    wire new_AGEMA_signal_12126 ;
    wire new_AGEMA_signal_12127 ;
    wire new_AGEMA_signal_12128 ;
    wire new_AGEMA_signal_12129 ;
    wire new_AGEMA_signal_12130 ;
    wire new_AGEMA_signal_12131 ;
    wire new_AGEMA_signal_12132 ;
    wire new_AGEMA_signal_12133 ;
    wire new_AGEMA_signal_12134 ;
    wire new_AGEMA_signal_12135 ;
    wire new_AGEMA_signal_12136 ;
    wire new_AGEMA_signal_12137 ;
    wire new_AGEMA_signal_12138 ;
    wire new_AGEMA_signal_12139 ;
    wire new_AGEMA_signal_12140 ;
    wire new_AGEMA_signal_12141 ;
    wire new_AGEMA_signal_12142 ;
    wire new_AGEMA_signal_12143 ;
    wire new_AGEMA_signal_12144 ;
    wire new_AGEMA_signal_12145 ;
    wire new_AGEMA_signal_12146 ;
    wire new_AGEMA_signal_12147 ;
    wire new_AGEMA_signal_12148 ;
    wire new_AGEMA_signal_12149 ;
    wire new_AGEMA_signal_12150 ;
    wire new_AGEMA_signal_12151 ;
    wire new_AGEMA_signal_12152 ;
    wire new_AGEMA_signal_12153 ;
    wire new_AGEMA_signal_12154 ;
    wire new_AGEMA_signal_12155 ;
    wire new_AGEMA_signal_12156 ;
    wire new_AGEMA_signal_12157 ;
    wire new_AGEMA_signal_12158 ;
    wire new_AGEMA_signal_12159 ;
    wire new_AGEMA_signal_12160 ;
    wire new_AGEMA_signal_12161 ;
    wire new_AGEMA_signal_12162 ;
    wire new_AGEMA_signal_12163 ;
    wire new_AGEMA_signal_12164 ;
    wire new_AGEMA_signal_12165 ;
    wire new_AGEMA_signal_12166 ;
    wire new_AGEMA_signal_12167 ;
    wire new_AGEMA_signal_12168 ;
    wire new_AGEMA_signal_12169 ;
    wire new_AGEMA_signal_12170 ;
    wire new_AGEMA_signal_12171 ;
    wire new_AGEMA_signal_12172 ;
    wire new_AGEMA_signal_12173 ;
    wire new_AGEMA_signal_12174 ;
    wire new_AGEMA_signal_12175 ;
    wire new_AGEMA_signal_12176 ;
    wire new_AGEMA_signal_12177 ;
    wire new_AGEMA_signal_12178 ;
    wire new_AGEMA_signal_12179 ;
    wire new_AGEMA_signal_12180 ;
    wire new_AGEMA_signal_12181 ;
    wire new_AGEMA_signal_12182 ;
    wire new_AGEMA_signal_12183 ;
    wire new_AGEMA_signal_12184 ;
    wire new_AGEMA_signal_12185 ;
    wire new_AGEMA_signal_12186 ;
    wire new_AGEMA_signal_12187 ;
    wire new_AGEMA_signal_12188 ;
    wire new_AGEMA_signal_12189 ;
    wire new_AGEMA_signal_12190 ;
    wire new_AGEMA_signal_12191 ;
    wire new_AGEMA_signal_12192 ;
    wire new_AGEMA_signal_12193 ;
    wire new_AGEMA_signal_12194 ;
    wire new_AGEMA_signal_12195 ;
    wire new_AGEMA_signal_12196 ;
    wire new_AGEMA_signal_12197 ;
    wire new_AGEMA_signal_12198 ;
    wire new_AGEMA_signal_12199 ;
    wire new_AGEMA_signal_12200 ;
    wire new_AGEMA_signal_12201 ;
    wire new_AGEMA_signal_12202 ;
    wire new_AGEMA_signal_12203 ;
    wire new_AGEMA_signal_12204 ;
    wire new_AGEMA_signal_12205 ;
    wire new_AGEMA_signal_12206 ;
    wire new_AGEMA_signal_12207 ;
    wire new_AGEMA_signal_12208 ;
    wire new_AGEMA_signal_12209 ;
    wire new_AGEMA_signal_12210 ;
    wire new_AGEMA_signal_12211 ;
    wire new_AGEMA_signal_12212 ;
    wire new_AGEMA_signal_12213 ;
    wire new_AGEMA_signal_12214 ;
    wire new_AGEMA_signal_12215 ;
    wire new_AGEMA_signal_12216 ;
    wire new_AGEMA_signal_12217 ;
    wire new_AGEMA_signal_12218 ;
    wire new_AGEMA_signal_12219 ;
    wire new_AGEMA_signal_12220 ;
    wire new_AGEMA_signal_12221 ;
    wire new_AGEMA_signal_12222 ;
    wire new_AGEMA_signal_12223 ;
    wire new_AGEMA_signal_12224 ;
    wire new_AGEMA_signal_12225 ;
    wire new_AGEMA_signal_12226 ;
    wire new_AGEMA_signal_12227 ;
    wire new_AGEMA_signal_12228 ;
    wire new_AGEMA_signal_12229 ;
    wire new_AGEMA_signal_12230 ;
    wire new_AGEMA_signal_12231 ;
    wire new_AGEMA_signal_12232 ;
    wire new_AGEMA_signal_12233 ;
    wire new_AGEMA_signal_12234 ;
    wire new_AGEMA_signal_12235 ;
    wire new_AGEMA_signal_12236 ;
    wire new_AGEMA_signal_12237 ;
    wire new_AGEMA_signal_12238 ;
    wire new_AGEMA_signal_12239 ;
    wire new_AGEMA_signal_12240 ;
    wire new_AGEMA_signal_12241 ;
    wire new_AGEMA_signal_12242 ;
    wire new_AGEMA_signal_12243 ;
    wire new_AGEMA_signal_12244 ;
    wire new_AGEMA_signal_12245 ;
    wire new_AGEMA_signal_12246 ;
    wire new_AGEMA_signal_12247 ;
    wire new_AGEMA_signal_12248 ;
    wire new_AGEMA_signal_12249 ;
    wire new_AGEMA_signal_12250 ;
    wire new_AGEMA_signal_12251 ;
    wire new_AGEMA_signal_12252 ;
    wire new_AGEMA_signal_12253 ;
    wire new_AGEMA_signal_12254 ;
    wire new_AGEMA_signal_12255 ;
    wire new_AGEMA_signal_12256 ;
    wire new_AGEMA_signal_12257 ;
    wire new_AGEMA_signal_12258 ;
    wire new_AGEMA_signal_12259 ;
    wire new_AGEMA_signal_12260 ;
    wire new_AGEMA_signal_12261 ;
    wire new_AGEMA_signal_12262 ;
    wire new_AGEMA_signal_12263 ;
    wire new_AGEMA_signal_12264 ;
    wire new_AGEMA_signal_12265 ;
    wire new_AGEMA_signal_12266 ;
    wire new_AGEMA_signal_12267 ;
    wire new_AGEMA_signal_12268 ;
    wire new_AGEMA_signal_12269 ;
    wire new_AGEMA_signal_12270 ;
    wire new_AGEMA_signal_12271 ;
    wire new_AGEMA_signal_12272 ;
    wire new_AGEMA_signal_12273 ;
    wire new_AGEMA_signal_12274 ;
    wire new_AGEMA_signal_12275 ;
    wire new_AGEMA_signal_12276 ;
    wire new_AGEMA_signal_12277 ;
    wire new_AGEMA_signal_12278 ;
    wire new_AGEMA_signal_12279 ;
    wire new_AGEMA_signal_12280 ;
    wire new_AGEMA_signal_12281 ;
    wire new_AGEMA_signal_12282 ;
    wire new_AGEMA_signal_12283 ;
    wire new_AGEMA_signal_12284 ;
    wire new_AGEMA_signal_12285 ;
    wire new_AGEMA_signal_12286 ;
    wire new_AGEMA_signal_12287 ;
    wire new_AGEMA_signal_12288 ;
    wire new_AGEMA_signal_12289 ;
    wire new_AGEMA_signal_12290 ;
    wire new_AGEMA_signal_12291 ;
    wire new_AGEMA_signal_12292 ;
    wire new_AGEMA_signal_12293 ;
    wire new_AGEMA_signal_12294 ;
    wire new_AGEMA_signal_12295 ;
    wire new_AGEMA_signal_12296 ;
    wire new_AGEMA_signal_12297 ;
    wire new_AGEMA_signal_12298 ;
    wire new_AGEMA_signal_12299 ;
    wire new_AGEMA_signal_12300 ;
    wire new_AGEMA_signal_12301 ;
    wire new_AGEMA_signal_12302 ;
    wire new_AGEMA_signal_12303 ;
    wire new_AGEMA_signal_12304 ;
    wire new_AGEMA_signal_12305 ;
    wire new_AGEMA_signal_12306 ;
    wire new_AGEMA_signal_12307 ;
    wire new_AGEMA_signal_12308 ;
    wire new_AGEMA_signal_12309 ;
    wire new_AGEMA_signal_12310 ;
    wire new_AGEMA_signal_12311 ;
    wire new_AGEMA_signal_12312 ;
    wire new_AGEMA_signal_12313 ;
    wire new_AGEMA_signal_12314 ;
    wire new_AGEMA_signal_12315 ;
    wire new_AGEMA_signal_12316 ;
    wire new_AGEMA_signal_12317 ;
    wire new_AGEMA_signal_12318 ;
    wire new_AGEMA_signal_12319 ;
    wire new_AGEMA_signal_12320 ;
    wire new_AGEMA_signal_12321 ;
    wire new_AGEMA_signal_12322 ;
    wire new_AGEMA_signal_12323 ;
    wire new_AGEMA_signal_12324 ;
    wire new_AGEMA_signal_12325 ;
    wire new_AGEMA_signal_12326 ;
    wire new_AGEMA_signal_12327 ;
    wire new_AGEMA_signal_12328 ;
    wire new_AGEMA_signal_12329 ;
    wire new_AGEMA_signal_12330 ;
    wire new_AGEMA_signal_12331 ;
    wire new_AGEMA_signal_12332 ;
    wire new_AGEMA_signal_12333 ;
    wire new_AGEMA_signal_12334 ;
    wire new_AGEMA_signal_12335 ;
    wire new_AGEMA_signal_12336 ;
    wire new_AGEMA_signal_12337 ;
    wire new_AGEMA_signal_12338 ;
    wire new_AGEMA_signal_12339 ;
    wire new_AGEMA_signal_12340 ;
    wire new_AGEMA_signal_12341 ;
    wire new_AGEMA_signal_12342 ;
    wire new_AGEMA_signal_12343 ;
    wire new_AGEMA_signal_12344 ;
    wire new_AGEMA_signal_12345 ;
    wire new_AGEMA_signal_12346 ;
    wire new_AGEMA_signal_12347 ;
    wire new_AGEMA_signal_12348 ;
    wire new_AGEMA_signal_12349 ;
    wire new_AGEMA_signal_12350 ;
    wire new_AGEMA_signal_12351 ;
    wire new_AGEMA_signal_12352 ;
    wire new_AGEMA_signal_12353 ;
    wire new_AGEMA_signal_12354 ;
    wire new_AGEMA_signal_12355 ;
    wire new_AGEMA_signal_12356 ;
    wire new_AGEMA_signal_12357 ;
    wire new_AGEMA_signal_12358 ;
    wire new_AGEMA_signal_12359 ;
    wire new_AGEMA_signal_12360 ;
    wire new_AGEMA_signal_12361 ;
    wire new_AGEMA_signal_12362 ;
    wire new_AGEMA_signal_12363 ;
    wire new_AGEMA_signal_12364 ;
    wire new_AGEMA_signal_12365 ;
    wire new_AGEMA_signal_12366 ;
    wire new_AGEMA_signal_12367 ;
    wire new_AGEMA_signal_12368 ;
    wire new_AGEMA_signal_12369 ;
    wire new_AGEMA_signal_12370 ;
    wire new_AGEMA_signal_12371 ;
    wire new_AGEMA_signal_12372 ;
    wire new_AGEMA_signal_12373 ;
    wire new_AGEMA_signal_12374 ;
    wire new_AGEMA_signal_12375 ;
    wire new_AGEMA_signal_12376 ;
    wire new_AGEMA_signal_12377 ;
    wire new_AGEMA_signal_12378 ;
    wire new_AGEMA_signal_12379 ;
    wire new_AGEMA_signal_12380 ;
    wire new_AGEMA_signal_12381 ;
    wire new_AGEMA_signal_12382 ;
    wire new_AGEMA_signal_12383 ;
    wire new_AGEMA_signal_12384 ;
    wire new_AGEMA_signal_12385 ;
    wire new_AGEMA_signal_12386 ;
    wire new_AGEMA_signal_12387 ;
    wire new_AGEMA_signal_12388 ;
    wire new_AGEMA_signal_12389 ;
    wire new_AGEMA_signal_12390 ;
    wire new_AGEMA_signal_12391 ;
    wire new_AGEMA_signal_12392 ;
    wire new_AGEMA_signal_12393 ;
    wire new_AGEMA_signal_12394 ;
    wire new_AGEMA_signal_12395 ;
    wire new_AGEMA_signal_12396 ;
    wire new_AGEMA_signal_12397 ;
    wire new_AGEMA_signal_12398 ;
    wire new_AGEMA_signal_12399 ;
    wire new_AGEMA_signal_12400 ;
    wire new_AGEMA_signal_12401 ;
    wire new_AGEMA_signal_12402 ;
    wire new_AGEMA_signal_12403 ;
    wire new_AGEMA_signal_12404 ;
    wire new_AGEMA_signal_12405 ;
    wire new_AGEMA_signal_12406 ;
    wire new_AGEMA_signal_12407 ;
    wire new_AGEMA_signal_12408 ;
    wire new_AGEMA_signal_12409 ;
    wire new_AGEMA_signal_12410 ;
    wire new_AGEMA_signal_12411 ;
    wire new_AGEMA_signal_12412 ;
    wire new_AGEMA_signal_12413 ;
    wire new_AGEMA_signal_12414 ;
    wire new_AGEMA_signal_12415 ;
    wire new_AGEMA_signal_12416 ;
    wire new_AGEMA_signal_12417 ;
    wire new_AGEMA_signal_12418 ;
    wire new_AGEMA_signal_12419 ;
    wire new_AGEMA_signal_12420 ;
    wire new_AGEMA_signal_12421 ;
    wire new_AGEMA_signal_12422 ;
    wire new_AGEMA_signal_12423 ;
    wire new_AGEMA_signal_12424 ;
    wire new_AGEMA_signal_12425 ;
    wire new_AGEMA_signal_12426 ;
    wire new_AGEMA_signal_12427 ;
    wire new_AGEMA_signal_12428 ;
    wire new_AGEMA_signal_12429 ;
    wire new_AGEMA_signal_12430 ;
    wire new_AGEMA_signal_12431 ;
    wire new_AGEMA_signal_12432 ;
    wire new_AGEMA_signal_12433 ;
    wire new_AGEMA_signal_12434 ;
    wire new_AGEMA_signal_12435 ;
    wire new_AGEMA_signal_12436 ;
    wire new_AGEMA_signal_12437 ;
    wire new_AGEMA_signal_12438 ;
    wire new_AGEMA_signal_12439 ;
    wire new_AGEMA_signal_12440 ;
    wire new_AGEMA_signal_12441 ;
    wire new_AGEMA_signal_12442 ;
    wire new_AGEMA_signal_12443 ;
    wire new_AGEMA_signal_12444 ;
    wire new_AGEMA_signal_12445 ;
    wire new_AGEMA_signal_12446 ;
    wire new_AGEMA_signal_12447 ;
    wire new_AGEMA_signal_12448 ;
    wire new_AGEMA_signal_12449 ;
    wire new_AGEMA_signal_12450 ;
    wire new_AGEMA_signal_12451 ;
    wire new_AGEMA_signal_12452 ;
    wire new_AGEMA_signal_12453 ;
    wire new_AGEMA_signal_12454 ;
    wire new_AGEMA_signal_12455 ;
    wire new_AGEMA_signal_12456 ;
    wire new_AGEMA_signal_12457 ;
    wire new_AGEMA_signal_12458 ;
    wire new_AGEMA_signal_12459 ;
    wire new_AGEMA_signal_12460 ;
    wire new_AGEMA_signal_12461 ;
    wire new_AGEMA_signal_12462 ;
    wire new_AGEMA_signal_12463 ;
    wire new_AGEMA_signal_12464 ;
    wire new_AGEMA_signal_12465 ;
    wire new_AGEMA_signal_12466 ;
    wire new_AGEMA_signal_12467 ;
    wire new_AGEMA_signal_12468 ;
    wire new_AGEMA_signal_12469 ;
    wire new_AGEMA_signal_12470 ;
    wire new_AGEMA_signal_12471 ;
    wire new_AGEMA_signal_12472 ;
    wire new_AGEMA_signal_12473 ;
    wire new_AGEMA_signal_12474 ;
    wire new_AGEMA_signal_12475 ;
    wire new_AGEMA_signal_12476 ;
    wire new_AGEMA_signal_12477 ;
    wire new_AGEMA_signal_12478 ;
    wire new_AGEMA_signal_12479 ;
    wire new_AGEMA_signal_12480 ;
    wire new_AGEMA_signal_12481 ;
    wire new_AGEMA_signal_12482 ;
    wire new_AGEMA_signal_12483 ;
    wire new_AGEMA_signal_12484 ;
    wire new_AGEMA_signal_12485 ;
    wire new_AGEMA_signal_12486 ;
    wire new_AGEMA_signal_12487 ;
    wire new_AGEMA_signal_12488 ;
    wire new_AGEMA_signal_12489 ;
    wire new_AGEMA_signal_12490 ;
    wire new_AGEMA_signal_12491 ;
    wire new_AGEMA_signal_12492 ;
    wire new_AGEMA_signal_12493 ;
    wire new_AGEMA_signal_12494 ;
    wire new_AGEMA_signal_12495 ;
    wire new_AGEMA_signal_12496 ;
    wire new_AGEMA_signal_12497 ;
    wire new_AGEMA_signal_12498 ;
    wire new_AGEMA_signal_12499 ;
    wire new_AGEMA_signal_12500 ;
    wire new_AGEMA_signal_12501 ;
    wire new_AGEMA_signal_12502 ;
    wire new_AGEMA_signal_12503 ;
    wire new_AGEMA_signal_12504 ;
    wire new_AGEMA_signal_12505 ;
    wire new_AGEMA_signal_12506 ;
    wire new_AGEMA_signal_12507 ;
    wire new_AGEMA_signal_12508 ;
    wire new_AGEMA_signal_12509 ;
    wire new_AGEMA_signal_12510 ;
    wire new_AGEMA_signal_12511 ;
    wire new_AGEMA_signal_12512 ;
    wire new_AGEMA_signal_12513 ;
    wire new_AGEMA_signal_12514 ;
    wire new_AGEMA_signal_12515 ;
    wire new_AGEMA_signal_12516 ;
    wire new_AGEMA_signal_12517 ;
    wire new_AGEMA_signal_12518 ;
    wire new_AGEMA_signal_12519 ;
    wire new_AGEMA_signal_12520 ;
    wire new_AGEMA_signal_12521 ;
    wire new_AGEMA_signal_12522 ;
    wire new_AGEMA_signal_12523 ;
    wire new_AGEMA_signal_12524 ;
    wire new_AGEMA_signal_12525 ;
    wire new_AGEMA_signal_12526 ;
    wire new_AGEMA_signal_12527 ;
    wire new_AGEMA_signal_12528 ;
    wire new_AGEMA_signal_12529 ;
    wire new_AGEMA_signal_12530 ;
    wire new_AGEMA_signal_12531 ;
    wire new_AGEMA_signal_12532 ;
    wire new_AGEMA_signal_12533 ;
    wire new_AGEMA_signal_12534 ;
    wire new_AGEMA_signal_12535 ;
    wire new_AGEMA_signal_12536 ;
    wire new_AGEMA_signal_12537 ;
    wire new_AGEMA_signal_12538 ;
    wire new_AGEMA_signal_12539 ;
    wire new_AGEMA_signal_12540 ;
    wire new_AGEMA_signal_12541 ;
    wire new_AGEMA_signal_12542 ;
    wire new_AGEMA_signal_12543 ;
    wire new_AGEMA_signal_12544 ;
    wire new_AGEMA_signal_12545 ;
    wire new_AGEMA_signal_12546 ;
    wire new_AGEMA_signal_12547 ;
    wire new_AGEMA_signal_12548 ;
    wire new_AGEMA_signal_12549 ;
    wire new_AGEMA_signal_12550 ;
    wire new_AGEMA_signal_12551 ;
    wire new_AGEMA_signal_12552 ;
    wire new_AGEMA_signal_12553 ;
    wire new_AGEMA_signal_12554 ;
    wire new_AGEMA_signal_12555 ;
    wire new_AGEMA_signal_12556 ;
    wire new_AGEMA_signal_12557 ;
    wire new_AGEMA_signal_12558 ;
    wire new_AGEMA_signal_12559 ;
    wire new_AGEMA_signal_12560 ;
    wire new_AGEMA_signal_12561 ;
    wire new_AGEMA_signal_12562 ;
    wire new_AGEMA_signal_12563 ;
    wire new_AGEMA_signal_12564 ;
    wire new_AGEMA_signal_12565 ;
    wire new_AGEMA_signal_12566 ;
    wire new_AGEMA_signal_12567 ;
    wire new_AGEMA_signal_12568 ;
    wire new_AGEMA_signal_12569 ;
    wire new_AGEMA_signal_12570 ;
    wire new_AGEMA_signal_12571 ;
    wire new_AGEMA_signal_12572 ;
    wire new_AGEMA_signal_12573 ;
    wire new_AGEMA_signal_12574 ;
    wire new_AGEMA_signal_12575 ;
    wire new_AGEMA_signal_12576 ;
    wire new_AGEMA_signal_12577 ;
    wire new_AGEMA_signal_12578 ;
    wire new_AGEMA_signal_12579 ;
    wire new_AGEMA_signal_12580 ;
    wire new_AGEMA_signal_12581 ;
    wire new_AGEMA_signal_12582 ;
    wire new_AGEMA_signal_12583 ;
    wire new_AGEMA_signal_12584 ;
    wire new_AGEMA_signal_12585 ;
    wire new_AGEMA_signal_12586 ;
    wire new_AGEMA_signal_12587 ;
    wire new_AGEMA_signal_12588 ;
    wire new_AGEMA_signal_12589 ;
    wire new_AGEMA_signal_12590 ;
    wire new_AGEMA_signal_12591 ;
    wire new_AGEMA_signal_12592 ;
    wire new_AGEMA_signal_12593 ;
    wire new_AGEMA_signal_12594 ;
    wire new_AGEMA_signal_12595 ;
    wire new_AGEMA_signal_12596 ;
    wire new_AGEMA_signal_12597 ;
    wire new_AGEMA_signal_12598 ;
    wire new_AGEMA_signal_12599 ;
    wire new_AGEMA_signal_12600 ;
    wire new_AGEMA_signal_12601 ;
    wire new_AGEMA_signal_12602 ;
    wire new_AGEMA_signal_12603 ;
    wire new_AGEMA_signal_12604 ;
    wire new_AGEMA_signal_12605 ;
    wire new_AGEMA_signal_12606 ;
    wire new_AGEMA_signal_12607 ;
    wire new_AGEMA_signal_12608 ;
    wire new_AGEMA_signal_12609 ;
    wire new_AGEMA_signal_12610 ;
    wire new_AGEMA_signal_12611 ;
    wire new_AGEMA_signal_12612 ;
    wire new_AGEMA_signal_12613 ;
    wire new_AGEMA_signal_12614 ;
    wire new_AGEMA_signal_12615 ;
    wire new_AGEMA_signal_12616 ;
    wire new_AGEMA_signal_12617 ;
    wire new_AGEMA_signal_12618 ;
    wire new_AGEMA_signal_12619 ;
    wire new_AGEMA_signal_12620 ;
    wire new_AGEMA_signal_12621 ;
    wire new_AGEMA_signal_12622 ;
    wire new_AGEMA_signal_12623 ;
    wire new_AGEMA_signal_12624 ;
    wire new_AGEMA_signal_12625 ;
    wire new_AGEMA_signal_12626 ;
    wire new_AGEMA_signal_12627 ;
    wire new_AGEMA_signal_12628 ;
    wire new_AGEMA_signal_12629 ;
    wire new_AGEMA_signal_12630 ;
    wire new_AGEMA_signal_12631 ;
    wire new_AGEMA_signal_12632 ;
    wire new_AGEMA_signal_12633 ;
    wire new_AGEMA_signal_12634 ;
    wire new_AGEMA_signal_12635 ;
    wire new_AGEMA_signal_12636 ;
    wire new_AGEMA_signal_12637 ;
    wire new_AGEMA_signal_12638 ;
    wire new_AGEMA_signal_12639 ;
    wire new_AGEMA_signal_12640 ;
    wire new_AGEMA_signal_12641 ;
    wire new_AGEMA_signal_12642 ;
    wire new_AGEMA_signal_12643 ;
    wire new_AGEMA_signal_12644 ;
    wire new_AGEMA_signal_12645 ;
    wire new_AGEMA_signal_12646 ;
    wire new_AGEMA_signal_12647 ;
    wire new_AGEMA_signal_12648 ;
    wire new_AGEMA_signal_12649 ;
    wire new_AGEMA_signal_12650 ;
    wire new_AGEMA_signal_12651 ;
    wire new_AGEMA_signal_12652 ;
    wire new_AGEMA_signal_12653 ;
    wire new_AGEMA_signal_12654 ;
    wire new_AGEMA_signal_12655 ;
    wire new_AGEMA_signal_12656 ;
    wire new_AGEMA_signal_12657 ;
    wire new_AGEMA_signal_12658 ;
    wire new_AGEMA_signal_12659 ;
    wire new_AGEMA_signal_12660 ;
    wire new_AGEMA_signal_12661 ;
    wire new_AGEMA_signal_12662 ;
    wire new_AGEMA_signal_12663 ;
    wire new_AGEMA_signal_12664 ;
    wire new_AGEMA_signal_12665 ;
    wire new_AGEMA_signal_12666 ;
    wire new_AGEMA_signal_12667 ;
    wire new_AGEMA_signal_12668 ;
    wire new_AGEMA_signal_12669 ;
    wire new_AGEMA_signal_12670 ;
    wire new_AGEMA_signal_12671 ;
    wire new_AGEMA_signal_12672 ;
    wire new_AGEMA_signal_12673 ;
    wire new_AGEMA_signal_12674 ;
    wire new_AGEMA_signal_12675 ;
    wire new_AGEMA_signal_12676 ;
    wire new_AGEMA_signal_12677 ;
    wire new_AGEMA_signal_12678 ;
    wire new_AGEMA_signal_12679 ;
    wire new_AGEMA_signal_12680 ;
    wire new_AGEMA_signal_12681 ;
    wire new_AGEMA_signal_12682 ;
    wire new_AGEMA_signal_12683 ;
    wire new_AGEMA_signal_12684 ;
    wire new_AGEMA_signal_12685 ;
    wire new_AGEMA_signal_12686 ;
    wire new_AGEMA_signal_12687 ;
    wire new_AGEMA_signal_12688 ;
    wire new_AGEMA_signal_12689 ;
    wire new_AGEMA_signal_12690 ;
    wire new_AGEMA_signal_12691 ;
    wire new_AGEMA_signal_12692 ;
    wire new_AGEMA_signal_12693 ;
    wire new_AGEMA_signal_12694 ;
    wire new_AGEMA_signal_12695 ;
    wire new_AGEMA_signal_12696 ;
    wire new_AGEMA_signal_12697 ;
    wire new_AGEMA_signal_12698 ;
    wire new_AGEMA_signal_12699 ;
    wire new_AGEMA_signal_12700 ;
    wire new_AGEMA_signal_12701 ;
    wire new_AGEMA_signal_12702 ;
    wire new_AGEMA_signal_12703 ;
    wire new_AGEMA_signal_12704 ;
    wire new_AGEMA_signal_12705 ;
    wire new_AGEMA_signal_12706 ;
    wire new_AGEMA_signal_12707 ;
    wire new_AGEMA_signal_12708 ;
    wire new_AGEMA_signal_12709 ;
    wire new_AGEMA_signal_12710 ;
    wire new_AGEMA_signal_12711 ;
    wire new_AGEMA_signal_12712 ;
    wire new_AGEMA_signal_12713 ;
    wire new_AGEMA_signal_12714 ;
    wire new_AGEMA_signal_12715 ;
    wire new_AGEMA_signal_12716 ;
    wire new_AGEMA_signal_12717 ;
    wire new_AGEMA_signal_12718 ;
    wire new_AGEMA_signal_12719 ;
    wire new_AGEMA_signal_12720 ;
    wire new_AGEMA_signal_12721 ;
    wire new_AGEMA_signal_12722 ;
    wire new_AGEMA_signal_12723 ;
    wire new_AGEMA_signal_12724 ;
    wire new_AGEMA_signal_12725 ;
    wire new_AGEMA_signal_12726 ;
    wire new_AGEMA_signal_12727 ;
    wire new_AGEMA_signal_12728 ;
    wire new_AGEMA_signal_12729 ;
    wire new_AGEMA_signal_12730 ;
    wire new_AGEMA_signal_12731 ;
    wire new_AGEMA_signal_12732 ;
    wire new_AGEMA_signal_12733 ;
    wire new_AGEMA_signal_12734 ;
    wire new_AGEMA_signal_12735 ;
    wire new_AGEMA_signal_12736 ;
    wire new_AGEMA_signal_12737 ;
    wire new_AGEMA_signal_12738 ;
    wire new_AGEMA_signal_12739 ;
    wire new_AGEMA_signal_12740 ;
    wire new_AGEMA_signal_12741 ;
    wire new_AGEMA_signal_12742 ;
    wire new_AGEMA_signal_12743 ;
    wire new_AGEMA_signal_12744 ;
    wire new_AGEMA_signal_12745 ;
    wire new_AGEMA_signal_12746 ;
    wire new_AGEMA_signal_12747 ;
    wire new_AGEMA_signal_12748 ;
    wire new_AGEMA_signal_12749 ;
    wire new_AGEMA_signal_12750 ;
    wire new_AGEMA_signal_12751 ;
    wire new_AGEMA_signal_12752 ;
    wire new_AGEMA_signal_12753 ;
    wire new_AGEMA_signal_12754 ;
    wire new_AGEMA_signal_12755 ;
    wire new_AGEMA_signal_12756 ;
    wire new_AGEMA_signal_12757 ;
    wire new_AGEMA_signal_12758 ;
    wire new_AGEMA_signal_12759 ;
    wire new_AGEMA_signal_12760 ;
    wire new_AGEMA_signal_12761 ;
    wire new_AGEMA_signal_12762 ;
    wire new_AGEMA_signal_12763 ;
    wire new_AGEMA_signal_12764 ;
    wire new_AGEMA_signal_12765 ;
    wire new_AGEMA_signal_12766 ;
    wire new_AGEMA_signal_12767 ;
    wire new_AGEMA_signal_12768 ;
    wire new_AGEMA_signal_12769 ;
    wire new_AGEMA_signal_12770 ;
    wire new_AGEMA_signal_12771 ;
    wire new_AGEMA_signal_12772 ;
    wire new_AGEMA_signal_12773 ;
    wire new_AGEMA_signal_12774 ;
    wire new_AGEMA_signal_12775 ;
    wire new_AGEMA_signal_12776 ;
    wire new_AGEMA_signal_12777 ;
    wire new_AGEMA_signal_12778 ;
    wire new_AGEMA_signal_12779 ;
    wire new_AGEMA_signal_12780 ;
    wire new_AGEMA_signal_12781 ;
    wire new_AGEMA_signal_12782 ;
    wire new_AGEMA_signal_12783 ;
    wire new_AGEMA_signal_12784 ;
    wire new_AGEMA_signal_12785 ;
    wire new_AGEMA_signal_12786 ;
    wire new_AGEMA_signal_12787 ;
    wire new_AGEMA_signal_12788 ;
    wire new_AGEMA_signal_12789 ;
    wire new_AGEMA_signal_12790 ;
    wire new_AGEMA_signal_12791 ;
    wire new_AGEMA_signal_12792 ;
    wire new_AGEMA_signal_12793 ;
    wire new_AGEMA_signal_12794 ;
    wire new_AGEMA_signal_12795 ;
    wire new_AGEMA_signal_12796 ;
    wire new_AGEMA_signal_12797 ;
    wire new_AGEMA_signal_12798 ;
    wire new_AGEMA_signal_12799 ;
    wire new_AGEMA_signal_12800 ;
    wire new_AGEMA_signal_12801 ;
    wire new_AGEMA_signal_12802 ;
    wire new_AGEMA_signal_12803 ;
    wire new_AGEMA_signal_12804 ;
    wire new_AGEMA_signal_12805 ;
    wire new_AGEMA_signal_12806 ;
    wire new_AGEMA_signal_12807 ;
    wire new_AGEMA_signal_12808 ;
    wire new_AGEMA_signal_12809 ;
    wire new_AGEMA_signal_12810 ;
    wire new_AGEMA_signal_12811 ;
    wire new_AGEMA_signal_12812 ;
    wire new_AGEMA_signal_12813 ;
    wire new_AGEMA_signal_12814 ;
    wire new_AGEMA_signal_12815 ;
    wire new_AGEMA_signal_12816 ;
    wire new_AGEMA_signal_12817 ;
    wire new_AGEMA_signal_12818 ;
    wire new_AGEMA_signal_12819 ;
    wire new_AGEMA_signal_12820 ;
    wire new_AGEMA_signal_12821 ;
    wire new_AGEMA_signal_12822 ;
    wire new_AGEMA_signal_12823 ;
    wire new_AGEMA_signal_12824 ;
    wire new_AGEMA_signal_12825 ;
    wire new_AGEMA_signal_12826 ;
    wire new_AGEMA_signal_12827 ;
    wire new_AGEMA_signal_12828 ;
    wire new_AGEMA_signal_12829 ;
    wire new_AGEMA_signal_12830 ;
    wire new_AGEMA_signal_12831 ;
    wire new_AGEMA_signal_12832 ;
    wire new_AGEMA_signal_12833 ;
    wire new_AGEMA_signal_12834 ;
    wire new_AGEMA_signal_12835 ;
    wire new_AGEMA_signal_12836 ;
    wire new_AGEMA_signal_12837 ;
    wire new_AGEMA_signal_12838 ;
    wire new_AGEMA_signal_12839 ;
    wire new_AGEMA_signal_12840 ;
    wire new_AGEMA_signal_12841 ;
    wire new_AGEMA_signal_12842 ;
    wire new_AGEMA_signal_12843 ;
    wire new_AGEMA_signal_12844 ;
    wire new_AGEMA_signal_12845 ;
    wire new_AGEMA_signal_12846 ;
    wire new_AGEMA_signal_12847 ;
    wire new_AGEMA_signal_12848 ;
    wire new_AGEMA_signal_12849 ;
    wire new_AGEMA_signal_12850 ;
    wire new_AGEMA_signal_12851 ;
    wire new_AGEMA_signal_12852 ;
    wire new_AGEMA_signal_12853 ;
    wire new_AGEMA_signal_12854 ;
    wire new_AGEMA_signal_12855 ;
    wire new_AGEMA_signal_12856 ;
    wire new_AGEMA_signal_12857 ;
    wire new_AGEMA_signal_12858 ;
    wire new_AGEMA_signal_12859 ;
    wire new_AGEMA_signal_12860 ;
    wire new_AGEMA_signal_12861 ;
    wire new_AGEMA_signal_12862 ;
    wire new_AGEMA_signal_12863 ;
    wire new_AGEMA_signal_12864 ;
    wire new_AGEMA_signal_12865 ;
    wire new_AGEMA_signal_12866 ;
    wire new_AGEMA_signal_12867 ;
    wire new_AGEMA_signal_12868 ;
    wire new_AGEMA_signal_12869 ;
    wire new_AGEMA_signal_12870 ;
    wire new_AGEMA_signal_12871 ;
    wire new_AGEMA_signal_12872 ;
    wire new_AGEMA_signal_12873 ;
    wire new_AGEMA_signal_12874 ;
    wire new_AGEMA_signal_12875 ;
    wire new_AGEMA_signal_12876 ;
    wire new_AGEMA_signal_12877 ;
    wire new_AGEMA_signal_12878 ;
    wire new_AGEMA_signal_12879 ;
    wire new_AGEMA_signal_12880 ;
    wire new_AGEMA_signal_12881 ;
    wire new_AGEMA_signal_12882 ;
    wire new_AGEMA_signal_12883 ;
    wire new_AGEMA_signal_12884 ;
    wire new_AGEMA_signal_12885 ;
    wire new_AGEMA_signal_12886 ;
    wire new_AGEMA_signal_12887 ;
    wire new_AGEMA_signal_12888 ;
    wire new_AGEMA_signal_12889 ;
    wire new_AGEMA_signal_12890 ;
    wire new_AGEMA_signal_12891 ;
    wire new_AGEMA_signal_12892 ;
    wire new_AGEMA_signal_12893 ;
    wire new_AGEMA_signal_12894 ;
    wire new_AGEMA_signal_12895 ;
    wire new_AGEMA_signal_12896 ;
    wire new_AGEMA_signal_12897 ;
    wire new_AGEMA_signal_12898 ;
    wire new_AGEMA_signal_12899 ;
    wire new_AGEMA_signal_12900 ;
    wire new_AGEMA_signal_12901 ;
    wire new_AGEMA_signal_12902 ;
    wire new_AGEMA_signal_12903 ;
    wire new_AGEMA_signal_12904 ;
    wire new_AGEMA_signal_12905 ;
    wire new_AGEMA_signal_12906 ;
    wire new_AGEMA_signal_12907 ;
    wire new_AGEMA_signal_12908 ;
    wire new_AGEMA_signal_12909 ;
    wire new_AGEMA_signal_12910 ;
    wire new_AGEMA_signal_12911 ;
    wire new_AGEMA_signal_12912 ;
    wire new_AGEMA_signal_12913 ;
    wire new_AGEMA_signal_12914 ;
    wire new_AGEMA_signal_12915 ;
    wire new_AGEMA_signal_12916 ;
    wire new_AGEMA_signal_12917 ;
    wire new_AGEMA_signal_12918 ;
    wire new_AGEMA_signal_12919 ;
    wire new_AGEMA_signal_12920 ;
    wire new_AGEMA_signal_12921 ;
    wire new_AGEMA_signal_12922 ;
    wire new_AGEMA_signal_12923 ;
    wire new_AGEMA_signal_12924 ;
    wire new_AGEMA_signal_12925 ;
    wire new_AGEMA_signal_12926 ;
    wire new_AGEMA_signal_12927 ;
    wire new_AGEMA_signal_12928 ;
    wire new_AGEMA_signal_12929 ;
    wire new_AGEMA_signal_12930 ;
    wire new_AGEMA_signal_12931 ;
    wire new_AGEMA_signal_12932 ;
    wire new_AGEMA_signal_12933 ;
    wire new_AGEMA_signal_12934 ;
    wire new_AGEMA_signal_12935 ;
    wire new_AGEMA_signal_12936 ;
    wire new_AGEMA_signal_12937 ;
    wire new_AGEMA_signal_12938 ;
    wire new_AGEMA_signal_12939 ;
    wire new_AGEMA_signal_12940 ;
    wire new_AGEMA_signal_12941 ;
    wire new_AGEMA_signal_12942 ;
    wire new_AGEMA_signal_12943 ;
    wire new_AGEMA_signal_12944 ;
    wire new_AGEMA_signal_12945 ;
    wire new_AGEMA_signal_12946 ;
    wire new_AGEMA_signal_12947 ;
    wire new_AGEMA_signal_12948 ;
    wire new_AGEMA_signal_12949 ;
    wire new_AGEMA_signal_12950 ;
    wire new_AGEMA_signal_12951 ;
    wire new_AGEMA_signal_12952 ;
    wire new_AGEMA_signal_12953 ;
    wire new_AGEMA_signal_12954 ;
    wire new_AGEMA_signal_12955 ;
    wire new_AGEMA_signal_12956 ;
    wire new_AGEMA_signal_12957 ;
    wire new_AGEMA_signal_12958 ;
    wire new_AGEMA_signal_12959 ;
    wire new_AGEMA_signal_12960 ;
    wire new_AGEMA_signal_12961 ;
    wire new_AGEMA_signal_12962 ;
    wire new_AGEMA_signal_12963 ;
    wire new_AGEMA_signal_12964 ;
    wire new_AGEMA_signal_12965 ;
    wire new_AGEMA_signal_12966 ;
    wire new_AGEMA_signal_12967 ;
    wire new_AGEMA_signal_12968 ;
    wire new_AGEMA_signal_12969 ;
    wire new_AGEMA_signal_12970 ;
    wire new_AGEMA_signal_12971 ;
    wire new_AGEMA_signal_12972 ;
    wire new_AGEMA_signal_12973 ;
    wire new_AGEMA_signal_12974 ;
    wire new_AGEMA_signal_12975 ;
    wire new_AGEMA_signal_12976 ;
    wire new_AGEMA_signal_12977 ;
    wire new_AGEMA_signal_12978 ;
    wire new_AGEMA_signal_12979 ;
    wire new_AGEMA_signal_12980 ;
    wire new_AGEMA_signal_12981 ;
    wire new_AGEMA_signal_12982 ;
    wire new_AGEMA_signal_12983 ;
    wire new_AGEMA_signal_12984 ;
    wire new_AGEMA_signal_12985 ;
    wire new_AGEMA_signal_12986 ;
    wire new_AGEMA_signal_12987 ;
    wire new_AGEMA_signal_12988 ;
    wire new_AGEMA_signal_12989 ;
    wire new_AGEMA_signal_12990 ;
    wire new_AGEMA_signal_12991 ;
    wire new_AGEMA_signal_12992 ;
    wire new_AGEMA_signal_12993 ;
    wire new_AGEMA_signal_12994 ;
    wire new_AGEMA_signal_12995 ;
    wire new_AGEMA_signal_12996 ;
    wire new_AGEMA_signal_12997 ;
    wire new_AGEMA_signal_12998 ;
    wire new_AGEMA_signal_12999 ;
    wire new_AGEMA_signal_13000 ;
    wire new_AGEMA_signal_13001 ;
    wire new_AGEMA_signal_13002 ;
    wire new_AGEMA_signal_13003 ;
    wire new_AGEMA_signal_13004 ;
    wire new_AGEMA_signal_13005 ;
    wire new_AGEMA_signal_13006 ;
    wire new_AGEMA_signal_13007 ;
    wire new_AGEMA_signal_13008 ;
    wire new_AGEMA_signal_13009 ;
    wire new_AGEMA_signal_13010 ;
    wire new_AGEMA_signal_13011 ;
    wire new_AGEMA_signal_13012 ;
    wire new_AGEMA_signal_13013 ;
    wire new_AGEMA_signal_13014 ;
    wire new_AGEMA_signal_13015 ;
    wire new_AGEMA_signal_13016 ;
    wire new_AGEMA_signal_13017 ;
    wire new_AGEMA_signal_13018 ;
    wire new_AGEMA_signal_13019 ;
    wire new_AGEMA_signal_13020 ;
    wire new_AGEMA_signal_13021 ;
    wire new_AGEMA_signal_13022 ;
    wire new_AGEMA_signal_13023 ;
    wire new_AGEMA_signal_13024 ;
    wire new_AGEMA_signal_13025 ;
    wire new_AGEMA_signal_13026 ;
    wire new_AGEMA_signal_13027 ;
    wire new_AGEMA_signal_13028 ;
    wire new_AGEMA_signal_13029 ;
    wire new_AGEMA_signal_13030 ;
    wire new_AGEMA_signal_13031 ;
    wire new_AGEMA_signal_13032 ;
    wire new_AGEMA_signal_13033 ;
    wire new_AGEMA_signal_13034 ;
    wire new_AGEMA_signal_13035 ;
    wire new_AGEMA_signal_13036 ;
    wire new_AGEMA_signal_13037 ;
    wire new_AGEMA_signal_13038 ;
    wire new_AGEMA_signal_13039 ;
    wire new_AGEMA_signal_13040 ;
    wire new_AGEMA_signal_13041 ;
    wire new_AGEMA_signal_13042 ;
    wire new_AGEMA_signal_13043 ;
    wire new_AGEMA_signal_13044 ;
    wire new_AGEMA_signal_13045 ;
    wire new_AGEMA_signal_13046 ;
    wire new_AGEMA_signal_13047 ;
    wire new_AGEMA_signal_13048 ;
    wire new_AGEMA_signal_13049 ;
    wire new_AGEMA_signal_13050 ;
    wire new_AGEMA_signal_13051 ;
    wire new_AGEMA_signal_13052 ;
    wire new_AGEMA_signal_13053 ;
    wire new_AGEMA_signal_13054 ;
    wire new_AGEMA_signal_13055 ;
    wire new_AGEMA_signal_13056 ;
    wire new_AGEMA_signal_13057 ;
    wire new_AGEMA_signal_13058 ;
    wire new_AGEMA_signal_13059 ;
    wire new_AGEMA_signal_13060 ;
    wire new_AGEMA_signal_13061 ;
    wire new_AGEMA_signal_13062 ;
    wire new_AGEMA_signal_13063 ;
    wire new_AGEMA_signal_13064 ;
    wire new_AGEMA_signal_13065 ;
    wire new_AGEMA_signal_13066 ;
    wire new_AGEMA_signal_13067 ;
    wire new_AGEMA_signal_13068 ;
    wire new_AGEMA_signal_13069 ;
    wire new_AGEMA_signal_13070 ;
    wire new_AGEMA_signal_13071 ;
    wire new_AGEMA_signal_13072 ;
    wire new_AGEMA_signal_13073 ;
    wire new_AGEMA_signal_13074 ;
    wire new_AGEMA_signal_13075 ;
    wire new_AGEMA_signal_13076 ;
    wire new_AGEMA_signal_13077 ;
    wire new_AGEMA_signal_13078 ;
    wire new_AGEMA_signal_13079 ;
    wire new_AGEMA_signal_13080 ;
    wire new_AGEMA_signal_13081 ;
    wire new_AGEMA_signal_13082 ;
    wire new_AGEMA_signal_13083 ;
    wire new_AGEMA_signal_13084 ;
    wire new_AGEMA_signal_13085 ;
    wire new_AGEMA_signal_13086 ;
    wire new_AGEMA_signal_13087 ;
    wire new_AGEMA_signal_13088 ;
    wire new_AGEMA_signal_13089 ;
    wire new_AGEMA_signal_13090 ;
    wire new_AGEMA_signal_13091 ;
    wire new_AGEMA_signal_13092 ;
    wire new_AGEMA_signal_13093 ;
    wire new_AGEMA_signal_13094 ;
    wire new_AGEMA_signal_13095 ;
    wire new_AGEMA_signal_13096 ;
    wire new_AGEMA_signal_13097 ;
    wire new_AGEMA_signal_13098 ;
    wire new_AGEMA_signal_13099 ;
    wire new_AGEMA_signal_13100 ;
    wire new_AGEMA_signal_13101 ;
    wire new_AGEMA_signal_13102 ;
    wire new_AGEMA_signal_13103 ;
    wire new_AGEMA_signal_13104 ;
    wire new_AGEMA_signal_13105 ;
    wire new_AGEMA_signal_13106 ;
    wire new_AGEMA_signal_13107 ;
    wire new_AGEMA_signal_13108 ;
    wire new_AGEMA_signal_13109 ;
    wire new_AGEMA_signal_13110 ;
    wire new_AGEMA_signal_13111 ;
    wire new_AGEMA_signal_13112 ;
    wire new_AGEMA_signal_13113 ;
    wire new_AGEMA_signal_13114 ;
    wire new_AGEMA_signal_13115 ;
    wire new_AGEMA_signal_13116 ;
    wire new_AGEMA_signal_13117 ;
    wire new_AGEMA_signal_13118 ;
    wire new_AGEMA_signal_13119 ;
    wire new_AGEMA_signal_13120 ;
    wire new_AGEMA_signal_13121 ;
    wire new_AGEMA_signal_13122 ;
    wire new_AGEMA_signal_13123 ;
    wire new_AGEMA_signal_13124 ;
    wire new_AGEMA_signal_13125 ;
    wire new_AGEMA_signal_13126 ;
    wire new_AGEMA_signal_13127 ;
    wire new_AGEMA_signal_13128 ;
    wire new_AGEMA_signal_13129 ;
    wire new_AGEMA_signal_13130 ;
    wire new_AGEMA_signal_13131 ;
    wire new_AGEMA_signal_13132 ;
    wire new_AGEMA_signal_13133 ;
    wire new_AGEMA_signal_13134 ;
    wire new_AGEMA_signal_13135 ;
    wire new_AGEMA_signal_13136 ;
    wire new_AGEMA_signal_13137 ;
    wire new_AGEMA_signal_13138 ;
    wire new_AGEMA_signal_13139 ;
    wire new_AGEMA_signal_13140 ;
    wire new_AGEMA_signal_13141 ;
    wire new_AGEMA_signal_13142 ;
    wire new_AGEMA_signal_13143 ;
    wire new_AGEMA_signal_13144 ;
    wire new_AGEMA_signal_13145 ;
    wire new_AGEMA_signal_13146 ;
    wire new_AGEMA_signal_13147 ;
    wire new_AGEMA_signal_13148 ;
    wire new_AGEMA_signal_13149 ;
    wire new_AGEMA_signal_13150 ;
    wire new_AGEMA_signal_13151 ;
    wire new_AGEMA_signal_13152 ;
    wire new_AGEMA_signal_13153 ;
    wire new_AGEMA_signal_13154 ;
    wire new_AGEMA_signal_13155 ;
    wire new_AGEMA_signal_13156 ;
    wire new_AGEMA_signal_13157 ;
    wire new_AGEMA_signal_13158 ;
    wire new_AGEMA_signal_13159 ;
    wire new_AGEMA_signal_13160 ;
    wire new_AGEMA_signal_13161 ;
    wire new_AGEMA_signal_13162 ;
    wire new_AGEMA_signal_13163 ;
    wire new_AGEMA_signal_13164 ;
    wire new_AGEMA_signal_13165 ;
    wire new_AGEMA_signal_13166 ;
    wire new_AGEMA_signal_13167 ;
    wire new_AGEMA_signal_13168 ;
    wire new_AGEMA_signal_13169 ;
    wire new_AGEMA_signal_13170 ;
    wire new_AGEMA_signal_13171 ;
    wire new_AGEMA_signal_13172 ;
    wire new_AGEMA_signal_13173 ;
    wire new_AGEMA_signal_13174 ;
    wire new_AGEMA_signal_13175 ;
    wire new_AGEMA_signal_13176 ;
    wire new_AGEMA_signal_13177 ;
    wire new_AGEMA_signal_13178 ;
    wire new_AGEMA_signal_13179 ;
    wire new_AGEMA_signal_13180 ;
    wire new_AGEMA_signal_13181 ;
    wire new_AGEMA_signal_13182 ;
    wire new_AGEMA_signal_13183 ;
    wire new_AGEMA_signal_13184 ;
    wire new_AGEMA_signal_13185 ;
    wire new_AGEMA_signal_13186 ;
    wire new_AGEMA_signal_13187 ;
    wire new_AGEMA_signal_13188 ;
    wire new_AGEMA_signal_13189 ;
    wire new_AGEMA_signal_13190 ;
    wire new_AGEMA_signal_13191 ;
    wire new_AGEMA_signal_13192 ;
    wire new_AGEMA_signal_13193 ;
    wire new_AGEMA_signal_13194 ;
    wire new_AGEMA_signal_13195 ;
    wire new_AGEMA_signal_13196 ;
    wire new_AGEMA_signal_13197 ;
    wire new_AGEMA_signal_13198 ;
    wire new_AGEMA_signal_13199 ;
    wire new_AGEMA_signal_13200 ;
    wire new_AGEMA_signal_13201 ;
    wire new_AGEMA_signal_13202 ;
    wire new_AGEMA_signal_13203 ;
    wire new_AGEMA_signal_13204 ;
    wire new_AGEMA_signal_13205 ;
    wire new_AGEMA_signal_13206 ;
    wire new_AGEMA_signal_13207 ;
    wire new_AGEMA_signal_13208 ;
    wire new_AGEMA_signal_13209 ;
    wire new_AGEMA_signal_13210 ;
    wire new_AGEMA_signal_13211 ;
    wire new_AGEMA_signal_13212 ;
    wire new_AGEMA_signal_13213 ;
    wire new_AGEMA_signal_13214 ;
    wire new_AGEMA_signal_13215 ;
    wire new_AGEMA_signal_13216 ;
    wire new_AGEMA_signal_13217 ;
    wire new_AGEMA_signal_13218 ;
    wire new_AGEMA_signal_13219 ;
    wire new_AGEMA_signal_13220 ;
    wire new_AGEMA_signal_13221 ;
    wire new_AGEMA_signal_13222 ;
    wire new_AGEMA_signal_13223 ;
    wire new_AGEMA_signal_13224 ;
    wire new_AGEMA_signal_13225 ;
    wire new_AGEMA_signal_13226 ;
    wire new_AGEMA_signal_13227 ;
    wire new_AGEMA_signal_13228 ;
    wire new_AGEMA_signal_13229 ;
    wire new_AGEMA_signal_13230 ;
    wire new_AGEMA_signal_13231 ;
    wire new_AGEMA_signal_13232 ;
    wire new_AGEMA_signal_13233 ;
    wire new_AGEMA_signal_13234 ;
    wire new_AGEMA_signal_13235 ;
    wire new_AGEMA_signal_13236 ;
    wire new_AGEMA_signal_13237 ;
    wire new_AGEMA_signal_13238 ;
    wire new_AGEMA_signal_13239 ;
    wire new_AGEMA_signal_13240 ;
    wire new_AGEMA_signal_13241 ;
    wire new_AGEMA_signal_13242 ;
    wire new_AGEMA_signal_13243 ;
    wire new_AGEMA_signal_13244 ;
    wire new_AGEMA_signal_13245 ;
    wire new_AGEMA_signal_13246 ;
    wire new_AGEMA_signal_13247 ;
    wire new_AGEMA_signal_13248 ;
    wire new_AGEMA_signal_13249 ;
    wire new_AGEMA_signal_13250 ;
    wire new_AGEMA_signal_13251 ;
    wire new_AGEMA_signal_13252 ;
    wire new_AGEMA_signal_13253 ;
    wire new_AGEMA_signal_13254 ;
    wire new_AGEMA_signal_13255 ;
    wire new_AGEMA_signal_13256 ;
    wire new_AGEMA_signal_13257 ;
    wire new_AGEMA_signal_13258 ;
    wire new_AGEMA_signal_13259 ;
    wire new_AGEMA_signal_13260 ;
    wire new_AGEMA_signal_13261 ;
    wire new_AGEMA_signal_13262 ;
    wire new_AGEMA_signal_13263 ;
    wire new_AGEMA_signal_13264 ;
    wire new_AGEMA_signal_13265 ;
    wire new_AGEMA_signal_13266 ;
    wire new_AGEMA_signal_13267 ;
    wire new_AGEMA_signal_13268 ;
    wire new_AGEMA_signal_13269 ;
    wire new_AGEMA_signal_13270 ;
    wire new_AGEMA_signal_13271 ;
    wire new_AGEMA_signal_13272 ;
    wire new_AGEMA_signal_13273 ;
    wire new_AGEMA_signal_13274 ;
    wire new_AGEMA_signal_13275 ;
    wire new_AGEMA_signal_13276 ;
    wire new_AGEMA_signal_13277 ;
    wire new_AGEMA_signal_13278 ;
    wire new_AGEMA_signal_13279 ;
    wire new_AGEMA_signal_13280 ;
    wire new_AGEMA_signal_13281 ;
    wire new_AGEMA_signal_13282 ;
    wire new_AGEMA_signal_13283 ;
    wire new_AGEMA_signal_13284 ;
    wire new_AGEMA_signal_13285 ;
    wire new_AGEMA_signal_13286 ;
    wire new_AGEMA_signal_13287 ;
    wire new_AGEMA_signal_13288 ;
    wire new_AGEMA_signal_13289 ;
    wire new_AGEMA_signal_13290 ;
    wire new_AGEMA_signal_13291 ;
    wire new_AGEMA_signal_13292 ;
    wire new_AGEMA_signal_13293 ;
    wire new_AGEMA_signal_13294 ;
    wire new_AGEMA_signal_13295 ;
    wire new_AGEMA_signal_13296 ;
    wire new_AGEMA_signal_13297 ;
    wire new_AGEMA_signal_13298 ;
    wire new_AGEMA_signal_13299 ;
    wire new_AGEMA_signal_13300 ;
    wire new_AGEMA_signal_13301 ;
    wire new_AGEMA_signal_13302 ;
    wire new_AGEMA_signal_13303 ;
    wire new_AGEMA_signal_13304 ;
    wire new_AGEMA_signal_13305 ;
    wire new_AGEMA_signal_13306 ;
    wire new_AGEMA_signal_13307 ;
    wire new_AGEMA_signal_13308 ;
    wire new_AGEMA_signal_13309 ;
    wire new_AGEMA_signal_13310 ;
    wire new_AGEMA_signal_13311 ;
    wire new_AGEMA_signal_13312 ;
    wire new_AGEMA_signal_13313 ;
    wire new_AGEMA_signal_13314 ;
    wire new_AGEMA_signal_13315 ;
    wire new_AGEMA_signal_13316 ;
    wire new_AGEMA_signal_13317 ;
    wire new_AGEMA_signal_13318 ;
    wire new_AGEMA_signal_13319 ;
    wire new_AGEMA_signal_13320 ;
    wire new_AGEMA_signal_13321 ;
    wire new_AGEMA_signal_13322 ;
    wire new_AGEMA_signal_13323 ;
    wire new_AGEMA_signal_13324 ;
    wire new_AGEMA_signal_13325 ;
    wire new_AGEMA_signal_13326 ;
    wire new_AGEMA_signal_13327 ;
    wire new_AGEMA_signal_13328 ;
    wire new_AGEMA_signal_13329 ;
    wire new_AGEMA_signal_13330 ;
    wire new_AGEMA_signal_13331 ;
    wire new_AGEMA_signal_13332 ;
    wire new_AGEMA_signal_13333 ;
    wire new_AGEMA_signal_13334 ;
    wire new_AGEMA_signal_13335 ;
    wire new_AGEMA_signal_13336 ;
    wire new_AGEMA_signal_13337 ;
    wire new_AGEMA_signal_13338 ;
    wire new_AGEMA_signal_13339 ;
    wire new_AGEMA_signal_13340 ;
    wire new_AGEMA_signal_13341 ;
    wire new_AGEMA_signal_13342 ;
    wire new_AGEMA_signal_13343 ;
    wire new_AGEMA_signal_13344 ;
    wire new_AGEMA_signal_13345 ;
    wire new_AGEMA_signal_13346 ;
    wire new_AGEMA_signal_13347 ;
    wire new_AGEMA_signal_13348 ;
    wire new_AGEMA_signal_13349 ;
    wire new_AGEMA_signal_13350 ;
    wire new_AGEMA_signal_13351 ;
    wire new_AGEMA_signal_13352 ;
    wire new_AGEMA_signal_13353 ;
    wire new_AGEMA_signal_13354 ;
    wire new_AGEMA_signal_13355 ;
    wire new_AGEMA_signal_13356 ;
    wire new_AGEMA_signal_13357 ;
    wire new_AGEMA_signal_13358 ;
    wire new_AGEMA_signal_13359 ;
    wire new_AGEMA_signal_13360 ;
    wire new_AGEMA_signal_13361 ;
    wire new_AGEMA_signal_13362 ;
    wire new_AGEMA_signal_13363 ;
    wire new_AGEMA_signal_13364 ;
    wire new_AGEMA_signal_13365 ;
    wire new_AGEMA_signal_13366 ;
    wire new_AGEMA_signal_13367 ;
    wire new_AGEMA_signal_13368 ;
    wire new_AGEMA_signal_13369 ;
    wire new_AGEMA_signal_13370 ;
    wire new_AGEMA_signal_13371 ;
    wire new_AGEMA_signal_13372 ;
    wire new_AGEMA_signal_13373 ;
    wire new_AGEMA_signal_13374 ;
    wire new_AGEMA_signal_13375 ;
    wire new_AGEMA_signal_13376 ;
    wire new_AGEMA_signal_13377 ;
    wire new_AGEMA_signal_13378 ;
    wire new_AGEMA_signal_13379 ;
    wire new_AGEMA_signal_13380 ;
    wire new_AGEMA_signal_13381 ;
    wire new_AGEMA_signal_13382 ;
    wire new_AGEMA_signal_13383 ;
    wire new_AGEMA_signal_13384 ;
    wire new_AGEMA_signal_13385 ;
    wire new_AGEMA_signal_13386 ;
    wire new_AGEMA_signal_13387 ;
    wire new_AGEMA_signal_13388 ;
    wire new_AGEMA_signal_13389 ;
    wire new_AGEMA_signal_13390 ;
    wire new_AGEMA_signal_13391 ;
    wire new_AGEMA_signal_13392 ;
    wire new_AGEMA_signal_13393 ;
    wire new_AGEMA_signal_13394 ;
    wire new_AGEMA_signal_13395 ;
    wire new_AGEMA_signal_13396 ;
    wire new_AGEMA_signal_13397 ;
    wire new_AGEMA_signal_13398 ;
    wire new_AGEMA_signal_13399 ;
    wire new_AGEMA_signal_13400 ;
    wire new_AGEMA_signal_13401 ;
    wire new_AGEMA_signal_13402 ;
    wire new_AGEMA_signal_13403 ;
    wire new_AGEMA_signal_13404 ;
    wire new_AGEMA_signal_13405 ;
    wire new_AGEMA_signal_13406 ;
    wire new_AGEMA_signal_13407 ;
    wire new_AGEMA_signal_13408 ;
    wire new_AGEMA_signal_13409 ;
    wire new_AGEMA_signal_13410 ;
    wire new_AGEMA_signal_13411 ;
    wire new_AGEMA_signal_13412 ;
    wire new_AGEMA_signal_13413 ;
    wire new_AGEMA_signal_13414 ;
    wire new_AGEMA_signal_13415 ;
    wire new_AGEMA_signal_13416 ;
    wire new_AGEMA_signal_13417 ;
    wire new_AGEMA_signal_13418 ;
    wire new_AGEMA_signal_13419 ;
    wire new_AGEMA_signal_13420 ;
    wire new_AGEMA_signal_13421 ;
    wire new_AGEMA_signal_13422 ;
    wire new_AGEMA_signal_13423 ;
    wire new_AGEMA_signal_13424 ;
    wire new_AGEMA_signal_13425 ;
    wire new_AGEMA_signal_13426 ;
    wire new_AGEMA_signal_13427 ;
    wire new_AGEMA_signal_13428 ;
    wire new_AGEMA_signal_13429 ;
    wire new_AGEMA_signal_13430 ;
    wire new_AGEMA_signal_13431 ;
    wire new_AGEMA_signal_13432 ;
    wire new_AGEMA_signal_13433 ;
    wire new_AGEMA_signal_13434 ;
    wire new_AGEMA_signal_13435 ;
    wire new_AGEMA_signal_13436 ;
    wire new_AGEMA_signal_13437 ;
    wire new_AGEMA_signal_13438 ;
    wire new_AGEMA_signal_13439 ;
    wire new_AGEMA_signal_13440 ;
    wire new_AGEMA_signal_13441 ;
    wire new_AGEMA_signal_13442 ;
    wire new_AGEMA_signal_13443 ;
    wire new_AGEMA_signal_13444 ;
    wire new_AGEMA_signal_13445 ;
    wire new_AGEMA_signal_13446 ;
    wire new_AGEMA_signal_13447 ;
    wire new_AGEMA_signal_13448 ;
    wire new_AGEMA_signal_13449 ;
    wire new_AGEMA_signal_13450 ;
    wire new_AGEMA_signal_13451 ;
    wire new_AGEMA_signal_13452 ;
    wire new_AGEMA_signal_13453 ;
    wire new_AGEMA_signal_13454 ;
    wire new_AGEMA_signal_13455 ;
    wire new_AGEMA_signal_13456 ;
    wire new_AGEMA_signal_13457 ;
    wire new_AGEMA_signal_13458 ;
    wire new_AGEMA_signal_13459 ;
    wire new_AGEMA_signal_13460 ;
    wire new_AGEMA_signal_13461 ;
    wire new_AGEMA_signal_13462 ;
    wire new_AGEMA_signal_13463 ;
    wire new_AGEMA_signal_13464 ;
    wire new_AGEMA_signal_13465 ;
    wire new_AGEMA_signal_13466 ;
    wire new_AGEMA_signal_13467 ;
    wire new_AGEMA_signal_13468 ;
    wire new_AGEMA_signal_13469 ;
    wire new_AGEMA_signal_13470 ;
    wire new_AGEMA_signal_13471 ;
    wire new_AGEMA_signal_13472 ;
    wire new_AGEMA_signal_13473 ;
    wire new_AGEMA_signal_13474 ;
    wire new_AGEMA_signal_13475 ;
    wire new_AGEMA_signal_13476 ;
    wire new_AGEMA_signal_13477 ;
    wire new_AGEMA_signal_13478 ;
    wire new_AGEMA_signal_13479 ;
    wire new_AGEMA_signal_13480 ;
    wire new_AGEMA_signal_13481 ;
    wire new_AGEMA_signal_13482 ;
    wire new_AGEMA_signal_13483 ;
    wire new_AGEMA_signal_13484 ;
    wire new_AGEMA_signal_13485 ;
    wire new_AGEMA_signal_13486 ;
    wire new_AGEMA_signal_13487 ;
    wire new_AGEMA_signal_13488 ;
    wire new_AGEMA_signal_13489 ;
    wire new_AGEMA_signal_13490 ;
    wire new_AGEMA_signal_13491 ;
    wire new_AGEMA_signal_13492 ;
    wire new_AGEMA_signal_13493 ;
    wire new_AGEMA_signal_13494 ;
    wire new_AGEMA_signal_13495 ;
    wire new_AGEMA_signal_13496 ;
    wire new_AGEMA_signal_13497 ;
    wire new_AGEMA_signal_13498 ;
    wire new_AGEMA_signal_13499 ;
    wire new_AGEMA_signal_13500 ;
    wire new_AGEMA_signal_13501 ;
    wire new_AGEMA_signal_13502 ;
    wire new_AGEMA_signal_13503 ;
    wire new_AGEMA_signal_13504 ;
    wire new_AGEMA_signal_13505 ;
    wire new_AGEMA_signal_13506 ;
    wire new_AGEMA_signal_13507 ;
    wire new_AGEMA_signal_13508 ;
    wire new_AGEMA_signal_13509 ;
    wire new_AGEMA_signal_13510 ;
    wire new_AGEMA_signal_13511 ;
    wire new_AGEMA_signal_13512 ;
    wire new_AGEMA_signal_13513 ;
    wire new_AGEMA_signal_13514 ;
    wire new_AGEMA_signal_13515 ;
    wire new_AGEMA_signal_13516 ;
    wire new_AGEMA_signal_13517 ;
    wire new_AGEMA_signal_13518 ;
    wire new_AGEMA_signal_13519 ;
    wire new_AGEMA_signal_13520 ;
    wire new_AGEMA_signal_13521 ;
    wire new_AGEMA_signal_13522 ;
    wire new_AGEMA_signal_13523 ;
    wire new_AGEMA_signal_13524 ;
    wire new_AGEMA_signal_13525 ;
    wire new_AGEMA_signal_13526 ;
    wire new_AGEMA_signal_13527 ;
    wire new_AGEMA_signal_13528 ;
    wire new_AGEMA_signal_13529 ;
    wire new_AGEMA_signal_13530 ;
    wire new_AGEMA_signal_13531 ;
    wire new_AGEMA_signal_13532 ;
    wire new_AGEMA_signal_13533 ;
    wire new_AGEMA_signal_13534 ;
    wire new_AGEMA_signal_13535 ;
    wire new_AGEMA_signal_13536 ;
    wire new_AGEMA_signal_13537 ;
    wire new_AGEMA_signal_13538 ;
    wire new_AGEMA_signal_13539 ;
    wire new_AGEMA_signal_13540 ;
    wire new_AGEMA_signal_13541 ;
    wire new_AGEMA_signal_13542 ;
    wire new_AGEMA_signal_13543 ;
    wire new_AGEMA_signal_13544 ;
    wire new_AGEMA_signal_13545 ;
    wire new_AGEMA_signal_13546 ;
    wire new_AGEMA_signal_13547 ;
    wire new_AGEMA_signal_13548 ;
    wire new_AGEMA_signal_13549 ;
    wire new_AGEMA_signal_13550 ;
    wire new_AGEMA_signal_13551 ;
    wire new_AGEMA_signal_13552 ;
    wire new_AGEMA_signal_13553 ;
    wire new_AGEMA_signal_13554 ;
    wire new_AGEMA_signal_13555 ;
    wire new_AGEMA_signal_13556 ;
    wire new_AGEMA_signal_13557 ;
    wire new_AGEMA_signal_13558 ;
    wire new_AGEMA_signal_13559 ;
    wire new_AGEMA_signal_13560 ;
    wire new_AGEMA_signal_13561 ;
    wire new_AGEMA_signal_13562 ;
    wire new_AGEMA_signal_13563 ;
    wire new_AGEMA_signal_13564 ;
    wire new_AGEMA_signal_13565 ;
    wire new_AGEMA_signal_13566 ;
    wire new_AGEMA_signal_13567 ;
    wire new_AGEMA_signal_13568 ;
    wire new_AGEMA_signal_13569 ;
    wire new_AGEMA_signal_13570 ;
    wire new_AGEMA_signal_13571 ;
    wire new_AGEMA_signal_13572 ;
    wire new_AGEMA_signal_13573 ;
    wire new_AGEMA_signal_13574 ;
    wire new_AGEMA_signal_13575 ;
    wire new_AGEMA_signal_13576 ;
    wire new_AGEMA_signal_13577 ;
    wire new_AGEMA_signal_13578 ;
    wire new_AGEMA_signal_13579 ;
    wire new_AGEMA_signal_13580 ;
    wire new_AGEMA_signal_13581 ;
    wire new_AGEMA_signal_13582 ;
    wire new_AGEMA_signal_13583 ;
    wire new_AGEMA_signal_13584 ;
    wire new_AGEMA_signal_13585 ;
    wire new_AGEMA_signal_13586 ;
    wire new_AGEMA_signal_13587 ;
    wire new_AGEMA_signal_13588 ;
    wire new_AGEMA_signal_13589 ;
    wire new_AGEMA_signal_13590 ;
    wire new_AGEMA_signal_13591 ;
    wire new_AGEMA_signal_13592 ;
    wire new_AGEMA_signal_13593 ;
    wire new_AGEMA_signal_13594 ;
    wire new_AGEMA_signal_13595 ;
    wire new_AGEMA_signal_13596 ;
    wire new_AGEMA_signal_13597 ;
    wire new_AGEMA_signal_13598 ;
    wire new_AGEMA_signal_13599 ;
    wire new_AGEMA_signal_13600 ;
    wire new_AGEMA_signal_13601 ;
    wire new_AGEMA_signal_13602 ;
    wire new_AGEMA_signal_13603 ;
    wire new_AGEMA_signal_13604 ;
    wire new_AGEMA_signal_13605 ;
    wire new_AGEMA_signal_13606 ;
    wire new_AGEMA_signal_13607 ;
    wire new_AGEMA_signal_13608 ;
    wire new_AGEMA_signal_13609 ;
    wire new_AGEMA_signal_13610 ;
    wire new_AGEMA_signal_13611 ;
    wire new_AGEMA_signal_13612 ;
    wire new_AGEMA_signal_13613 ;
    wire new_AGEMA_signal_13614 ;
    wire new_AGEMA_signal_13615 ;
    wire new_AGEMA_signal_13616 ;
    wire new_AGEMA_signal_13617 ;
    wire new_AGEMA_signal_13618 ;
    wire new_AGEMA_signal_13619 ;
    wire new_AGEMA_signal_13620 ;
    wire new_AGEMA_signal_13621 ;
    wire new_AGEMA_signal_13622 ;
    wire new_AGEMA_signal_13623 ;
    wire new_AGEMA_signal_13624 ;
    wire new_AGEMA_signal_13625 ;
    wire new_AGEMA_signal_13626 ;
    wire new_AGEMA_signal_13627 ;
    wire new_AGEMA_signal_13628 ;
    wire new_AGEMA_signal_13629 ;
    wire new_AGEMA_signal_13630 ;
    wire new_AGEMA_signal_13631 ;
    wire new_AGEMA_signal_13632 ;
    wire new_AGEMA_signal_13633 ;
    wire new_AGEMA_signal_13634 ;
    wire new_AGEMA_signal_13635 ;
    wire new_AGEMA_signal_13636 ;
    wire new_AGEMA_signal_13637 ;
    wire new_AGEMA_signal_13638 ;
    wire new_AGEMA_signal_13639 ;
    wire new_AGEMA_signal_13640 ;
    wire new_AGEMA_signal_13641 ;
    wire new_AGEMA_signal_13642 ;
    wire new_AGEMA_signal_13643 ;
    wire new_AGEMA_signal_13644 ;
    wire new_AGEMA_signal_13645 ;
    wire new_AGEMA_signal_13646 ;
    wire new_AGEMA_signal_13647 ;
    wire new_AGEMA_signal_13648 ;
    wire new_AGEMA_signal_13649 ;
    wire new_AGEMA_signal_13650 ;
    wire new_AGEMA_signal_13651 ;
    wire new_AGEMA_signal_13652 ;
    wire new_AGEMA_signal_13653 ;
    wire new_AGEMA_signal_13654 ;
    wire new_AGEMA_signal_13655 ;
    wire new_AGEMA_signal_13656 ;
    wire new_AGEMA_signal_13657 ;
    wire new_AGEMA_signal_13658 ;
    wire new_AGEMA_signal_13659 ;
    wire new_AGEMA_signal_13660 ;
    wire new_AGEMA_signal_13661 ;
    wire new_AGEMA_signal_13662 ;
    wire new_AGEMA_signal_13663 ;
    wire new_AGEMA_signal_13664 ;
    wire new_AGEMA_signal_13665 ;
    wire new_AGEMA_signal_13666 ;
    wire new_AGEMA_signal_13667 ;
    wire new_AGEMA_signal_13668 ;
    wire new_AGEMA_signal_13669 ;
    wire new_AGEMA_signal_13670 ;
    wire new_AGEMA_signal_13671 ;
    wire new_AGEMA_signal_13672 ;
    wire new_AGEMA_signal_13673 ;
    wire new_AGEMA_signal_13674 ;
    wire new_AGEMA_signal_13675 ;
    wire new_AGEMA_signal_13676 ;
    wire new_AGEMA_signal_13677 ;
    wire new_AGEMA_signal_13678 ;
    wire new_AGEMA_signal_13679 ;
    wire new_AGEMA_signal_13680 ;
    wire new_AGEMA_signal_13681 ;
    wire new_AGEMA_signal_13682 ;
    wire new_AGEMA_signal_13683 ;
    wire new_AGEMA_signal_13684 ;
    wire new_AGEMA_signal_13685 ;
    wire new_AGEMA_signal_13686 ;
    wire new_AGEMA_signal_13687 ;
    wire new_AGEMA_signal_13688 ;
    wire new_AGEMA_signal_13689 ;
    wire new_AGEMA_signal_13690 ;
    wire new_AGEMA_signal_13691 ;
    wire new_AGEMA_signal_13692 ;
    wire new_AGEMA_signal_13693 ;
    wire new_AGEMA_signal_13694 ;
    wire new_AGEMA_signal_13695 ;
    wire new_AGEMA_signal_13696 ;
    wire new_AGEMA_signal_13697 ;
    wire new_AGEMA_signal_13698 ;
    wire new_AGEMA_signal_13699 ;
    wire new_AGEMA_signal_13700 ;
    wire new_AGEMA_signal_13701 ;
    wire new_AGEMA_signal_13702 ;
    wire new_AGEMA_signal_13703 ;
    wire new_AGEMA_signal_13704 ;
    wire new_AGEMA_signal_13705 ;
    wire new_AGEMA_signal_13706 ;
    wire new_AGEMA_signal_13707 ;
    wire new_AGEMA_signal_13708 ;
    wire new_AGEMA_signal_13709 ;
    wire new_AGEMA_signal_13710 ;
    wire new_AGEMA_signal_13711 ;
    wire new_AGEMA_signal_13712 ;
    wire new_AGEMA_signal_13713 ;
    wire new_AGEMA_signal_13714 ;
    wire new_AGEMA_signal_13715 ;
    wire new_AGEMA_signal_13716 ;
    wire new_AGEMA_signal_13717 ;
    wire new_AGEMA_signal_13718 ;
    wire new_AGEMA_signal_13719 ;
    wire new_AGEMA_signal_13720 ;
    wire new_AGEMA_signal_13721 ;
    wire new_AGEMA_signal_13722 ;
    wire new_AGEMA_signal_13723 ;
    wire new_AGEMA_signal_13724 ;
    wire new_AGEMA_signal_13725 ;
    wire new_AGEMA_signal_13726 ;
    wire new_AGEMA_signal_13727 ;
    wire new_AGEMA_signal_13728 ;
    wire new_AGEMA_signal_13729 ;
    wire new_AGEMA_signal_13730 ;
    wire new_AGEMA_signal_13731 ;
    wire new_AGEMA_signal_13732 ;
    wire new_AGEMA_signal_13733 ;
    wire new_AGEMA_signal_13734 ;
    wire new_AGEMA_signal_13735 ;
    wire new_AGEMA_signal_13736 ;
    wire new_AGEMA_signal_13737 ;
    wire new_AGEMA_signal_13738 ;
    wire new_AGEMA_signal_13739 ;
    wire new_AGEMA_signal_13740 ;
    wire new_AGEMA_signal_13741 ;
    wire new_AGEMA_signal_13742 ;
    wire new_AGEMA_signal_13743 ;
    wire new_AGEMA_signal_13744 ;
    wire new_AGEMA_signal_13745 ;
    wire new_AGEMA_signal_13746 ;
    wire new_AGEMA_signal_13747 ;
    wire new_AGEMA_signal_13748 ;
    wire new_AGEMA_signal_13749 ;
    wire new_AGEMA_signal_13750 ;
    wire new_AGEMA_signal_13751 ;
    wire new_AGEMA_signal_13752 ;
    wire new_AGEMA_signal_13753 ;
    wire new_AGEMA_signal_13754 ;
    wire new_AGEMA_signal_13755 ;
    wire new_AGEMA_signal_13756 ;
    wire new_AGEMA_signal_13757 ;
    wire new_AGEMA_signal_13758 ;
    wire new_AGEMA_signal_13759 ;
    wire new_AGEMA_signal_13760 ;
    wire new_AGEMA_signal_13761 ;
    wire new_AGEMA_signal_13762 ;
    wire new_AGEMA_signal_13763 ;
    wire new_AGEMA_signal_13764 ;
    wire new_AGEMA_signal_13765 ;
    wire new_AGEMA_signal_13766 ;
    wire new_AGEMA_signal_13767 ;
    wire new_AGEMA_signal_13768 ;
    wire new_AGEMA_signal_13769 ;
    wire new_AGEMA_signal_13770 ;
    wire new_AGEMA_signal_13771 ;
    wire new_AGEMA_signal_13772 ;
    wire new_AGEMA_signal_13773 ;
    wire new_AGEMA_signal_13774 ;
    wire new_AGEMA_signal_13775 ;
    wire new_AGEMA_signal_13776 ;
    wire new_AGEMA_signal_13777 ;
    wire new_AGEMA_signal_13778 ;
    wire new_AGEMA_signal_13779 ;
    wire new_AGEMA_signal_13780 ;
    wire new_AGEMA_signal_13781 ;
    wire new_AGEMA_signal_13782 ;
    wire new_AGEMA_signal_13783 ;
    wire new_AGEMA_signal_13784 ;
    wire new_AGEMA_signal_13785 ;
    wire new_AGEMA_signal_13786 ;
    wire new_AGEMA_signal_13787 ;
    wire new_AGEMA_signal_13788 ;
    wire new_AGEMA_signal_13789 ;
    wire new_AGEMA_signal_13790 ;
    wire new_AGEMA_signal_13791 ;
    wire new_AGEMA_signal_13792 ;
    wire new_AGEMA_signal_13793 ;
    wire new_AGEMA_signal_13794 ;
    wire new_AGEMA_signal_13795 ;
    wire new_AGEMA_signal_13796 ;
    wire new_AGEMA_signal_13797 ;
    wire new_AGEMA_signal_13798 ;
    wire new_AGEMA_signal_13799 ;
    wire new_AGEMA_signal_13800 ;
    wire new_AGEMA_signal_13801 ;
    wire new_AGEMA_signal_13802 ;
    wire new_AGEMA_signal_13803 ;
    wire new_AGEMA_signal_13804 ;
    wire new_AGEMA_signal_13805 ;
    wire new_AGEMA_signal_13806 ;
    wire new_AGEMA_signal_13807 ;
    wire new_AGEMA_signal_13808 ;
    wire new_AGEMA_signal_13809 ;
    wire new_AGEMA_signal_13810 ;
    wire new_AGEMA_signal_13811 ;
    wire new_AGEMA_signal_13812 ;
    wire new_AGEMA_signal_13813 ;
    wire new_AGEMA_signal_13814 ;
    wire new_AGEMA_signal_13815 ;
    wire new_AGEMA_signal_13816 ;
    wire new_AGEMA_signal_13817 ;
    wire new_AGEMA_signal_13818 ;
    wire new_AGEMA_signal_13819 ;
    wire new_AGEMA_signal_13820 ;
    wire new_AGEMA_signal_13821 ;
    wire new_AGEMA_signal_13822 ;
    wire new_AGEMA_signal_13823 ;
    wire new_AGEMA_signal_13824 ;
    wire new_AGEMA_signal_13825 ;
    wire new_AGEMA_signal_13826 ;
    wire new_AGEMA_signal_13827 ;
    wire new_AGEMA_signal_13828 ;
    wire new_AGEMA_signal_13829 ;
    wire new_AGEMA_signal_13830 ;
    wire new_AGEMA_signal_13831 ;
    wire new_AGEMA_signal_13832 ;
    wire new_AGEMA_signal_13833 ;
    wire new_AGEMA_signal_13834 ;
    wire new_AGEMA_signal_13835 ;
    wire new_AGEMA_signal_13836 ;
    wire new_AGEMA_signal_13837 ;
    wire new_AGEMA_signal_13838 ;
    wire new_AGEMA_signal_13839 ;
    wire new_AGEMA_signal_13840 ;
    wire new_AGEMA_signal_13841 ;
    wire new_AGEMA_signal_13842 ;
    wire new_AGEMA_signal_13843 ;
    wire new_AGEMA_signal_13844 ;
    wire new_AGEMA_signal_13845 ;
    wire new_AGEMA_signal_13846 ;
    wire new_AGEMA_signal_13847 ;
    wire new_AGEMA_signal_13848 ;
    wire new_AGEMA_signal_13849 ;
    wire new_AGEMA_signal_13850 ;
    wire new_AGEMA_signal_13851 ;
    wire new_AGEMA_signal_13852 ;
    wire new_AGEMA_signal_13853 ;
    wire new_AGEMA_signal_13854 ;
    wire new_AGEMA_signal_13855 ;
    wire new_AGEMA_signal_13856 ;
    wire new_AGEMA_signal_13857 ;
    wire new_AGEMA_signal_13858 ;
    wire new_AGEMA_signal_13859 ;
    wire new_AGEMA_signal_13860 ;
    wire new_AGEMA_signal_13861 ;
    wire new_AGEMA_signal_13862 ;
    wire new_AGEMA_signal_13863 ;
    wire new_AGEMA_signal_13864 ;
    wire new_AGEMA_signal_13865 ;
    wire new_AGEMA_signal_13866 ;
    wire new_AGEMA_signal_13867 ;
    wire new_AGEMA_signal_13868 ;
    wire new_AGEMA_signal_13869 ;
    wire new_AGEMA_signal_13870 ;
    wire new_AGEMA_signal_13871 ;
    wire new_AGEMA_signal_13872 ;
    wire new_AGEMA_signal_13873 ;
    wire new_AGEMA_signal_13874 ;
    wire new_AGEMA_signal_13875 ;
    wire new_AGEMA_signal_13876 ;
    wire new_AGEMA_signal_13877 ;
    wire new_AGEMA_signal_13878 ;
    wire new_AGEMA_signal_13879 ;
    wire new_AGEMA_signal_13880 ;
    wire new_AGEMA_signal_13881 ;
    wire new_AGEMA_signal_13882 ;
    wire new_AGEMA_signal_13883 ;
    wire new_AGEMA_signal_13884 ;
    wire new_AGEMA_signal_13885 ;
    wire new_AGEMA_signal_13886 ;
    wire new_AGEMA_signal_13887 ;
    wire new_AGEMA_signal_13888 ;
    wire new_AGEMA_signal_13889 ;
    wire new_AGEMA_signal_13890 ;
    wire new_AGEMA_signal_13891 ;
    wire new_AGEMA_signal_13892 ;
    wire new_AGEMA_signal_13893 ;
    wire new_AGEMA_signal_13894 ;
    wire new_AGEMA_signal_13895 ;
    wire new_AGEMA_signal_13896 ;
    wire new_AGEMA_signal_13897 ;
    wire new_AGEMA_signal_13898 ;
    wire new_AGEMA_signal_13899 ;
    wire new_AGEMA_signal_13900 ;
    wire new_AGEMA_signal_13901 ;
    wire new_AGEMA_signal_13902 ;
    wire new_AGEMA_signal_13903 ;
    wire new_AGEMA_signal_13904 ;
    wire new_AGEMA_signal_13905 ;
    wire new_AGEMA_signal_13906 ;
    wire new_AGEMA_signal_13907 ;
    wire new_AGEMA_signal_13908 ;
    wire new_AGEMA_signal_13909 ;
    wire new_AGEMA_signal_13910 ;
    wire new_AGEMA_signal_13911 ;
    wire new_AGEMA_signal_13912 ;
    wire new_AGEMA_signal_13913 ;
    wire new_AGEMA_signal_13914 ;
    wire new_AGEMA_signal_13915 ;
    wire new_AGEMA_signal_13916 ;
    wire new_AGEMA_signal_13917 ;
    wire new_AGEMA_signal_13918 ;
    wire new_AGEMA_signal_13919 ;
    wire new_AGEMA_signal_13920 ;
    wire new_AGEMA_signal_13921 ;
    wire new_AGEMA_signal_13922 ;
    wire new_AGEMA_signal_13923 ;
    wire new_AGEMA_signal_13924 ;
    wire new_AGEMA_signal_13925 ;
    wire new_AGEMA_signal_13926 ;
    wire new_AGEMA_signal_13927 ;
    wire new_AGEMA_signal_13928 ;
    wire new_AGEMA_signal_13929 ;
    wire new_AGEMA_signal_13930 ;
    wire new_AGEMA_signal_13931 ;
    wire new_AGEMA_signal_13932 ;
    wire new_AGEMA_signal_13933 ;
    wire new_AGEMA_signal_13934 ;
    wire new_AGEMA_signal_13935 ;
    wire new_AGEMA_signal_13936 ;
    wire new_AGEMA_signal_13937 ;
    wire new_AGEMA_signal_13938 ;
    wire new_AGEMA_signal_13939 ;
    wire new_AGEMA_signal_13940 ;
    wire new_AGEMA_signal_13941 ;
    wire new_AGEMA_signal_13942 ;
    wire new_AGEMA_signal_13943 ;
    wire new_AGEMA_signal_13944 ;
    wire new_AGEMA_signal_13945 ;
    wire new_AGEMA_signal_13946 ;
    wire new_AGEMA_signal_13947 ;
    wire new_AGEMA_signal_13948 ;
    wire new_AGEMA_signal_13949 ;
    wire new_AGEMA_signal_13950 ;
    wire new_AGEMA_signal_13951 ;
    wire new_AGEMA_signal_13952 ;
    wire new_AGEMA_signal_13953 ;
    wire new_AGEMA_signal_13954 ;
    wire new_AGEMA_signal_13955 ;
    wire new_AGEMA_signal_13956 ;
    wire new_AGEMA_signal_13957 ;
    wire new_AGEMA_signal_13958 ;
    wire new_AGEMA_signal_13959 ;
    wire new_AGEMA_signal_13960 ;
    wire new_AGEMA_signal_13961 ;
    wire new_AGEMA_signal_13962 ;
    wire new_AGEMA_signal_13963 ;
    wire new_AGEMA_signal_13964 ;
    wire new_AGEMA_signal_13965 ;
    wire new_AGEMA_signal_13966 ;
    wire new_AGEMA_signal_13967 ;
    wire new_AGEMA_signal_13968 ;
    wire new_AGEMA_signal_13969 ;
    wire new_AGEMA_signal_13970 ;
    wire new_AGEMA_signal_13971 ;
    wire new_AGEMA_signal_13972 ;
    wire new_AGEMA_signal_13973 ;
    wire new_AGEMA_signal_13974 ;
    wire new_AGEMA_signal_13975 ;
    wire new_AGEMA_signal_13976 ;
    wire new_AGEMA_signal_13977 ;
    wire new_AGEMA_signal_13978 ;
    wire new_AGEMA_signal_13979 ;
    wire new_AGEMA_signal_13980 ;
    wire new_AGEMA_signal_13981 ;
    wire new_AGEMA_signal_13982 ;
    wire new_AGEMA_signal_13983 ;
    wire new_AGEMA_signal_13984 ;
    wire new_AGEMA_signal_13985 ;
    wire new_AGEMA_signal_13986 ;
    wire new_AGEMA_signal_13987 ;
    wire new_AGEMA_signal_13988 ;
    wire new_AGEMA_signal_13989 ;
    wire new_AGEMA_signal_13990 ;
    wire new_AGEMA_signal_13991 ;
    wire new_AGEMA_signal_13992 ;
    wire new_AGEMA_signal_13993 ;
    wire new_AGEMA_signal_13994 ;
    wire new_AGEMA_signal_13995 ;
    wire new_AGEMA_signal_13996 ;
    wire new_AGEMA_signal_13997 ;
    wire new_AGEMA_signal_13998 ;
    wire new_AGEMA_signal_13999 ;
    wire new_AGEMA_signal_14000 ;
    wire new_AGEMA_signal_14001 ;
    wire new_AGEMA_signal_14002 ;
    wire new_AGEMA_signal_14003 ;
    wire new_AGEMA_signal_14004 ;
    wire new_AGEMA_signal_14005 ;
    wire new_AGEMA_signal_14006 ;
    wire new_AGEMA_signal_14007 ;
    wire new_AGEMA_signal_14008 ;
    wire new_AGEMA_signal_14009 ;
    wire new_AGEMA_signal_14010 ;
    wire new_AGEMA_signal_14011 ;
    wire new_AGEMA_signal_14012 ;
    wire new_AGEMA_signal_14013 ;
    wire new_AGEMA_signal_14014 ;
    wire new_AGEMA_signal_14015 ;
    wire new_AGEMA_signal_14016 ;
    wire new_AGEMA_signal_14017 ;
    wire new_AGEMA_signal_14018 ;
    wire new_AGEMA_signal_14019 ;
    wire new_AGEMA_signal_14020 ;
    wire new_AGEMA_signal_14021 ;
    wire new_AGEMA_signal_14022 ;
    wire new_AGEMA_signal_14023 ;
    wire new_AGEMA_signal_14024 ;
    wire new_AGEMA_signal_14025 ;
    wire new_AGEMA_signal_14026 ;
    wire new_AGEMA_signal_14027 ;
    wire new_AGEMA_signal_14028 ;
    wire new_AGEMA_signal_14029 ;
    wire new_AGEMA_signal_14030 ;
    wire new_AGEMA_signal_14031 ;
    wire new_AGEMA_signal_14032 ;
    wire new_AGEMA_signal_14033 ;
    wire new_AGEMA_signal_14034 ;
    wire new_AGEMA_signal_14035 ;
    wire new_AGEMA_signal_14036 ;
    wire new_AGEMA_signal_14037 ;
    wire new_AGEMA_signal_14038 ;
    wire new_AGEMA_signal_14039 ;
    wire new_AGEMA_signal_14040 ;
    wire new_AGEMA_signal_14041 ;
    wire new_AGEMA_signal_14042 ;
    wire new_AGEMA_signal_14043 ;
    wire new_AGEMA_signal_14044 ;
    wire new_AGEMA_signal_14045 ;
    wire new_AGEMA_signal_14046 ;
    wire new_AGEMA_signal_14047 ;
    wire new_AGEMA_signal_14048 ;
    wire new_AGEMA_signal_14049 ;
    wire new_AGEMA_signal_14050 ;
    wire new_AGEMA_signal_14051 ;
    wire new_AGEMA_signal_14052 ;
    wire new_AGEMA_signal_14053 ;
    wire new_AGEMA_signal_14054 ;
    wire new_AGEMA_signal_14055 ;
    wire new_AGEMA_signal_14056 ;
    wire new_AGEMA_signal_14057 ;
    wire new_AGEMA_signal_14058 ;
    wire new_AGEMA_signal_14059 ;
    wire new_AGEMA_signal_14060 ;
    wire new_AGEMA_signal_14061 ;
    wire new_AGEMA_signal_14062 ;
    wire new_AGEMA_signal_14063 ;
    wire new_AGEMA_signal_14064 ;
    wire new_AGEMA_signal_14065 ;
    wire new_AGEMA_signal_14066 ;
    wire new_AGEMA_signal_14067 ;
    wire new_AGEMA_signal_14068 ;
    wire new_AGEMA_signal_14069 ;
    wire new_AGEMA_signal_14070 ;
    wire new_AGEMA_signal_14071 ;
    wire new_AGEMA_signal_14072 ;
    wire new_AGEMA_signal_14073 ;
    wire new_AGEMA_signal_14074 ;
    wire new_AGEMA_signal_14075 ;
    wire new_AGEMA_signal_14076 ;
    wire new_AGEMA_signal_14077 ;
    wire new_AGEMA_signal_14078 ;
    wire new_AGEMA_signal_14079 ;
    wire new_AGEMA_signal_14080 ;
    wire new_AGEMA_signal_14081 ;
    wire new_AGEMA_signal_14082 ;
    wire new_AGEMA_signal_14083 ;
    wire new_AGEMA_signal_14084 ;
    wire new_AGEMA_signal_14085 ;
    wire new_AGEMA_signal_14086 ;
    wire new_AGEMA_signal_14087 ;
    wire new_AGEMA_signal_14088 ;
    wire new_AGEMA_signal_14089 ;
    wire new_AGEMA_signal_14090 ;
    wire new_AGEMA_signal_14091 ;
    wire new_AGEMA_signal_14092 ;
    wire new_AGEMA_signal_14093 ;
    wire new_AGEMA_signal_14094 ;
    wire new_AGEMA_signal_14095 ;
    wire new_AGEMA_signal_14096 ;
    wire new_AGEMA_signal_14097 ;
    wire new_AGEMA_signal_14098 ;
    wire new_AGEMA_signal_14099 ;
    wire new_AGEMA_signal_14100 ;
    wire new_AGEMA_signal_14101 ;
    wire new_AGEMA_signal_14102 ;
    wire new_AGEMA_signal_14103 ;
    wire new_AGEMA_signal_14104 ;
    wire new_AGEMA_signal_14105 ;
    wire new_AGEMA_signal_14106 ;
    wire new_AGEMA_signal_14107 ;
    wire new_AGEMA_signal_14108 ;
    wire new_AGEMA_signal_14109 ;
    wire new_AGEMA_signal_14110 ;
    wire new_AGEMA_signal_14111 ;
    wire new_AGEMA_signal_14112 ;
    wire new_AGEMA_signal_14113 ;
    wire new_AGEMA_signal_14114 ;
    wire new_AGEMA_signal_14115 ;
    wire new_AGEMA_signal_14116 ;
    wire new_AGEMA_signal_14117 ;
    wire new_AGEMA_signal_14118 ;
    wire new_AGEMA_signal_14119 ;
    wire new_AGEMA_signal_14120 ;
    wire new_AGEMA_signal_14121 ;
    wire new_AGEMA_signal_14122 ;
    wire new_AGEMA_signal_14123 ;
    wire new_AGEMA_signal_14124 ;
    wire new_AGEMA_signal_14125 ;
    wire new_AGEMA_signal_14126 ;
    wire new_AGEMA_signal_14127 ;
    wire new_AGEMA_signal_14128 ;
    wire new_AGEMA_signal_14129 ;
    wire new_AGEMA_signal_14130 ;
    wire new_AGEMA_signal_14131 ;
    wire new_AGEMA_signal_14132 ;
    wire new_AGEMA_signal_14133 ;
    wire new_AGEMA_signal_14134 ;
    wire new_AGEMA_signal_14135 ;
    wire new_AGEMA_signal_14136 ;
    wire new_AGEMA_signal_14137 ;
    wire new_AGEMA_signal_14138 ;
    wire new_AGEMA_signal_14139 ;
    wire new_AGEMA_signal_14140 ;
    wire new_AGEMA_signal_14141 ;
    wire new_AGEMA_signal_14142 ;
    wire new_AGEMA_signal_14143 ;
    wire new_AGEMA_signal_14144 ;
    wire new_AGEMA_signal_14145 ;
    wire new_AGEMA_signal_14146 ;
    wire new_AGEMA_signal_14147 ;
    wire new_AGEMA_signal_14148 ;
    wire new_AGEMA_signal_14149 ;
    wire new_AGEMA_signal_14150 ;
    wire new_AGEMA_signal_14151 ;
    wire new_AGEMA_signal_14152 ;
    wire new_AGEMA_signal_14153 ;
    wire new_AGEMA_signal_14154 ;
    wire new_AGEMA_signal_14155 ;
    wire new_AGEMA_signal_14156 ;
    wire new_AGEMA_signal_14157 ;
    wire new_AGEMA_signal_14158 ;
    wire new_AGEMA_signal_14159 ;
    wire new_AGEMA_signal_14160 ;
    wire new_AGEMA_signal_14161 ;
    wire new_AGEMA_signal_14162 ;
    wire new_AGEMA_signal_14163 ;
    wire new_AGEMA_signal_14164 ;
    wire new_AGEMA_signal_14165 ;
    wire new_AGEMA_signal_14166 ;
    wire new_AGEMA_signal_14167 ;
    wire new_AGEMA_signal_14168 ;
    wire new_AGEMA_signal_14169 ;
    wire new_AGEMA_signal_14170 ;
    wire new_AGEMA_signal_14171 ;
    wire new_AGEMA_signal_14172 ;
    wire new_AGEMA_signal_14173 ;
    wire new_AGEMA_signal_14174 ;
    wire new_AGEMA_signal_14175 ;
    wire new_AGEMA_signal_14176 ;
    wire new_AGEMA_signal_14177 ;
    wire new_AGEMA_signal_14178 ;
    wire new_AGEMA_signal_14179 ;
    wire new_AGEMA_signal_14180 ;
    wire new_AGEMA_signal_14181 ;
    wire new_AGEMA_signal_14182 ;
    wire new_AGEMA_signal_14183 ;
    wire new_AGEMA_signal_14184 ;
    wire new_AGEMA_signal_14185 ;
    wire new_AGEMA_signal_14186 ;
    wire new_AGEMA_signal_14187 ;
    wire new_AGEMA_signal_14188 ;
    wire new_AGEMA_signal_14189 ;
    wire new_AGEMA_signal_14190 ;
    wire new_AGEMA_signal_14191 ;
    wire new_AGEMA_signal_14192 ;
    wire new_AGEMA_signal_14193 ;
    wire new_AGEMA_signal_14194 ;
    wire new_AGEMA_signal_14195 ;
    wire new_AGEMA_signal_14196 ;
    wire new_AGEMA_signal_14197 ;
    wire new_AGEMA_signal_14198 ;
    wire new_AGEMA_signal_14199 ;
    wire new_AGEMA_signal_14200 ;
    wire new_AGEMA_signal_14201 ;
    wire new_AGEMA_signal_14202 ;
    wire new_AGEMA_signal_14203 ;
    wire new_AGEMA_signal_14204 ;
    wire new_AGEMA_signal_14205 ;
    wire new_AGEMA_signal_14206 ;
    wire new_AGEMA_signal_14207 ;
    wire new_AGEMA_signal_14208 ;
    wire new_AGEMA_signal_14209 ;
    wire new_AGEMA_signal_14210 ;
    wire new_AGEMA_signal_14211 ;
    wire new_AGEMA_signal_14212 ;
    wire new_AGEMA_signal_14213 ;
    wire new_AGEMA_signal_14214 ;
    wire new_AGEMA_signal_14215 ;
    wire new_AGEMA_signal_14216 ;
    wire new_AGEMA_signal_14217 ;
    wire new_AGEMA_signal_14218 ;
    wire new_AGEMA_signal_14219 ;
    wire new_AGEMA_signal_14220 ;
    wire new_AGEMA_signal_14221 ;
    wire new_AGEMA_signal_14222 ;
    wire new_AGEMA_signal_14223 ;
    wire new_AGEMA_signal_14224 ;
    wire new_AGEMA_signal_14225 ;
    wire new_AGEMA_signal_14226 ;
    wire new_AGEMA_signal_14227 ;
    wire new_AGEMA_signal_14228 ;
    wire new_AGEMA_signal_14229 ;
    wire new_AGEMA_signal_14230 ;
    wire new_AGEMA_signal_14231 ;
    wire new_AGEMA_signal_14232 ;
    wire new_AGEMA_signal_14233 ;
    wire new_AGEMA_signal_14234 ;
    wire new_AGEMA_signal_14235 ;
    wire new_AGEMA_signal_14236 ;
    wire new_AGEMA_signal_14237 ;
    wire new_AGEMA_signal_14238 ;
    wire new_AGEMA_signal_14239 ;
    wire new_AGEMA_signal_14240 ;
    wire new_AGEMA_signal_14241 ;
    wire new_AGEMA_signal_14242 ;
    wire new_AGEMA_signal_14243 ;
    wire new_AGEMA_signal_14244 ;
    wire new_AGEMA_signal_14245 ;
    wire new_AGEMA_signal_14246 ;
    wire new_AGEMA_signal_14247 ;
    wire new_AGEMA_signal_14248 ;
    wire new_AGEMA_signal_14249 ;
    wire new_AGEMA_signal_14250 ;
    wire new_AGEMA_signal_14251 ;
    wire new_AGEMA_signal_14252 ;
    wire new_AGEMA_signal_14253 ;
    wire new_AGEMA_signal_14254 ;
    wire new_AGEMA_signal_14255 ;
    wire new_AGEMA_signal_14256 ;
    wire new_AGEMA_signal_14257 ;
    wire new_AGEMA_signal_14258 ;
    wire new_AGEMA_signal_14259 ;
    wire new_AGEMA_signal_14260 ;
    wire new_AGEMA_signal_14261 ;
    wire new_AGEMA_signal_14262 ;
    wire new_AGEMA_signal_14263 ;
    wire new_AGEMA_signal_14264 ;
    wire new_AGEMA_signal_14265 ;
    wire new_AGEMA_signal_14266 ;
    wire new_AGEMA_signal_14267 ;
    wire new_AGEMA_signal_14268 ;
    wire new_AGEMA_signal_14269 ;
    wire new_AGEMA_signal_14270 ;
    wire new_AGEMA_signal_14271 ;
    wire new_AGEMA_signal_14272 ;
    wire new_AGEMA_signal_14273 ;
    wire new_AGEMA_signal_14274 ;
    wire new_AGEMA_signal_14275 ;
    wire new_AGEMA_signal_14276 ;
    wire new_AGEMA_signal_14277 ;
    wire new_AGEMA_signal_14278 ;
    wire new_AGEMA_signal_14279 ;
    wire new_AGEMA_signal_14280 ;
    wire new_AGEMA_signal_14281 ;
    wire new_AGEMA_signal_14282 ;
    wire new_AGEMA_signal_14283 ;
    wire new_AGEMA_signal_14284 ;
    wire new_AGEMA_signal_14285 ;
    wire new_AGEMA_signal_14286 ;
    wire new_AGEMA_signal_14287 ;
    wire new_AGEMA_signal_14288 ;
    wire new_AGEMA_signal_14289 ;
    wire new_AGEMA_signal_14290 ;
    wire new_AGEMA_signal_14291 ;
    wire new_AGEMA_signal_14292 ;
    wire new_AGEMA_signal_14293 ;
    wire new_AGEMA_signal_14294 ;
    wire new_AGEMA_signal_14295 ;
    wire new_AGEMA_signal_14296 ;
    wire new_AGEMA_signal_14297 ;
    wire new_AGEMA_signal_14298 ;
    wire new_AGEMA_signal_14299 ;
    wire new_AGEMA_signal_14300 ;
    wire new_AGEMA_signal_14301 ;
    wire new_AGEMA_signal_14302 ;
    wire new_AGEMA_signal_14303 ;
    wire new_AGEMA_signal_14304 ;
    wire new_AGEMA_signal_14305 ;
    wire new_AGEMA_signal_14306 ;
    wire new_AGEMA_signal_14307 ;
    wire new_AGEMA_signal_14308 ;
    wire new_AGEMA_signal_14309 ;
    wire new_AGEMA_signal_14310 ;
    wire new_AGEMA_signal_14311 ;
    wire new_AGEMA_signal_14312 ;
    wire new_AGEMA_signal_14313 ;
    wire new_AGEMA_signal_14314 ;
    wire new_AGEMA_signal_14315 ;
    wire new_AGEMA_signal_14316 ;
    wire new_AGEMA_signal_14317 ;
    wire new_AGEMA_signal_14318 ;
    wire new_AGEMA_signal_14319 ;
    wire new_AGEMA_signal_14320 ;
    wire new_AGEMA_signal_14321 ;
    wire new_AGEMA_signal_14322 ;
    wire new_AGEMA_signal_14323 ;
    wire new_AGEMA_signal_14324 ;
    wire new_AGEMA_signal_14325 ;
    wire new_AGEMA_signal_14326 ;
    wire new_AGEMA_signal_14327 ;
    wire new_AGEMA_signal_14328 ;
    wire new_AGEMA_signal_14329 ;
    wire new_AGEMA_signal_14330 ;
    wire new_AGEMA_signal_14331 ;
    wire new_AGEMA_signal_14332 ;
    wire new_AGEMA_signal_14333 ;
    wire new_AGEMA_signal_14334 ;
    wire new_AGEMA_signal_14335 ;
    wire new_AGEMA_signal_14336 ;
    wire new_AGEMA_signal_14337 ;
    wire new_AGEMA_signal_14338 ;
    wire new_AGEMA_signal_14339 ;
    wire new_AGEMA_signal_14340 ;
    wire new_AGEMA_signal_14341 ;
    wire new_AGEMA_signal_14342 ;
    wire new_AGEMA_signal_14343 ;
    wire new_AGEMA_signal_14344 ;
    wire new_AGEMA_signal_14345 ;
    wire new_AGEMA_signal_14346 ;
    wire new_AGEMA_signal_14347 ;
    wire new_AGEMA_signal_14348 ;
    wire new_AGEMA_signal_14349 ;
    wire new_AGEMA_signal_14350 ;
    wire new_AGEMA_signal_14351 ;
    wire new_AGEMA_signal_14352 ;
    wire new_AGEMA_signal_14353 ;
    wire new_AGEMA_signal_14354 ;
    wire new_AGEMA_signal_14355 ;
    wire new_AGEMA_signal_14356 ;
    wire new_AGEMA_signal_14357 ;
    wire new_AGEMA_signal_14358 ;
    wire new_AGEMA_signal_14359 ;
    wire new_AGEMA_signal_14360 ;
    wire new_AGEMA_signal_14361 ;
    wire new_AGEMA_signal_14362 ;
    wire new_AGEMA_signal_14363 ;
    wire new_AGEMA_signal_14364 ;
    wire new_AGEMA_signal_14365 ;
    wire new_AGEMA_signal_14366 ;
    wire new_AGEMA_signal_14367 ;
    wire new_AGEMA_signal_14368 ;
    wire new_AGEMA_signal_14369 ;
    wire new_AGEMA_signal_14370 ;
    wire new_AGEMA_signal_14371 ;
    wire new_AGEMA_signal_14372 ;
    wire new_AGEMA_signal_14373 ;
    wire new_AGEMA_signal_14374 ;
    wire new_AGEMA_signal_14375 ;
    wire new_AGEMA_signal_14376 ;
    wire new_AGEMA_signal_14377 ;
    wire new_AGEMA_signal_14378 ;
    wire new_AGEMA_signal_14379 ;
    wire new_AGEMA_signal_14380 ;
    wire new_AGEMA_signal_14381 ;
    wire new_AGEMA_signal_14382 ;
    wire new_AGEMA_signal_14383 ;
    wire new_AGEMA_signal_14384 ;
    wire new_AGEMA_signal_14385 ;
    wire new_AGEMA_signal_14386 ;
    wire new_AGEMA_signal_14387 ;
    wire new_AGEMA_signal_14388 ;
    wire new_AGEMA_signal_14389 ;
    wire new_AGEMA_signal_14390 ;
    wire new_AGEMA_signal_14391 ;
    wire new_AGEMA_signal_14392 ;
    wire new_AGEMA_signal_14393 ;
    wire new_AGEMA_signal_14394 ;
    wire new_AGEMA_signal_14395 ;
    wire new_AGEMA_signal_14396 ;
    wire new_AGEMA_signal_14397 ;
    wire new_AGEMA_signal_14398 ;
    wire new_AGEMA_signal_14399 ;
    wire new_AGEMA_signal_14400 ;
    wire new_AGEMA_signal_14401 ;
    wire new_AGEMA_signal_14402 ;
    wire new_AGEMA_signal_14403 ;
    wire new_AGEMA_signal_14404 ;
    wire new_AGEMA_signal_14405 ;
    wire new_AGEMA_signal_14406 ;
    wire new_AGEMA_signal_14407 ;
    wire new_AGEMA_signal_14408 ;
    wire new_AGEMA_signal_14409 ;
    wire new_AGEMA_signal_14410 ;
    wire new_AGEMA_signal_14411 ;
    wire new_AGEMA_signal_14412 ;
    wire new_AGEMA_signal_14413 ;
    wire new_AGEMA_signal_14414 ;
    wire new_AGEMA_signal_14415 ;
    wire new_AGEMA_signal_14416 ;
    wire new_AGEMA_signal_14417 ;
    wire new_AGEMA_signal_14418 ;
    wire new_AGEMA_signal_14419 ;
    wire new_AGEMA_signal_14420 ;
    wire new_AGEMA_signal_14421 ;
    wire new_AGEMA_signal_14422 ;
    wire new_AGEMA_signal_14423 ;
    wire new_AGEMA_signal_14424 ;
    wire new_AGEMA_signal_14425 ;
    wire new_AGEMA_signal_14426 ;
    wire new_AGEMA_signal_14427 ;
    wire new_AGEMA_signal_14428 ;
    wire new_AGEMA_signal_14429 ;
    wire new_AGEMA_signal_14430 ;
    wire new_AGEMA_signal_14431 ;
    wire new_AGEMA_signal_14432 ;
    wire new_AGEMA_signal_14433 ;
    wire new_AGEMA_signal_14434 ;
    wire new_AGEMA_signal_14435 ;
    wire new_AGEMA_signal_14436 ;
    wire new_AGEMA_signal_14437 ;
    wire new_AGEMA_signal_14438 ;
    wire new_AGEMA_signal_14439 ;
    wire new_AGEMA_signal_14440 ;
    wire new_AGEMA_signal_14441 ;
    wire new_AGEMA_signal_14442 ;
    wire new_AGEMA_signal_14443 ;
    wire new_AGEMA_signal_14444 ;
    wire new_AGEMA_signal_14445 ;
    wire new_AGEMA_signal_14446 ;
    wire new_AGEMA_signal_14447 ;
    wire new_AGEMA_signal_14448 ;
    wire new_AGEMA_signal_14449 ;
    wire new_AGEMA_signal_14450 ;
    wire new_AGEMA_signal_14451 ;
    wire new_AGEMA_signal_14452 ;
    wire new_AGEMA_signal_14453 ;
    wire new_AGEMA_signal_14454 ;
    wire new_AGEMA_signal_14455 ;
    wire new_AGEMA_signal_14456 ;
    wire new_AGEMA_signal_14457 ;
    wire new_AGEMA_signal_14458 ;
    wire new_AGEMA_signal_14459 ;
    wire new_AGEMA_signal_14460 ;
    wire new_AGEMA_signal_14461 ;
    wire new_AGEMA_signal_14462 ;
    wire new_AGEMA_signal_14463 ;
    wire new_AGEMA_signal_14464 ;
    wire new_AGEMA_signal_14465 ;
    wire new_AGEMA_signal_14466 ;
    wire new_AGEMA_signal_14467 ;
    wire new_AGEMA_signal_14468 ;
    wire new_AGEMA_signal_14469 ;
    wire new_AGEMA_signal_14470 ;
    wire new_AGEMA_signal_14471 ;
    wire new_AGEMA_signal_14472 ;
    wire new_AGEMA_signal_14473 ;
    wire new_AGEMA_signal_14474 ;
    wire new_AGEMA_signal_14475 ;
    wire new_AGEMA_signal_14476 ;
    wire new_AGEMA_signal_14477 ;
    wire new_AGEMA_signal_14478 ;
    wire new_AGEMA_signal_14479 ;
    wire new_AGEMA_signal_14480 ;
    wire new_AGEMA_signal_14481 ;
    wire new_AGEMA_signal_14482 ;
    wire new_AGEMA_signal_14483 ;
    wire new_AGEMA_signal_14484 ;
    wire new_AGEMA_signal_14485 ;
    wire new_AGEMA_signal_14486 ;
    wire new_AGEMA_signal_14487 ;
    wire new_AGEMA_signal_14488 ;
    wire new_AGEMA_signal_14489 ;
    wire new_AGEMA_signal_14490 ;
    wire new_AGEMA_signal_14491 ;
    wire new_AGEMA_signal_14492 ;
    wire new_AGEMA_signal_14493 ;
    wire new_AGEMA_signal_14494 ;
    wire new_AGEMA_signal_14495 ;
    wire new_AGEMA_signal_14496 ;
    wire new_AGEMA_signal_14497 ;
    wire new_AGEMA_signal_14498 ;
    wire new_AGEMA_signal_14499 ;
    wire new_AGEMA_signal_14500 ;
    wire new_AGEMA_signal_14501 ;
    wire new_AGEMA_signal_14502 ;
    wire new_AGEMA_signal_14503 ;
    wire new_AGEMA_signal_14504 ;
    wire new_AGEMA_signal_14505 ;
    wire new_AGEMA_signal_14506 ;
    wire new_AGEMA_signal_14507 ;
    wire new_AGEMA_signal_14508 ;
    wire new_AGEMA_signal_14509 ;
    wire new_AGEMA_signal_14510 ;
    wire new_AGEMA_signal_14511 ;
    wire new_AGEMA_signal_14512 ;
    wire new_AGEMA_signal_14513 ;
    wire new_AGEMA_signal_14514 ;
    wire new_AGEMA_signal_14515 ;
    wire new_AGEMA_signal_14516 ;
    wire new_AGEMA_signal_14517 ;
    wire new_AGEMA_signal_14518 ;
    wire new_AGEMA_signal_14519 ;
    wire new_AGEMA_signal_14520 ;
    wire new_AGEMA_signal_14521 ;
    wire new_AGEMA_signal_14522 ;
    wire new_AGEMA_signal_14523 ;
    wire new_AGEMA_signal_14524 ;
    wire new_AGEMA_signal_14525 ;
    wire new_AGEMA_signal_14526 ;
    wire new_AGEMA_signal_14527 ;
    wire new_AGEMA_signal_14528 ;
    wire new_AGEMA_signal_14529 ;
    wire new_AGEMA_signal_14530 ;
    wire new_AGEMA_signal_14531 ;
    wire new_AGEMA_signal_14532 ;
    wire new_AGEMA_signal_14533 ;
    wire new_AGEMA_signal_14534 ;
    wire new_AGEMA_signal_14535 ;
    wire new_AGEMA_signal_14536 ;
    wire new_AGEMA_signal_14537 ;
    wire new_AGEMA_signal_14538 ;
    wire new_AGEMA_signal_14539 ;
    wire new_AGEMA_signal_14540 ;
    wire new_AGEMA_signal_14541 ;
    wire new_AGEMA_signal_14542 ;
    wire new_AGEMA_signal_14543 ;
    wire new_AGEMA_signal_14544 ;
    wire new_AGEMA_signal_14545 ;
    wire new_AGEMA_signal_14546 ;
    wire new_AGEMA_signal_14547 ;
    wire new_AGEMA_signal_14548 ;
    wire new_AGEMA_signal_14549 ;
    wire new_AGEMA_signal_14550 ;
    wire new_AGEMA_signal_14551 ;
    wire new_AGEMA_signal_14552 ;
    wire new_AGEMA_signal_14553 ;
    wire new_AGEMA_signal_14554 ;
    wire new_AGEMA_signal_14555 ;
    wire new_AGEMA_signal_14556 ;
    wire new_AGEMA_signal_14557 ;
    wire new_AGEMA_signal_14558 ;
    wire new_AGEMA_signal_14559 ;
    wire new_AGEMA_signal_14560 ;
    wire new_AGEMA_signal_14561 ;
    wire new_AGEMA_signal_14562 ;
    wire new_AGEMA_signal_14563 ;
    wire new_AGEMA_signal_14564 ;
    wire new_AGEMA_signal_14565 ;
    wire new_AGEMA_signal_14566 ;
    wire new_AGEMA_signal_14567 ;
    wire new_AGEMA_signal_14568 ;
    wire new_AGEMA_signal_14569 ;
    wire new_AGEMA_signal_14570 ;
    wire new_AGEMA_signal_14571 ;
    wire new_AGEMA_signal_14572 ;
    wire new_AGEMA_signal_14573 ;
    wire new_AGEMA_signal_14574 ;
    wire new_AGEMA_signal_14575 ;
    wire new_AGEMA_signal_14576 ;
    wire new_AGEMA_signal_14577 ;
    wire new_AGEMA_signal_14578 ;
    wire new_AGEMA_signal_14579 ;
    wire new_AGEMA_signal_14580 ;
    wire new_AGEMA_signal_14581 ;
    wire new_AGEMA_signal_14582 ;
    wire new_AGEMA_signal_14583 ;
    wire new_AGEMA_signal_14584 ;
    wire new_AGEMA_signal_14585 ;
    wire new_AGEMA_signal_14586 ;
    wire new_AGEMA_signal_14587 ;
    wire new_AGEMA_signal_14588 ;
    wire new_AGEMA_signal_14589 ;
    wire new_AGEMA_signal_14590 ;
    wire new_AGEMA_signal_14591 ;
    wire new_AGEMA_signal_14592 ;
    wire new_AGEMA_signal_14593 ;
    wire new_AGEMA_signal_14594 ;
    wire new_AGEMA_signal_14595 ;
    wire new_AGEMA_signal_14596 ;
    wire new_AGEMA_signal_14597 ;
    wire new_AGEMA_signal_14598 ;
    wire new_AGEMA_signal_14599 ;
    wire new_AGEMA_signal_14600 ;
    wire new_AGEMA_signal_14601 ;
    wire new_AGEMA_signal_14602 ;
    wire new_AGEMA_signal_14603 ;
    wire new_AGEMA_signal_14604 ;
    wire new_AGEMA_signal_14605 ;
    wire new_AGEMA_signal_14606 ;
    wire new_AGEMA_signal_14607 ;
    wire new_AGEMA_signal_14608 ;
    wire new_AGEMA_signal_14609 ;
    wire new_AGEMA_signal_14610 ;
    wire new_AGEMA_signal_14611 ;
    wire new_AGEMA_signal_14612 ;
    wire new_AGEMA_signal_14613 ;
    wire new_AGEMA_signal_14614 ;
    wire new_AGEMA_signal_14615 ;
    wire new_AGEMA_signal_14616 ;
    wire new_AGEMA_signal_14617 ;
    wire new_AGEMA_signal_14618 ;
    wire new_AGEMA_signal_14619 ;
    wire new_AGEMA_signal_14620 ;
    wire new_AGEMA_signal_14621 ;
    wire new_AGEMA_signal_14622 ;
    wire new_AGEMA_signal_14623 ;
    wire new_AGEMA_signal_14624 ;
    wire new_AGEMA_signal_14625 ;
    wire new_AGEMA_signal_14626 ;
    wire new_AGEMA_signal_14627 ;
    wire new_AGEMA_signal_14628 ;
    wire new_AGEMA_signal_14629 ;
    wire new_AGEMA_signal_14630 ;
    wire new_AGEMA_signal_14631 ;
    wire new_AGEMA_signal_14632 ;
    wire new_AGEMA_signal_14633 ;
    wire new_AGEMA_signal_14634 ;
    wire new_AGEMA_signal_14635 ;
    wire new_AGEMA_signal_14636 ;
    wire new_AGEMA_signal_14637 ;
    wire new_AGEMA_signal_14638 ;
    wire new_AGEMA_signal_14639 ;
    wire new_AGEMA_signal_14640 ;
    wire new_AGEMA_signal_14641 ;
    wire new_AGEMA_signal_14642 ;
    wire new_AGEMA_signal_14643 ;
    wire new_AGEMA_signal_14644 ;
    wire new_AGEMA_signal_14645 ;
    wire new_AGEMA_signal_14646 ;
    wire new_AGEMA_signal_14647 ;
    wire new_AGEMA_signal_14648 ;
    wire new_AGEMA_signal_14649 ;
    wire new_AGEMA_signal_14650 ;
    wire new_AGEMA_signal_14651 ;
    wire new_AGEMA_signal_14652 ;
    wire new_AGEMA_signal_14653 ;
    wire new_AGEMA_signal_14654 ;
    wire new_AGEMA_signal_14655 ;
    wire new_AGEMA_signal_14656 ;
    wire new_AGEMA_signal_14657 ;
    wire new_AGEMA_signal_14658 ;
    wire new_AGEMA_signal_14659 ;
    wire new_AGEMA_signal_14660 ;
    wire new_AGEMA_signal_14661 ;
    wire new_AGEMA_signal_14662 ;
    wire new_AGEMA_signal_14663 ;
    wire new_AGEMA_signal_14664 ;
    wire new_AGEMA_signal_14665 ;
    wire new_AGEMA_signal_14666 ;
    wire new_AGEMA_signal_14667 ;
    wire new_AGEMA_signal_14668 ;
    wire new_AGEMA_signal_14669 ;
    wire new_AGEMA_signal_14670 ;
    wire new_AGEMA_signal_14671 ;
    wire new_AGEMA_signal_14672 ;
    wire new_AGEMA_signal_14673 ;
    wire new_AGEMA_signal_14674 ;
    wire new_AGEMA_signal_14675 ;
    wire new_AGEMA_signal_14676 ;
    wire new_AGEMA_signal_14677 ;
    wire new_AGEMA_signal_14678 ;
    wire new_AGEMA_signal_14679 ;
    wire new_AGEMA_signal_14680 ;
    wire new_AGEMA_signal_14681 ;
    wire new_AGEMA_signal_14682 ;
    wire new_AGEMA_signal_14683 ;
    wire new_AGEMA_signal_14684 ;
    wire new_AGEMA_signal_14685 ;
    wire new_AGEMA_signal_14686 ;
    wire new_AGEMA_signal_14687 ;
    wire new_AGEMA_signal_14688 ;
    wire new_AGEMA_signal_14689 ;
    wire new_AGEMA_signal_14690 ;
    wire new_AGEMA_signal_14691 ;
    wire new_AGEMA_signal_14692 ;
    wire new_AGEMA_signal_14693 ;
    wire new_AGEMA_signal_14694 ;
    wire new_AGEMA_signal_14695 ;
    wire new_AGEMA_signal_14696 ;
    wire new_AGEMA_signal_14697 ;
    wire new_AGEMA_signal_14698 ;
    wire new_AGEMA_signal_14699 ;
    wire new_AGEMA_signal_14700 ;
    wire new_AGEMA_signal_14701 ;
    wire new_AGEMA_signal_14702 ;
    wire new_AGEMA_signal_14703 ;
    wire new_AGEMA_signal_14704 ;
    wire new_AGEMA_signal_14705 ;
    wire new_AGEMA_signal_14706 ;
    wire new_AGEMA_signal_14707 ;
    wire new_AGEMA_signal_14708 ;
    wire new_AGEMA_signal_14709 ;
    wire new_AGEMA_signal_14710 ;
    wire new_AGEMA_signal_14711 ;
    wire new_AGEMA_signal_14712 ;
    wire new_AGEMA_signal_14713 ;
    wire new_AGEMA_signal_14714 ;
    wire new_AGEMA_signal_14715 ;
    wire new_AGEMA_signal_14716 ;
    wire new_AGEMA_signal_14717 ;
    wire new_AGEMA_signal_14718 ;
    wire new_AGEMA_signal_14719 ;
    wire new_AGEMA_signal_14720 ;
    wire new_AGEMA_signal_14721 ;
    wire new_AGEMA_signal_14722 ;
    wire new_AGEMA_signal_14723 ;
    wire new_AGEMA_signal_14724 ;
    wire new_AGEMA_signal_14725 ;
    wire new_AGEMA_signal_14726 ;
    wire new_AGEMA_signal_14727 ;
    wire new_AGEMA_signal_14728 ;
    wire new_AGEMA_signal_14729 ;
    wire new_AGEMA_signal_14730 ;
    wire new_AGEMA_signal_14731 ;
    wire new_AGEMA_signal_14732 ;
    wire new_AGEMA_signal_14733 ;
    wire new_AGEMA_signal_14734 ;
    wire new_AGEMA_signal_14735 ;
    wire new_AGEMA_signal_14736 ;
    wire new_AGEMA_signal_14737 ;
    wire new_AGEMA_signal_14738 ;
    wire new_AGEMA_signal_14739 ;
    wire new_AGEMA_signal_14740 ;
    wire new_AGEMA_signal_14741 ;
    wire new_AGEMA_signal_14742 ;
    wire new_AGEMA_signal_14743 ;
    wire new_AGEMA_signal_14744 ;
    wire new_AGEMA_signal_14745 ;
    wire new_AGEMA_signal_14746 ;
    wire new_AGEMA_signal_14747 ;
    wire new_AGEMA_signal_14748 ;
    wire new_AGEMA_signal_14749 ;
    wire new_AGEMA_signal_14750 ;
    wire new_AGEMA_signal_14751 ;
    wire new_AGEMA_signal_14752 ;
    wire new_AGEMA_signal_14753 ;
    wire new_AGEMA_signal_14754 ;
    wire new_AGEMA_signal_14755 ;
    wire new_AGEMA_signal_14756 ;
    wire new_AGEMA_signal_14757 ;
    wire new_AGEMA_signal_14758 ;
    wire new_AGEMA_signal_14759 ;
    wire new_AGEMA_signal_14760 ;
    wire new_AGEMA_signal_14761 ;
    wire new_AGEMA_signal_14762 ;
    wire new_AGEMA_signal_14763 ;
    wire new_AGEMA_signal_14764 ;
    wire new_AGEMA_signal_14765 ;
    wire new_AGEMA_signal_14766 ;
    wire new_AGEMA_signal_14767 ;
    wire new_AGEMA_signal_14768 ;
    wire new_AGEMA_signal_14769 ;
    wire new_AGEMA_signal_14770 ;
    wire new_AGEMA_signal_14771 ;
    wire new_AGEMA_signal_14772 ;
    wire new_AGEMA_signal_14773 ;
    wire new_AGEMA_signal_14774 ;
    wire new_AGEMA_signal_14775 ;
    wire new_AGEMA_signal_14776 ;
    wire new_AGEMA_signal_14777 ;
    wire new_AGEMA_signal_14778 ;
    wire new_AGEMA_signal_14779 ;
    wire new_AGEMA_signal_14780 ;
    wire new_AGEMA_signal_14781 ;
    wire new_AGEMA_signal_14782 ;
    wire new_AGEMA_signal_14783 ;
    wire new_AGEMA_signal_14784 ;
    wire new_AGEMA_signal_14785 ;
    wire new_AGEMA_signal_14786 ;
    wire new_AGEMA_signal_14787 ;
    wire new_AGEMA_signal_14788 ;
    wire new_AGEMA_signal_14789 ;
    wire new_AGEMA_signal_14790 ;
    wire new_AGEMA_signal_14791 ;
    wire new_AGEMA_signal_14792 ;
    wire new_AGEMA_signal_14793 ;
    wire new_AGEMA_signal_14794 ;
    wire new_AGEMA_signal_14795 ;
    wire new_AGEMA_signal_14796 ;
    wire new_AGEMA_signal_14797 ;
    wire new_AGEMA_signal_14798 ;
    wire new_AGEMA_signal_14799 ;
    wire new_AGEMA_signal_14800 ;
    wire new_AGEMA_signal_14801 ;
    wire new_AGEMA_signal_14802 ;
    wire new_AGEMA_signal_14803 ;
    wire new_AGEMA_signal_14804 ;
    wire new_AGEMA_signal_14805 ;
    wire new_AGEMA_signal_14806 ;
    wire new_AGEMA_signal_14807 ;
    wire new_AGEMA_signal_14808 ;
    wire new_AGEMA_signal_14809 ;
    wire new_AGEMA_signal_14810 ;
    wire new_AGEMA_signal_14811 ;
    wire new_AGEMA_signal_14812 ;
    wire new_AGEMA_signal_14813 ;
    wire new_AGEMA_signal_14814 ;
    wire new_AGEMA_signal_14815 ;
    wire new_AGEMA_signal_14816 ;
    wire new_AGEMA_signal_14817 ;
    wire new_AGEMA_signal_14818 ;
    wire new_AGEMA_signal_14819 ;
    wire new_AGEMA_signal_14820 ;
    wire new_AGEMA_signal_14821 ;
    wire new_AGEMA_signal_14822 ;
    wire new_AGEMA_signal_14823 ;
    wire new_AGEMA_signal_14824 ;
    wire new_AGEMA_signal_14825 ;
    wire new_AGEMA_signal_14826 ;
    wire new_AGEMA_signal_14827 ;
    wire new_AGEMA_signal_14828 ;
    wire new_AGEMA_signal_14829 ;
    wire new_AGEMA_signal_14830 ;
    wire new_AGEMA_signal_14831 ;
    wire new_AGEMA_signal_14832 ;
    wire new_AGEMA_signal_14833 ;
    wire new_AGEMA_signal_14834 ;
    wire new_AGEMA_signal_14835 ;
    wire new_AGEMA_signal_14836 ;
    wire new_AGEMA_signal_14837 ;
    wire new_AGEMA_signal_14838 ;
    wire new_AGEMA_signal_14839 ;
    wire new_AGEMA_signal_14840 ;
    wire new_AGEMA_signal_14841 ;
    wire new_AGEMA_signal_14842 ;
    wire new_AGEMA_signal_14843 ;
    wire new_AGEMA_signal_14844 ;
    wire new_AGEMA_signal_14845 ;
    wire new_AGEMA_signal_14846 ;
    wire new_AGEMA_signal_14847 ;
    wire new_AGEMA_signal_14848 ;
    wire new_AGEMA_signal_14849 ;
    wire new_AGEMA_signal_14850 ;
    wire new_AGEMA_signal_14851 ;
    wire new_AGEMA_signal_14852 ;
    wire new_AGEMA_signal_14853 ;
    wire new_AGEMA_signal_14854 ;
    wire new_AGEMA_signal_14855 ;
    wire new_AGEMA_signal_14856 ;
    wire new_AGEMA_signal_14857 ;
    wire new_AGEMA_signal_14858 ;
    wire new_AGEMA_signal_14859 ;
    wire new_AGEMA_signal_14860 ;
    wire new_AGEMA_signal_14861 ;
    wire new_AGEMA_signal_14862 ;
    wire new_AGEMA_signal_14863 ;
    wire new_AGEMA_signal_14864 ;
    wire new_AGEMA_signal_14865 ;
    wire new_AGEMA_signal_14866 ;
    wire new_AGEMA_signal_14867 ;
    wire new_AGEMA_signal_14868 ;
    wire new_AGEMA_signal_14869 ;
    wire new_AGEMA_signal_14870 ;
    wire new_AGEMA_signal_14871 ;
    wire new_AGEMA_signal_14872 ;
    wire new_AGEMA_signal_14873 ;
    wire new_AGEMA_signal_14874 ;
    wire new_AGEMA_signal_14875 ;
    wire new_AGEMA_signal_14876 ;
    wire new_AGEMA_signal_14877 ;
    wire new_AGEMA_signal_14878 ;
    wire new_AGEMA_signal_14879 ;
    wire new_AGEMA_signal_14880 ;
    wire new_AGEMA_signal_14881 ;
    wire new_AGEMA_signal_14882 ;
    wire new_AGEMA_signal_14883 ;
    wire new_AGEMA_signal_14884 ;
    wire new_AGEMA_signal_14885 ;
    wire new_AGEMA_signal_14886 ;
    wire new_AGEMA_signal_14887 ;
    wire new_AGEMA_signal_14888 ;
    wire new_AGEMA_signal_14889 ;
    wire new_AGEMA_signal_14890 ;
    wire new_AGEMA_signal_14891 ;
    wire new_AGEMA_signal_14892 ;
    wire new_AGEMA_signal_14893 ;
    wire new_AGEMA_signal_14894 ;
    wire new_AGEMA_signal_14895 ;
    wire new_AGEMA_signal_14896 ;
    wire new_AGEMA_signal_14897 ;
    wire new_AGEMA_signal_14898 ;
    wire new_AGEMA_signal_14899 ;
    wire new_AGEMA_signal_14900 ;
    wire new_AGEMA_signal_14901 ;
    wire new_AGEMA_signal_14902 ;
    wire new_AGEMA_signal_14903 ;
    wire new_AGEMA_signal_14904 ;
    wire new_AGEMA_signal_14905 ;
    wire new_AGEMA_signal_14906 ;
    wire new_AGEMA_signal_14907 ;
    wire new_AGEMA_signal_14908 ;
    wire new_AGEMA_signal_14909 ;
    wire new_AGEMA_signal_14910 ;
    wire new_AGEMA_signal_14911 ;
    wire new_AGEMA_signal_14912 ;
    wire new_AGEMA_signal_14913 ;
    wire new_AGEMA_signal_14914 ;
    wire new_AGEMA_signal_14915 ;
    wire new_AGEMA_signal_14916 ;
    wire new_AGEMA_signal_14917 ;
    wire new_AGEMA_signal_14918 ;
    wire new_AGEMA_signal_14919 ;
    wire new_AGEMA_signal_14920 ;
    wire new_AGEMA_signal_14921 ;
    wire new_AGEMA_signal_14922 ;
    wire new_AGEMA_signal_14923 ;
    wire new_AGEMA_signal_14924 ;
    wire new_AGEMA_signal_14925 ;
    wire new_AGEMA_signal_14926 ;
    wire new_AGEMA_signal_14927 ;
    wire new_AGEMA_signal_14928 ;
    wire new_AGEMA_signal_14929 ;
    wire new_AGEMA_signal_14930 ;
    wire new_AGEMA_signal_14931 ;
    wire new_AGEMA_signal_14932 ;
    wire new_AGEMA_signal_14933 ;
    wire new_AGEMA_signal_14934 ;
    wire new_AGEMA_signal_14935 ;
    wire new_AGEMA_signal_14936 ;
    wire new_AGEMA_signal_14937 ;
    wire new_AGEMA_signal_14938 ;
    wire new_AGEMA_signal_14939 ;
    wire new_AGEMA_signal_14940 ;
    wire new_AGEMA_signal_14941 ;
    wire new_AGEMA_signal_14942 ;
    wire new_AGEMA_signal_14943 ;
    wire new_AGEMA_signal_14944 ;
    wire new_AGEMA_signal_14945 ;
    wire new_AGEMA_signal_14946 ;
    wire new_AGEMA_signal_14947 ;
    wire new_AGEMA_signal_14948 ;
    wire new_AGEMA_signal_14949 ;
    wire new_AGEMA_signal_14950 ;
    wire new_AGEMA_signal_14951 ;
    wire new_AGEMA_signal_14952 ;
    wire new_AGEMA_signal_14953 ;
    wire new_AGEMA_signal_14954 ;
    wire new_AGEMA_signal_14955 ;
    wire new_AGEMA_signal_14956 ;
    wire new_AGEMA_signal_14957 ;
    wire new_AGEMA_signal_14958 ;
    wire new_AGEMA_signal_14959 ;
    wire new_AGEMA_signal_14960 ;
    wire new_AGEMA_signal_14961 ;
    wire new_AGEMA_signal_14962 ;
    wire new_AGEMA_signal_14963 ;
    wire new_AGEMA_signal_14964 ;
    wire new_AGEMA_signal_14965 ;
    wire new_AGEMA_signal_14966 ;
    wire new_AGEMA_signal_14967 ;
    wire new_AGEMA_signal_14968 ;
    wire new_AGEMA_signal_14969 ;
    wire new_AGEMA_signal_14970 ;
    wire new_AGEMA_signal_14971 ;
    wire new_AGEMA_signal_14972 ;
    wire new_AGEMA_signal_14973 ;
    wire new_AGEMA_signal_14974 ;
    wire new_AGEMA_signal_14975 ;
    wire new_AGEMA_signal_14976 ;
    wire new_AGEMA_signal_14977 ;
    wire new_AGEMA_signal_14978 ;
    wire new_AGEMA_signal_14979 ;
    wire new_AGEMA_signal_14980 ;
    wire new_AGEMA_signal_14981 ;
    wire new_AGEMA_signal_14982 ;
    wire new_AGEMA_signal_14983 ;
    wire new_AGEMA_signal_14984 ;
    wire new_AGEMA_signal_14985 ;
    wire new_AGEMA_signal_14986 ;
    wire new_AGEMA_signal_14987 ;
    wire new_AGEMA_signal_14988 ;
    wire new_AGEMA_signal_14989 ;
    wire new_AGEMA_signal_14990 ;
    wire new_AGEMA_signal_14991 ;
    wire new_AGEMA_signal_14992 ;
    wire new_AGEMA_signal_14993 ;
    wire new_AGEMA_signal_14994 ;
    wire new_AGEMA_signal_14995 ;
    wire new_AGEMA_signal_14996 ;
    wire new_AGEMA_signal_14997 ;
    wire new_AGEMA_signal_14998 ;
    wire new_AGEMA_signal_14999 ;
    wire new_AGEMA_signal_15000 ;
    wire new_AGEMA_signal_15001 ;
    wire new_AGEMA_signal_15002 ;
    wire new_AGEMA_signal_15003 ;
    wire new_AGEMA_signal_15004 ;
    wire new_AGEMA_signal_15005 ;
    wire new_AGEMA_signal_15006 ;
    wire new_AGEMA_signal_15007 ;
    wire new_AGEMA_signal_15008 ;
    wire new_AGEMA_signal_15009 ;
    wire new_AGEMA_signal_15010 ;
    wire new_AGEMA_signal_15011 ;
    wire new_AGEMA_signal_15012 ;
    wire new_AGEMA_signal_15013 ;
    wire new_AGEMA_signal_15014 ;
    wire new_AGEMA_signal_15015 ;
    wire new_AGEMA_signal_15016 ;
    wire new_AGEMA_signal_15017 ;
    wire new_AGEMA_signal_15018 ;
    wire new_AGEMA_signal_15019 ;
    wire new_AGEMA_signal_15020 ;
    wire new_AGEMA_signal_15021 ;
    wire new_AGEMA_signal_15022 ;
    wire new_AGEMA_signal_15023 ;
    wire new_AGEMA_signal_15024 ;
    wire new_AGEMA_signal_15025 ;
    wire new_AGEMA_signal_15026 ;
    wire new_AGEMA_signal_15027 ;
    wire new_AGEMA_signal_15028 ;
    wire new_AGEMA_signal_15029 ;
    wire new_AGEMA_signal_15030 ;
    wire new_AGEMA_signal_15031 ;
    wire new_AGEMA_signal_15032 ;
    wire new_AGEMA_signal_15033 ;
    wire new_AGEMA_signal_15034 ;
    wire new_AGEMA_signal_15035 ;
    wire new_AGEMA_signal_15036 ;
    wire new_AGEMA_signal_15037 ;
    wire new_AGEMA_signal_15038 ;
    wire new_AGEMA_signal_15039 ;
    wire new_AGEMA_signal_15040 ;
    wire new_AGEMA_signal_15041 ;
    wire new_AGEMA_signal_15042 ;
    wire new_AGEMA_signal_15043 ;
    wire new_AGEMA_signal_15044 ;
    wire new_AGEMA_signal_15045 ;
    wire new_AGEMA_signal_15046 ;
    wire new_AGEMA_signal_15047 ;
    wire new_AGEMA_signal_15048 ;
    wire new_AGEMA_signal_15049 ;
    wire new_AGEMA_signal_15050 ;
    wire new_AGEMA_signal_15051 ;
    wire new_AGEMA_signal_15052 ;
    wire new_AGEMA_signal_15053 ;
    wire new_AGEMA_signal_15054 ;
    wire new_AGEMA_signal_15055 ;
    wire new_AGEMA_signal_15056 ;
    wire new_AGEMA_signal_15057 ;
    wire new_AGEMA_signal_15058 ;
    wire new_AGEMA_signal_15059 ;
    wire new_AGEMA_signal_15060 ;
    wire new_AGEMA_signal_15061 ;
    wire new_AGEMA_signal_15062 ;
    wire new_AGEMA_signal_15063 ;
    wire new_AGEMA_signal_15064 ;
    wire new_AGEMA_signal_15065 ;
    wire new_AGEMA_signal_15066 ;
    wire new_AGEMA_signal_15067 ;
    wire new_AGEMA_signal_15068 ;
    wire new_AGEMA_signal_15069 ;
    wire new_AGEMA_signal_15070 ;
    wire new_AGEMA_signal_15071 ;
    wire new_AGEMA_signal_15072 ;
    wire new_AGEMA_signal_15073 ;
    wire new_AGEMA_signal_15074 ;
    wire new_AGEMA_signal_15075 ;
    wire new_AGEMA_signal_15076 ;
    wire new_AGEMA_signal_15077 ;
    wire new_AGEMA_signal_15078 ;
    wire new_AGEMA_signal_15079 ;
    wire new_AGEMA_signal_15080 ;
    wire new_AGEMA_signal_15081 ;
    wire new_AGEMA_signal_15082 ;
    wire new_AGEMA_signal_15083 ;
    wire new_AGEMA_signal_15084 ;
    wire new_AGEMA_signal_15085 ;
    wire new_AGEMA_signal_15086 ;
    wire new_AGEMA_signal_15087 ;
    wire new_AGEMA_signal_15088 ;
    wire new_AGEMA_signal_15089 ;
    wire new_AGEMA_signal_15090 ;
    wire new_AGEMA_signal_15091 ;
    wire new_AGEMA_signal_15092 ;
    wire new_AGEMA_signal_15093 ;
    wire new_AGEMA_signal_15094 ;
    wire new_AGEMA_signal_15095 ;
    wire new_AGEMA_signal_15096 ;
    wire new_AGEMA_signal_15097 ;
    wire new_AGEMA_signal_15098 ;
    wire new_AGEMA_signal_15099 ;
    wire new_AGEMA_signal_15100 ;
    wire new_AGEMA_signal_15101 ;
    wire new_AGEMA_signal_15102 ;
    wire new_AGEMA_signal_15103 ;
    wire new_AGEMA_signal_15104 ;
    wire new_AGEMA_signal_15105 ;
    wire new_AGEMA_signal_15106 ;
    wire new_AGEMA_signal_15107 ;
    wire new_AGEMA_signal_15108 ;
    wire new_AGEMA_signal_15109 ;
    wire new_AGEMA_signal_15110 ;
    wire new_AGEMA_signal_15111 ;
    wire new_AGEMA_signal_15112 ;
    wire new_AGEMA_signal_15113 ;
    wire new_AGEMA_signal_15114 ;
    wire new_AGEMA_signal_15115 ;
    wire new_AGEMA_signal_15116 ;
    wire new_AGEMA_signal_15117 ;
    wire new_AGEMA_signal_15118 ;
    wire new_AGEMA_signal_15119 ;
    wire new_AGEMA_signal_15120 ;
    wire new_AGEMA_signal_15121 ;
    wire new_AGEMA_signal_15122 ;
    wire new_AGEMA_signal_15123 ;
    wire new_AGEMA_signal_15124 ;
    wire new_AGEMA_signal_15125 ;
    wire new_AGEMA_signal_15126 ;
    wire new_AGEMA_signal_15127 ;
    wire new_AGEMA_signal_15128 ;
    wire new_AGEMA_signal_15129 ;
    wire new_AGEMA_signal_15130 ;
    wire new_AGEMA_signal_15131 ;
    wire new_AGEMA_signal_15132 ;
    wire new_AGEMA_signal_15133 ;
    wire new_AGEMA_signal_15134 ;
    wire new_AGEMA_signal_15135 ;
    wire new_AGEMA_signal_15136 ;
    wire new_AGEMA_signal_15137 ;
    wire new_AGEMA_signal_15138 ;
    wire new_AGEMA_signal_15139 ;
    wire new_AGEMA_signal_15140 ;
    wire new_AGEMA_signal_15141 ;
    wire new_AGEMA_signal_15142 ;
    wire new_AGEMA_signal_15143 ;
    wire new_AGEMA_signal_15144 ;
    wire new_AGEMA_signal_15145 ;
    wire new_AGEMA_signal_15146 ;
    wire new_AGEMA_signal_15147 ;
    wire new_AGEMA_signal_15148 ;
    wire new_AGEMA_signal_15149 ;
    wire new_AGEMA_signal_15150 ;
    wire new_AGEMA_signal_15151 ;
    wire new_AGEMA_signal_15152 ;
    wire new_AGEMA_signal_15153 ;
    wire new_AGEMA_signal_15154 ;
    wire new_AGEMA_signal_15155 ;
    wire new_AGEMA_signal_15156 ;
    wire new_AGEMA_signal_15157 ;
    wire new_AGEMA_signal_15158 ;
    wire new_AGEMA_signal_15159 ;
    wire new_AGEMA_signal_15160 ;
    wire new_AGEMA_signal_15161 ;
    wire new_AGEMA_signal_15162 ;
    wire new_AGEMA_signal_15163 ;
    wire new_AGEMA_signal_15164 ;
    wire new_AGEMA_signal_15165 ;
    wire new_AGEMA_signal_15166 ;
    wire new_AGEMA_signal_15167 ;
    wire new_AGEMA_signal_15168 ;
    wire new_AGEMA_signal_15169 ;
    wire new_AGEMA_signal_15170 ;
    wire new_AGEMA_signal_15171 ;
    wire new_AGEMA_signal_15172 ;
    wire new_AGEMA_signal_15173 ;
    wire new_AGEMA_signal_15174 ;
    wire new_AGEMA_signal_15175 ;
    wire new_AGEMA_signal_15176 ;
    wire new_AGEMA_signal_15177 ;
    wire new_AGEMA_signal_15178 ;
    wire new_AGEMA_signal_15179 ;
    wire new_AGEMA_signal_15180 ;
    wire new_AGEMA_signal_15181 ;
    wire new_AGEMA_signal_15182 ;
    wire new_AGEMA_signal_15183 ;
    wire new_AGEMA_signal_15184 ;
    wire new_AGEMA_signal_15185 ;
    wire new_AGEMA_signal_15186 ;
    wire new_AGEMA_signal_15187 ;
    wire new_AGEMA_signal_15188 ;
    wire new_AGEMA_signal_15189 ;
    wire new_AGEMA_signal_15190 ;
    wire new_AGEMA_signal_15191 ;
    wire new_AGEMA_signal_15192 ;
    wire new_AGEMA_signal_15193 ;
    wire new_AGEMA_signal_15194 ;
    wire new_AGEMA_signal_15195 ;
    wire new_AGEMA_signal_15196 ;
    wire new_AGEMA_signal_15197 ;
    wire new_AGEMA_signal_15198 ;
    wire new_AGEMA_signal_15199 ;
    wire new_AGEMA_signal_15200 ;
    wire new_AGEMA_signal_15201 ;
    wire new_AGEMA_signal_15202 ;
    wire new_AGEMA_signal_15203 ;
    wire new_AGEMA_signal_15204 ;
    wire new_AGEMA_signal_15205 ;
    wire new_AGEMA_signal_15206 ;
    wire new_AGEMA_signal_15207 ;
    wire new_AGEMA_signal_15208 ;
    wire new_AGEMA_signal_15209 ;
    wire new_AGEMA_signal_15210 ;
    wire new_AGEMA_signal_15211 ;
    wire new_AGEMA_signal_15212 ;
    wire new_AGEMA_signal_15213 ;
    wire new_AGEMA_signal_15214 ;
    wire new_AGEMA_signal_15215 ;
    wire new_AGEMA_signal_15216 ;
    wire new_AGEMA_signal_15217 ;
    wire new_AGEMA_signal_15218 ;
    wire new_AGEMA_signal_15219 ;
    wire new_AGEMA_signal_15220 ;
    wire new_AGEMA_signal_15221 ;
    wire new_AGEMA_signal_15222 ;
    wire new_AGEMA_signal_15223 ;
    wire new_AGEMA_signal_15224 ;
    wire new_AGEMA_signal_15225 ;
    wire new_AGEMA_signal_15226 ;
    wire new_AGEMA_signal_15227 ;
    wire new_AGEMA_signal_15228 ;
    wire new_AGEMA_signal_15229 ;
    wire new_AGEMA_signal_15230 ;
    wire new_AGEMA_signal_15231 ;
    wire new_AGEMA_signal_15232 ;
    wire new_AGEMA_signal_15233 ;
    wire new_AGEMA_signal_15234 ;
    wire new_AGEMA_signal_15235 ;
    wire new_AGEMA_signal_15236 ;
    wire new_AGEMA_signal_15237 ;
    wire new_AGEMA_signal_15238 ;
    wire new_AGEMA_signal_15239 ;
    wire new_AGEMA_signal_15240 ;
    wire new_AGEMA_signal_15241 ;
    wire new_AGEMA_signal_15242 ;
    wire new_AGEMA_signal_15243 ;
    wire new_AGEMA_signal_15244 ;
    wire new_AGEMA_signal_15245 ;
    wire new_AGEMA_signal_15246 ;
    wire new_AGEMA_signal_15247 ;
    wire new_AGEMA_signal_15248 ;
    wire new_AGEMA_signal_15249 ;
    wire new_AGEMA_signal_15250 ;
    wire new_AGEMA_signal_15251 ;
    wire new_AGEMA_signal_15252 ;
    wire new_AGEMA_signal_15253 ;
    wire new_AGEMA_signal_15254 ;
    wire new_AGEMA_signal_15255 ;
    wire new_AGEMA_signal_15256 ;
    wire new_AGEMA_signal_15257 ;
    wire new_AGEMA_signal_15258 ;
    wire new_AGEMA_signal_15259 ;
    wire new_AGEMA_signal_15260 ;
    wire new_AGEMA_signal_15261 ;
    wire new_AGEMA_signal_15262 ;
    wire new_AGEMA_signal_15263 ;
    wire new_AGEMA_signal_15264 ;
    wire new_AGEMA_signal_15265 ;
    wire new_AGEMA_signal_15266 ;
    wire new_AGEMA_signal_15267 ;
    wire new_AGEMA_signal_15268 ;
    wire new_AGEMA_signal_15269 ;
    wire new_AGEMA_signal_15270 ;
    wire new_AGEMA_signal_15271 ;
    wire new_AGEMA_signal_15272 ;
    wire new_AGEMA_signal_15273 ;
    wire new_AGEMA_signal_15274 ;
    wire new_AGEMA_signal_15275 ;
    wire new_AGEMA_signal_15276 ;
    wire new_AGEMA_signal_15277 ;
    wire new_AGEMA_signal_15278 ;
    wire new_AGEMA_signal_15279 ;
    wire new_AGEMA_signal_15280 ;
    wire new_AGEMA_signal_15281 ;
    wire new_AGEMA_signal_15282 ;
    wire new_AGEMA_signal_15283 ;
    wire new_AGEMA_signal_15284 ;
    wire new_AGEMA_signal_15285 ;
    wire new_AGEMA_signal_15286 ;
    wire new_AGEMA_signal_15287 ;
    wire new_AGEMA_signal_15288 ;
    wire new_AGEMA_signal_15289 ;
    wire new_AGEMA_signal_15290 ;
    wire new_AGEMA_signal_15291 ;
    wire new_AGEMA_signal_15292 ;
    wire new_AGEMA_signal_15293 ;
    wire new_AGEMA_signal_15294 ;
    wire new_AGEMA_signal_15295 ;
    wire new_AGEMA_signal_15296 ;
    wire new_AGEMA_signal_15297 ;
    wire new_AGEMA_signal_15298 ;
    wire new_AGEMA_signal_15299 ;
    wire new_AGEMA_signal_15300 ;
    wire new_AGEMA_signal_15301 ;
    wire new_AGEMA_signal_15302 ;
    wire new_AGEMA_signal_15303 ;
    wire new_AGEMA_signal_15304 ;
    wire new_AGEMA_signal_15305 ;
    wire new_AGEMA_signal_15306 ;
    wire new_AGEMA_signal_15307 ;
    wire new_AGEMA_signal_15308 ;
    wire new_AGEMA_signal_15309 ;
    wire new_AGEMA_signal_15310 ;
    wire new_AGEMA_signal_15311 ;
    wire new_AGEMA_signal_15312 ;
    wire new_AGEMA_signal_15313 ;
    wire new_AGEMA_signal_15314 ;
    wire new_AGEMA_signal_15315 ;
    wire new_AGEMA_signal_15316 ;
    wire new_AGEMA_signal_15317 ;
    wire new_AGEMA_signal_15318 ;
    wire new_AGEMA_signal_15319 ;
    wire new_AGEMA_signal_15320 ;
    wire new_AGEMA_signal_15321 ;
    wire new_AGEMA_signal_15322 ;
    wire new_AGEMA_signal_15323 ;
    wire new_AGEMA_signal_15324 ;
    wire new_AGEMA_signal_15325 ;
    wire new_AGEMA_signal_15326 ;
    wire new_AGEMA_signal_15327 ;
    wire new_AGEMA_signal_15328 ;
    wire new_AGEMA_signal_15329 ;
    wire new_AGEMA_signal_15330 ;
    wire new_AGEMA_signal_15331 ;
    wire new_AGEMA_signal_15332 ;
    wire new_AGEMA_signal_15333 ;
    wire new_AGEMA_signal_15334 ;
    wire new_AGEMA_signal_15335 ;
    wire new_AGEMA_signal_15336 ;
    wire new_AGEMA_signal_15337 ;
    wire new_AGEMA_signal_15338 ;
    wire new_AGEMA_signal_15339 ;
    wire new_AGEMA_signal_15340 ;
    wire new_AGEMA_signal_15341 ;
    wire new_AGEMA_signal_15342 ;
    wire new_AGEMA_signal_15343 ;
    wire new_AGEMA_signal_15344 ;
    wire new_AGEMA_signal_15345 ;
    wire new_AGEMA_signal_15346 ;
    wire new_AGEMA_signal_15347 ;
    wire new_AGEMA_signal_15348 ;
    wire new_AGEMA_signal_15349 ;
    wire new_AGEMA_signal_15350 ;
    wire new_AGEMA_signal_15351 ;
    wire new_AGEMA_signal_15352 ;
    wire new_AGEMA_signal_15353 ;
    wire new_AGEMA_signal_15354 ;
    wire new_AGEMA_signal_15355 ;
    wire new_AGEMA_signal_15356 ;
    wire new_AGEMA_signal_15357 ;
    wire new_AGEMA_signal_15358 ;
    wire new_AGEMA_signal_15359 ;
    wire new_AGEMA_signal_15360 ;
    wire new_AGEMA_signal_15361 ;
    wire new_AGEMA_signal_15362 ;
    wire new_AGEMA_signal_15363 ;
    wire new_AGEMA_signal_15364 ;
    wire new_AGEMA_signal_15365 ;
    wire new_AGEMA_signal_15366 ;
    wire new_AGEMA_signal_15367 ;
    wire new_AGEMA_signal_15368 ;
    wire new_AGEMA_signal_15369 ;
    wire new_AGEMA_signal_15370 ;
    wire new_AGEMA_signal_15371 ;
    wire new_AGEMA_signal_15372 ;
    wire new_AGEMA_signal_15373 ;
    wire new_AGEMA_signal_15374 ;
    wire new_AGEMA_signal_15375 ;
    wire new_AGEMA_signal_15376 ;
    wire new_AGEMA_signal_15377 ;
    wire new_AGEMA_signal_15378 ;
    wire new_AGEMA_signal_15379 ;
    wire new_AGEMA_signal_15380 ;
    wire new_AGEMA_signal_15381 ;
    wire new_AGEMA_signal_15382 ;
    wire new_AGEMA_signal_15383 ;
    wire new_AGEMA_signal_15384 ;
    wire new_AGEMA_signal_15385 ;
    wire new_AGEMA_signal_15386 ;
    wire new_AGEMA_signal_15387 ;
    wire new_AGEMA_signal_15388 ;
    wire new_AGEMA_signal_15389 ;
    wire new_AGEMA_signal_15390 ;
    wire new_AGEMA_signal_15391 ;
    wire new_AGEMA_signal_15392 ;
    wire new_AGEMA_signal_15393 ;
    wire new_AGEMA_signal_15394 ;
    wire new_AGEMA_signal_15395 ;
    wire new_AGEMA_signal_15396 ;
    wire new_AGEMA_signal_15397 ;
    wire new_AGEMA_signal_15398 ;
    wire new_AGEMA_signal_15399 ;
    wire new_AGEMA_signal_15400 ;
    wire new_AGEMA_signal_15401 ;
    wire new_AGEMA_signal_15402 ;
    wire new_AGEMA_signal_15403 ;
    wire new_AGEMA_signal_15404 ;
    wire new_AGEMA_signal_15405 ;
    wire new_AGEMA_signal_15406 ;
    wire new_AGEMA_signal_15407 ;
    wire new_AGEMA_signal_15408 ;
    wire new_AGEMA_signal_15409 ;
    wire new_AGEMA_signal_15410 ;
    wire new_AGEMA_signal_15411 ;
    wire new_AGEMA_signal_15412 ;
    wire new_AGEMA_signal_15413 ;
    wire new_AGEMA_signal_15414 ;
    wire new_AGEMA_signal_15415 ;
    wire new_AGEMA_signal_15416 ;
    wire new_AGEMA_signal_15417 ;
    wire new_AGEMA_signal_15418 ;
    wire new_AGEMA_signal_15419 ;
    wire new_AGEMA_signal_15420 ;
    wire new_AGEMA_signal_15421 ;
    wire new_AGEMA_signal_15422 ;
    wire new_AGEMA_signal_15423 ;
    wire new_AGEMA_signal_15424 ;
    wire new_AGEMA_signal_15425 ;
    wire new_AGEMA_signal_15426 ;
    wire new_AGEMA_signal_15427 ;
    wire new_AGEMA_signal_15428 ;
    wire new_AGEMA_signal_15429 ;
    wire new_AGEMA_signal_15430 ;
    wire new_AGEMA_signal_15431 ;
    wire new_AGEMA_signal_15432 ;
    wire new_AGEMA_signal_15433 ;
    wire new_AGEMA_signal_15434 ;
    wire new_AGEMA_signal_15435 ;
    wire new_AGEMA_signal_15436 ;
    wire new_AGEMA_signal_15437 ;
    wire new_AGEMA_signal_15438 ;
    wire new_AGEMA_signal_15439 ;
    wire new_AGEMA_signal_15440 ;
    wire new_AGEMA_signal_15441 ;
    wire new_AGEMA_signal_15442 ;
    wire new_AGEMA_signal_15443 ;
    wire new_AGEMA_signal_15444 ;
    wire new_AGEMA_signal_15445 ;
    wire new_AGEMA_signal_15446 ;
    wire new_AGEMA_signal_15447 ;
    wire new_AGEMA_signal_15448 ;
    wire new_AGEMA_signal_15449 ;
    wire new_AGEMA_signal_15450 ;
    wire new_AGEMA_signal_15451 ;
    wire new_AGEMA_signal_15452 ;
    wire new_AGEMA_signal_15453 ;
    wire new_AGEMA_signal_15454 ;
    wire new_AGEMA_signal_15455 ;
    wire new_AGEMA_signal_15456 ;
    wire new_AGEMA_signal_15457 ;
    wire new_AGEMA_signal_15458 ;
    wire new_AGEMA_signal_15459 ;
    wire new_AGEMA_signal_15460 ;
    wire new_AGEMA_signal_15461 ;
    wire new_AGEMA_signal_15462 ;
    wire new_AGEMA_signal_15463 ;
    wire new_AGEMA_signal_15464 ;
    wire new_AGEMA_signal_15465 ;
    wire new_AGEMA_signal_15466 ;
    wire new_AGEMA_signal_15467 ;
    wire new_AGEMA_signal_15468 ;
    wire new_AGEMA_signal_15469 ;
    wire new_AGEMA_signal_15470 ;
    wire new_AGEMA_signal_15471 ;
    wire new_AGEMA_signal_15472 ;
    wire new_AGEMA_signal_15473 ;
    wire new_AGEMA_signal_15474 ;
    wire new_AGEMA_signal_15475 ;
    wire new_AGEMA_signal_15476 ;
    wire new_AGEMA_signal_15477 ;
    wire new_AGEMA_signal_15478 ;
    wire new_AGEMA_signal_15479 ;
    wire new_AGEMA_signal_15480 ;
    wire new_AGEMA_signal_15481 ;
    wire new_AGEMA_signal_15482 ;
    wire new_AGEMA_signal_15483 ;
    wire new_AGEMA_signal_15484 ;
    wire new_AGEMA_signal_15485 ;
    wire new_AGEMA_signal_15486 ;
    wire new_AGEMA_signal_15487 ;
    wire new_AGEMA_signal_15488 ;
    wire new_AGEMA_signal_15489 ;
    wire new_AGEMA_signal_15490 ;
    wire new_AGEMA_signal_15491 ;
    wire new_AGEMA_signal_15492 ;
    wire new_AGEMA_signal_15493 ;
    wire new_AGEMA_signal_15494 ;
    wire new_AGEMA_signal_15495 ;
    wire new_AGEMA_signal_15496 ;
    wire new_AGEMA_signal_15497 ;
    wire new_AGEMA_signal_15498 ;
    wire new_AGEMA_signal_15499 ;
    wire new_AGEMA_signal_15500 ;
    wire new_AGEMA_signal_15501 ;
    wire new_AGEMA_signal_15502 ;
    wire new_AGEMA_signal_15503 ;
    wire new_AGEMA_signal_15504 ;
    wire new_AGEMA_signal_15505 ;
    wire new_AGEMA_signal_15506 ;
    wire new_AGEMA_signal_15507 ;
    wire new_AGEMA_signal_15508 ;
    wire new_AGEMA_signal_15509 ;
    wire new_AGEMA_signal_15510 ;
    wire new_AGEMA_signal_15511 ;
    wire new_AGEMA_signal_15512 ;
    wire new_AGEMA_signal_15513 ;
    wire new_AGEMA_signal_15514 ;
    wire new_AGEMA_signal_15515 ;
    wire new_AGEMA_signal_15516 ;
    wire new_AGEMA_signal_15517 ;
    wire new_AGEMA_signal_15518 ;
    wire new_AGEMA_signal_15519 ;
    wire new_AGEMA_signal_15520 ;
    wire new_AGEMA_signal_15521 ;
    wire new_AGEMA_signal_15522 ;
    wire new_AGEMA_signal_15523 ;
    wire new_AGEMA_signal_15524 ;
    wire new_AGEMA_signal_15525 ;
    wire new_AGEMA_signal_15526 ;
    wire new_AGEMA_signal_15527 ;
    wire new_AGEMA_signal_15528 ;
    wire new_AGEMA_signal_15529 ;
    wire new_AGEMA_signal_15530 ;
    wire new_AGEMA_signal_15531 ;
    wire new_AGEMA_signal_15532 ;
    wire new_AGEMA_signal_15533 ;
    wire new_AGEMA_signal_15534 ;
    wire new_AGEMA_signal_15535 ;
    wire new_AGEMA_signal_15536 ;
    wire new_AGEMA_signal_15537 ;
    wire new_AGEMA_signal_15538 ;
    wire new_AGEMA_signal_15539 ;
    wire new_AGEMA_signal_15540 ;
    wire new_AGEMA_signal_15541 ;
    wire new_AGEMA_signal_15542 ;
    wire new_AGEMA_signal_15543 ;
    wire new_AGEMA_signal_15544 ;
    wire new_AGEMA_signal_15545 ;
    wire new_AGEMA_signal_15546 ;
    wire new_AGEMA_signal_15547 ;
    wire new_AGEMA_signal_15548 ;
    wire new_AGEMA_signal_15549 ;
    wire new_AGEMA_signal_15550 ;
    wire new_AGEMA_signal_15551 ;
    wire new_AGEMA_signal_15552 ;
    wire new_AGEMA_signal_15553 ;
    wire new_AGEMA_signal_15554 ;
    wire new_AGEMA_signal_15555 ;
    wire new_AGEMA_signal_15556 ;
    wire new_AGEMA_signal_15557 ;
    wire new_AGEMA_signal_15558 ;
    wire new_AGEMA_signal_15559 ;
    wire new_AGEMA_signal_15560 ;
    wire new_AGEMA_signal_15561 ;
    wire new_AGEMA_signal_15562 ;
    wire new_AGEMA_signal_15563 ;
    wire new_AGEMA_signal_15564 ;
    wire new_AGEMA_signal_15565 ;
    wire new_AGEMA_signal_15566 ;
    wire new_AGEMA_signal_15567 ;
    wire new_AGEMA_signal_15568 ;
    wire new_AGEMA_signal_15569 ;
    wire new_AGEMA_signal_15570 ;
    wire new_AGEMA_signal_15571 ;
    wire new_AGEMA_signal_15572 ;
    wire new_AGEMA_signal_15573 ;
    wire new_AGEMA_signal_15574 ;
    wire new_AGEMA_signal_15575 ;
    wire new_AGEMA_signal_15576 ;
    wire new_AGEMA_signal_15577 ;
    wire new_AGEMA_signal_15578 ;
    wire new_AGEMA_signal_15579 ;
    wire new_AGEMA_signal_15580 ;
    wire new_AGEMA_signal_15581 ;
    wire new_AGEMA_signal_15582 ;
    wire new_AGEMA_signal_15583 ;
    wire new_AGEMA_signal_15584 ;
    wire new_AGEMA_signal_15585 ;
    wire new_AGEMA_signal_15586 ;
    wire new_AGEMA_signal_15587 ;
    wire new_AGEMA_signal_15588 ;
    wire new_AGEMA_signal_15589 ;
    wire new_AGEMA_signal_15590 ;
    wire new_AGEMA_signal_15591 ;
    wire new_AGEMA_signal_15592 ;
    wire new_AGEMA_signal_15593 ;
    wire new_AGEMA_signal_15594 ;
    wire new_AGEMA_signal_15595 ;
    wire new_AGEMA_signal_15596 ;
    wire new_AGEMA_signal_15597 ;
    wire new_AGEMA_signal_15598 ;
    wire new_AGEMA_signal_15599 ;
    wire new_AGEMA_signal_15600 ;
    wire new_AGEMA_signal_15601 ;
    wire new_AGEMA_signal_15602 ;
    wire new_AGEMA_signal_15603 ;
    wire new_AGEMA_signal_15604 ;
    wire new_AGEMA_signal_15605 ;
    wire new_AGEMA_signal_15606 ;
    wire new_AGEMA_signal_15607 ;
    wire new_AGEMA_signal_15608 ;
    wire new_AGEMA_signal_15609 ;
    wire new_AGEMA_signal_15610 ;
    wire new_AGEMA_signal_15611 ;
    wire new_AGEMA_signal_15612 ;
    wire new_AGEMA_signal_15613 ;
    wire new_AGEMA_signal_15614 ;
    wire new_AGEMA_signal_15615 ;
    wire new_AGEMA_signal_15616 ;
    wire new_AGEMA_signal_15617 ;
    wire new_AGEMA_signal_15618 ;
    wire new_AGEMA_signal_15619 ;
    wire new_AGEMA_signal_15620 ;
    wire new_AGEMA_signal_15621 ;
    wire new_AGEMA_signal_15622 ;
    wire new_AGEMA_signal_15623 ;
    wire new_AGEMA_signal_15624 ;
    wire new_AGEMA_signal_15625 ;
    wire new_AGEMA_signal_15626 ;
    wire new_AGEMA_signal_15627 ;
    wire new_AGEMA_signal_15628 ;
    wire new_AGEMA_signal_15629 ;
    wire new_AGEMA_signal_15630 ;
    wire new_AGEMA_signal_15631 ;
    wire new_AGEMA_signal_15632 ;
    wire new_AGEMA_signal_15633 ;
    wire new_AGEMA_signal_15634 ;
    wire new_AGEMA_signal_15635 ;
    wire new_AGEMA_signal_15636 ;
    wire new_AGEMA_signal_15637 ;
    wire new_AGEMA_signal_15638 ;
    wire new_AGEMA_signal_15639 ;
    wire new_AGEMA_signal_15640 ;
    wire new_AGEMA_signal_15641 ;
    wire new_AGEMA_signal_15642 ;
    wire new_AGEMA_signal_15643 ;
    wire new_AGEMA_signal_15644 ;
    wire new_AGEMA_signal_15645 ;
    wire new_AGEMA_signal_15646 ;
    wire new_AGEMA_signal_15647 ;
    wire new_AGEMA_signal_15648 ;
    wire new_AGEMA_signal_15649 ;
    wire new_AGEMA_signal_15650 ;
    wire new_AGEMA_signal_15651 ;
    wire new_AGEMA_signal_15652 ;
    wire new_AGEMA_signal_15653 ;
    wire new_AGEMA_signal_15654 ;
    wire new_AGEMA_signal_15655 ;
    wire new_AGEMA_signal_15656 ;
    wire new_AGEMA_signal_15657 ;
    wire new_AGEMA_signal_15658 ;
    wire new_AGEMA_signal_15659 ;
    wire new_AGEMA_signal_15660 ;
    wire new_AGEMA_signal_15661 ;
    wire new_AGEMA_signal_15662 ;
    wire new_AGEMA_signal_15663 ;
    wire new_AGEMA_signal_15664 ;
    wire new_AGEMA_signal_15665 ;
    wire new_AGEMA_signal_15666 ;
    wire new_AGEMA_signal_15667 ;
    wire new_AGEMA_signal_15668 ;
    wire new_AGEMA_signal_15669 ;
    wire new_AGEMA_signal_15670 ;
    wire new_AGEMA_signal_15671 ;
    wire new_AGEMA_signal_15672 ;
    wire new_AGEMA_signal_15673 ;
    wire new_AGEMA_signal_15674 ;
    wire new_AGEMA_signal_15675 ;
    wire new_AGEMA_signal_15676 ;
    wire new_AGEMA_signal_15677 ;
    wire new_AGEMA_signal_15678 ;
    wire new_AGEMA_signal_15679 ;
    wire new_AGEMA_signal_15680 ;
    wire new_AGEMA_signal_15681 ;
    wire new_AGEMA_signal_15682 ;
    wire new_AGEMA_signal_15683 ;
    wire new_AGEMA_signal_15684 ;
    wire new_AGEMA_signal_15685 ;
    wire new_AGEMA_signal_15686 ;
    wire new_AGEMA_signal_15687 ;
    wire new_AGEMA_signal_15688 ;
    wire new_AGEMA_signal_15689 ;
    wire new_AGEMA_signal_15690 ;
    wire new_AGEMA_signal_15691 ;
    wire new_AGEMA_signal_15692 ;
    wire new_AGEMA_signal_15693 ;
    wire new_AGEMA_signal_15694 ;
    wire new_AGEMA_signal_15695 ;
    wire new_AGEMA_signal_15696 ;
    wire new_AGEMA_signal_15697 ;
    wire new_AGEMA_signal_15698 ;
    wire new_AGEMA_signal_15699 ;
    wire new_AGEMA_signal_15700 ;
    wire new_AGEMA_signal_15701 ;
    wire new_AGEMA_signal_15702 ;
    wire new_AGEMA_signal_15703 ;
    wire new_AGEMA_signal_15704 ;
    wire new_AGEMA_signal_15705 ;
    wire new_AGEMA_signal_15706 ;
    wire new_AGEMA_signal_15707 ;
    wire new_AGEMA_signal_15708 ;
    wire new_AGEMA_signal_15709 ;
    wire new_AGEMA_signal_15710 ;
    wire new_AGEMA_signal_15711 ;
    wire new_AGEMA_signal_15712 ;
    wire new_AGEMA_signal_15713 ;
    wire new_AGEMA_signal_15714 ;
    wire new_AGEMA_signal_15715 ;
    wire new_AGEMA_signal_15716 ;
    wire new_AGEMA_signal_15717 ;
    wire new_AGEMA_signal_15718 ;
    wire new_AGEMA_signal_15719 ;
    wire new_AGEMA_signal_15720 ;
    wire new_AGEMA_signal_15721 ;
    wire new_AGEMA_signal_15722 ;
    wire new_AGEMA_signal_15723 ;
    wire new_AGEMA_signal_15724 ;
    wire new_AGEMA_signal_15725 ;
    wire new_AGEMA_signal_15726 ;
    wire new_AGEMA_signal_15727 ;
    wire new_AGEMA_signal_15728 ;
    wire new_AGEMA_signal_15729 ;
    wire new_AGEMA_signal_15730 ;
    wire new_AGEMA_signal_15731 ;
    wire new_AGEMA_signal_15732 ;
    wire new_AGEMA_signal_15733 ;
    wire new_AGEMA_signal_15734 ;
    wire new_AGEMA_signal_15735 ;
    wire new_AGEMA_signal_15736 ;
    wire new_AGEMA_signal_15737 ;
    wire new_AGEMA_signal_15738 ;
    wire new_AGEMA_signal_15739 ;
    wire new_AGEMA_signal_15740 ;
    wire new_AGEMA_signal_15741 ;
    wire new_AGEMA_signal_15742 ;
    wire new_AGEMA_signal_15743 ;
    wire new_AGEMA_signal_15744 ;
    wire new_AGEMA_signal_15745 ;
    wire new_AGEMA_signal_15746 ;
    wire new_AGEMA_signal_15747 ;
    wire new_AGEMA_signal_15748 ;
    wire new_AGEMA_signal_15749 ;
    wire new_AGEMA_signal_15750 ;
    wire new_AGEMA_signal_15751 ;
    wire new_AGEMA_signal_15752 ;
    wire new_AGEMA_signal_15753 ;
    wire new_AGEMA_signal_15754 ;
    wire new_AGEMA_signal_15755 ;
    wire new_AGEMA_signal_15756 ;
    wire new_AGEMA_signal_15757 ;
    wire new_AGEMA_signal_15758 ;
    wire new_AGEMA_signal_15759 ;
    wire new_AGEMA_signal_15760 ;
    wire new_AGEMA_signal_15761 ;
    wire new_AGEMA_signal_15762 ;
    wire new_AGEMA_signal_15763 ;
    wire new_AGEMA_signal_15764 ;
    wire new_AGEMA_signal_15765 ;
    wire new_AGEMA_signal_15766 ;
    wire new_AGEMA_signal_15767 ;
    wire new_AGEMA_signal_15768 ;
    wire new_AGEMA_signal_15769 ;
    wire new_AGEMA_signal_15770 ;
    wire new_AGEMA_signal_15771 ;
    wire new_AGEMA_signal_15772 ;
    wire new_AGEMA_signal_15773 ;
    wire new_AGEMA_signal_15774 ;
    wire new_AGEMA_signal_15775 ;
    wire new_AGEMA_signal_15776 ;
    wire new_AGEMA_signal_15777 ;
    wire new_AGEMA_signal_15778 ;
    wire new_AGEMA_signal_15779 ;
    wire new_AGEMA_signal_15780 ;
    wire new_AGEMA_signal_15781 ;
    wire new_AGEMA_signal_15782 ;
    wire new_AGEMA_signal_15783 ;
    wire new_AGEMA_signal_15784 ;
    wire new_AGEMA_signal_15785 ;
    wire new_AGEMA_signal_15786 ;
    wire new_AGEMA_signal_15787 ;
    wire new_AGEMA_signal_15788 ;
    wire new_AGEMA_signal_15789 ;
    wire new_AGEMA_signal_15790 ;
    wire new_AGEMA_signal_15791 ;
    wire new_AGEMA_signal_15792 ;
    wire new_AGEMA_signal_15793 ;
    wire new_AGEMA_signal_15794 ;
    wire new_AGEMA_signal_15795 ;
    wire new_AGEMA_signal_15796 ;
    wire new_AGEMA_signal_15797 ;
    wire new_AGEMA_signal_15798 ;
    wire new_AGEMA_signal_15799 ;
    wire new_AGEMA_signal_15800 ;
    wire new_AGEMA_signal_15801 ;
    wire new_AGEMA_signal_15802 ;
    wire new_AGEMA_signal_15803 ;
    wire new_AGEMA_signal_15804 ;
    wire new_AGEMA_signal_15805 ;
    wire new_AGEMA_signal_15806 ;
    wire new_AGEMA_signal_15807 ;
    wire new_AGEMA_signal_15808 ;
    wire new_AGEMA_signal_15809 ;
    wire new_AGEMA_signal_15810 ;
    wire new_AGEMA_signal_15811 ;
    wire new_AGEMA_signal_15812 ;
    wire new_AGEMA_signal_15813 ;
    wire new_AGEMA_signal_15814 ;
    wire new_AGEMA_signal_15815 ;
    wire new_AGEMA_signal_15816 ;
    wire new_AGEMA_signal_15817 ;
    wire new_AGEMA_signal_15818 ;
    wire new_AGEMA_signal_15819 ;
    wire new_AGEMA_signal_15820 ;
    wire new_AGEMA_signal_15821 ;
    wire new_AGEMA_signal_15822 ;
    wire new_AGEMA_signal_15823 ;
    wire new_AGEMA_signal_15824 ;
    wire new_AGEMA_signal_15825 ;
    wire new_AGEMA_signal_15826 ;
    wire new_AGEMA_signal_15827 ;
    wire new_AGEMA_signal_15828 ;
    wire new_AGEMA_signal_15829 ;
    wire new_AGEMA_signal_15830 ;
    wire new_AGEMA_signal_15831 ;
    wire new_AGEMA_signal_15832 ;
    wire new_AGEMA_signal_15833 ;
    wire new_AGEMA_signal_15834 ;
    wire new_AGEMA_signal_15835 ;
    wire new_AGEMA_signal_15836 ;
    wire new_AGEMA_signal_15837 ;
    wire new_AGEMA_signal_15838 ;
    wire new_AGEMA_signal_15839 ;
    wire new_AGEMA_signal_15840 ;
    wire new_AGEMA_signal_15841 ;
    wire new_AGEMA_signal_15842 ;
    wire new_AGEMA_signal_15843 ;
    wire new_AGEMA_signal_15844 ;
    wire new_AGEMA_signal_15845 ;
    wire new_AGEMA_signal_15846 ;
    wire new_AGEMA_signal_15847 ;
    wire new_AGEMA_signal_15848 ;
    wire new_AGEMA_signal_15849 ;
    wire new_AGEMA_signal_15850 ;
    wire new_AGEMA_signal_15851 ;
    wire new_AGEMA_signal_15852 ;
    wire new_AGEMA_signal_15853 ;
    wire new_AGEMA_signal_15854 ;
    wire new_AGEMA_signal_15855 ;
    wire new_AGEMA_signal_15856 ;
    wire new_AGEMA_signal_15857 ;
    wire new_AGEMA_signal_15858 ;
    wire new_AGEMA_signal_15859 ;
    wire new_AGEMA_signal_15860 ;
    wire new_AGEMA_signal_15861 ;
    wire new_AGEMA_signal_15862 ;
    wire new_AGEMA_signal_15863 ;
    wire new_AGEMA_signal_15864 ;
    wire new_AGEMA_signal_15865 ;
    wire new_AGEMA_signal_15866 ;
    wire new_AGEMA_signal_15867 ;
    wire new_AGEMA_signal_15868 ;
    wire new_AGEMA_signal_15869 ;
    wire new_AGEMA_signal_15870 ;
    wire new_AGEMA_signal_15871 ;
    wire new_AGEMA_signal_15872 ;
    wire new_AGEMA_signal_15873 ;
    wire new_AGEMA_signal_15874 ;
    wire new_AGEMA_signal_15875 ;
    wire new_AGEMA_signal_15876 ;
    wire new_AGEMA_signal_15877 ;
    wire new_AGEMA_signal_15878 ;
    wire new_AGEMA_signal_15879 ;
    wire new_AGEMA_signal_15880 ;
    wire new_AGEMA_signal_15881 ;
    wire new_AGEMA_signal_15882 ;
    wire new_AGEMA_signal_15883 ;
    wire new_AGEMA_signal_15884 ;
    wire new_AGEMA_signal_15885 ;
    wire new_AGEMA_signal_15886 ;
    wire new_AGEMA_signal_15887 ;
    wire new_AGEMA_signal_15888 ;
    wire new_AGEMA_signal_15889 ;
    wire new_AGEMA_signal_15890 ;
    wire new_AGEMA_signal_15891 ;
    wire new_AGEMA_signal_15892 ;
    wire new_AGEMA_signal_15893 ;
    wire new_AGEMA_signal_15894 ;
    wire new_AGEMA_signal_15895 ;
    wire new_AGEMA_signal_15896 ;
    wire new_AGEMA_signal_15897 ;
    wire new_AGEMA_signal_15898 ;
    wire new_AGEMA_signal_15899 ;
    wire new_AGEMA_signal_15900 ;
    wire new_AGEMA_signal_15901 ;
    wire new_AGEMA_signal_15902 ;
    wire new_AGEMA_signal_15903 ;
    wire new_AGEMA_signal_15904 ;
    wire new_AGEMA_signal_15905 ;
    wire new_AGEMA_signal_15906 ;
    wire new_AGEMA_signal_15907 ;
    wire new_AGEMA_signal_15908 ;
    wire new_AGEMA_signal_15909 ;
    wire new_AGEMA_signal_15910 ;
    wire new_AGEMA_signal_15911 ;
    wire new_AGEMA_signal_15912 ;
    wire new_AGEMA_signal_15913 ;
    wire new_AGEMA_signal_15914 ;
    wire new_AGEMA_signal_15915 ;
    wire new_AGEMA_signal_15916 ;
    wire new_AGEMA_signal_15917 ;
    wire new_AGEMA_signal_15918 ;
    wire new_AGEMA_signal_15919 ;
    wire new_AGEMA_signal_15920 ;
    wire new_AGEMA_signal_15921 ;
    wire new_AGEMA_signal_15922 ;
    wire new_AGEMA_signal_15923 ;
    wire new_AGEMA_signal_15924 ;
    wire new_AGEMA_signal_15925 ;
    wire new_AGEMA_signal_15926 ;
    wire new_AGEMA_signal_15927 ;
    wire new_AGEMA_signal_15928 ;
    wire new_AGEMA_signal_15929 ;
    wire new_AGEMA_signal_15930 ;
    wire new_AGEMA_signal_15931 ;
    wire new_AGEMA_signal_15932 ;
    wire new_AGEMA_signal_15933 ;
    wire new_AGEMA_signal_15934 ;
    wire new_AGEMA_signal_15935 ;
    wire new_AGEMA_signal_15936 ;
    wire new_AGEMA_signal_15937 ;
    wire new_AGEMA_signal_15938 ;
    wire new_AGEMA_signal_15939 ;
    wire new_AGEMA_signal_15940 ;
    wire new_AGEMA_signal_15941 ;
    wire new_AGEMA_signal_15942 ;
    wire new_AGEMA_signal_15943 ;
    wire new_AGEMA_signal_15944 ;
    wire new_AGEMA_signal_15945 ;
    wire new_AGEMA_signal_15946 ;
    wire new_AGEMA_signal_15947 ;
    wire new_AGEMA_signal_15948 ;
    wire new_AGEMA_signal_15949 ;
    wire new_AGEMA_signal_15950 ;
    wire new_AGEMA_signal_15951 ;
    wire new_AGEMA_signal_15952 ;
    wire new_AGEMA_signal_15953 ;
    wire new_AGEMA_signal_15954 ;
    wire new_AGEMA_signal_15955 ;
    wire new_AGEMA_signal_15956 ;
    wire new_AGEMA_signal_15957 ;
    wire new_AGEMA_signal_15958 ;
    wire new_AGEMA_signal_15959 ;
    wire new_AGEMA_signal_15960 ;
    wire new_AGEMA_signal_15961 ;
    wire new_AGEMA_signal_15962 ;
    wire new_AGEMA_signal_15963 ;
    wire new_AGEMA_signal_15964 ;
    wire new_AGEMA_signal_15965 ;
    wire new_AGEMA_signal_15966 ;
    wire new_AGEMA_signal_15967 ;
    wire new_AGEMA_signal_15968 ;
    wire new_AGEMA_signal_15969 ;
    wire new_AGEMA_signal_15970 ;
    wire new_AGEMA_signal_15971 ;
    wire new_AGEMA_signal_15972 ;
    wire new_AGEMA_signal_15973 ;
    wire new_AGEMA_signal_15974 ;
    wire new_AGEMA_signal_15975 ;
    wire new_AGEMA_signal_15976 ;
    wire new_AGEMA_signal_15977 ;
    wire new_AGEMA_signal_15978 ;
    wire new_AGEMA_signal_15979 ;
    wire new_AGEMA_signal_15980 ;
    wire new_AGEMA_signal_15981 ;
    wire new_AGEMA_signal_15982 ;
    wire new_AGEMA_signal_15983 ;
    wire new_AGEMA_signal_15984 ;
    wire new_AGEMA_signal_15985 ;
    wire new_AGEMA_signal_15986 ;
    wire new_AGEMA_signal_15987 ;
    wire new_AGEMA_signal_15988 ;
    wire new_AGEMA_signal_15989 ;
    wire new_AGEMA_signal_15990 ;
    wire new_AGEMA_signal_15991 ;
    wire new_AGEMA_signal_15992 ;
    wire new_AGEMA_signal_15993 ;
    wire new_AGEMA_signal_15994 ;
    wire new_AGEMA_signal_15995 ;
    wire new_AGEMA_signal_15996 ;
    wire new_AGEMA_signal_15997 ;
    wire new_AGEMA_signal_15998 ;
    wire new_AGEMA_signal_15999 ;
    wire new_AGEMA_signal_16000 ;
    wire new_AGEMA_signal_16001 ;
    wire new_AGEMA_signal_16002 ;
    wire new_AGEMA_signal_16003 ;
    wire new_AGEMA_signal_16004 ;
    wire new_AGEMA_signal_16005 ;
    wire new_AGEMA_signal_16006 ;
    wire new_AGEMA_signal_16007 ;
    wire new_AGEMA_signal_16008 ;
    wire new_AGEMA_signal_16009 ;
    wire new_AGEMA_signal_16010 ;
    wire new_AGEMA_signal_16011 ;
    wire new_AGEMA_signal_16012 ;
    wire new_AGEMA_signal_16013 ;
    wire new_AGEMA_signal_16014 ;
    wire new_AGEMA_signal_16015 ;
    wire new_AGEMA_signal_16016 ;
    wire new_AGEMA_signal_16017 ;
    wire new_AGEMA_signal_16018 ;
    wire new_AGEMA_signal_16019 ;
    wire new_AGEMA_signal_16020 ;
    wire new_AGEMA_signal_16021 ;
    wire new_AGEMA_signal_16022 ;
    wire new_AGEMA_signal_16023 ;
    wire new_AGEMA_signal_16024 ;
    wire new_AGEMA_signal_16025 ;
    wire new_AGEMA_signal_16026 ;
    wire new_AGEMA_signal_16027 ;
    wire new_AGEMA_signal_16028 ;
    wire new_AGEMA_signal_16029 ;
    wire new_AGEMA_signal_16030 ;
    wire new_AGEMA_signal_16031 ;
    wire new_AGEMA_signal_16032 ;
    wire new_AGEMA_signal_16033 ;
    wire new_AGEMA_signal_16034 ;
    wire new_AGEMA_signal_16035 ;
    wire new_AGEMA_signal_16036 ;
    wire new_AGEMA_signal_16037 ;
    wire new_AGEMA_signal_16038 ;
    wire new_AGEMA_signal_16039 ;
    wire new_AGEMA_signal_16040 ;
    wire new_AGEMA_signal_16041 ;
    wire new_AGEMA_signal_16042 ;
    wire new_AGEMA_signal_16043 ;
    wire new_AGEMA_signal_16044 ;
    wire new_AGEMA_signal_16045 ;
    wire new_AGEMA_signal_16046 ;
    wire new_AGEMA_signal_16047 ;
    wire new_AGEMA_signal_16048 ;
    wire new_AGEMA_signal_16049 ;
    wire new_AGEMA_signal_16050 ;
    wire new_AGEMA_signal_16051 ;
    wire new_AGEMA_signal_16052 ;
    wire new_AGEMA_signal_16053 ;
    wire new_AGEMA_signal_16054 ;
    wire new_AGEMA_signal_16055 ;
    wire new_AGEMA_signal_16056 ;
    wire new_AGEMA_signal_16057 ;
    wire new_AGEMA_signal_16058 ;
    wire new_AGEMA_signal_16059 ;
    wire new_AGEMA_signal_16060 ;
    wire new_AGEMA_signal_16061 ;
    wire new_AGEMA_signal_16062 ;
    wire new_AGEMA_signal_16063 ;
    wire new_AGEMA_signal_16064 ;
    wire new_AGEMA_signal_16065 ;
    wire new_AGEMA_signal_16066 ;
    wire new_AGEMA_signal_16067 ;
    wire new_AGEMA_signal_16068 ;
    wire new_AGEMA_signal_16069 ;
    wire new_AGEMA_signal_16070 ;
    wire new_AGEMA_signal_16071 ;
    wire new_AGEMA_signal_16072 ;
    wire new_AGEMA_signal_16073 ;
    wire new_AGEMA_signal_16074 ;
    wire new_AGEMA_signal_16075 ;
    wire new_AGEMA_signal_16076 ;
    wire new_AGEMA_signal_16077 ;
    wire new_AGEMA_signal_16078 ;
    wire new_AGEMA_signal_16079 ;
    wire new_AGEMA_signal_16080 ;
    wire new_AGEMA_signal_16081 ;
    wire new_AGEMA_signal_16082 ;
    wire new_AGEMA_signal_16083 ;
    wire new_AGEMA_signal_16084 ;
    wire new_AGEMA_signal_16085 ;
    wire new_AGEMA_signal_16086 ;
    wire new_AGEMA_signal_16087 ;
    wire new_AGEMA_signal_16088 ;
    wire new_AGEMA_signal_16089 ;
    wire new_AGEMA_signal_16090 ;
    wire new_AGEMA_signal_16091 ;
    wire new_AGEMA_signal_16092 ;
    wire new_AGEMA_signal_16093 ;
    wire new_AGEMA_signal_16094 ;
    wire new_AGEMA_signal_16095 ;
    wire new_AGEMA_signal_16096 ;
    wire new_AGEMA_signal_16097 ;
    wire new_AGEMA_signal_16098 ;
    wire new_AGEMA_signal_16099 ;
    wire new_AGEMA_signal_16100 ;
    wire new_AGEMA_signal_16101 ;
    wire new_AGEMA_signal_16102 ;
    wire new_AGEMA_signal_16103 ;
    wire new_AGEMA_signal_16104 ;
    wire new_AGEMA_signal_16105 ;
    wire new_AGEMA_signal_16106 ;
    wire new_AGEMA_signal_16107 ;
    wire new_AGEMA_signal_16108 ;
    wire new_AGEMA_signal_16109 ;
    wire new_AGEMA_signal_16110 ;
    wire new_AGEMA_signal_16111 ;
    wire new_AGEMA_signal_16112 ;
    wire new_AGEMA_signal_16113 ;
    wire new_AGEMA_signal_16114 ;
    wire new_AGEMA_signal_16115 ;
    wire new_AGEMA_signal_16116 ;
    wire new_AGEMA_signal_16117 ;
    wire new_AGEMA_signal_16118 ;
    wire new_AGEMA_signal_16119 ;
    wire new_AGEMA_signal_16120 ;
    wire new_AGEMA_signal_16121 ;
    wire new_AGEMA_signal_16122 ;
    wire new_AGEMA_signal_16123 ;
    wire new_AGEMA_signal_16124 ;
    wire new_AGEMA_signal_16125 ;
    wire new_AGEMA_signal_16126 ;
    wire new_AGEMA_signal_16127 ;
    wire new_AGEMA_signal_16128 ;
    wire new_AGEMA_signal_16129 ;
    wire new_AGEMA_signal_16130 ;
    wire new_AGEMA_signal_16131 ;
    wire new_AGEMA_signal_16132 ;
    wire new_AGEMA_signal_16133 ;
    wire new_AGEMA_signal_16134 ;
    wire new_AGEMA_signal_16135 ;
    wire new_AGEMA_signal_16136 ;
    wire new_AGEMA_signal_16137 ;
    wire new_AGEMA_signal_16138 ;
    wire new_AGEMA_signal_16139 ;
    wire new_AGEMA_signal_16140 ;
    wire new_AGEMA_signal_16141 ;
    wire new_AGEMA_signal_16142 ;
    wire new_AGEMA_signal_16143 ;
    wire new_AGEMA_signal_16144 ;
    wire new_AGEMA_signal_16145 ;
    wire new_AGEMA_signal_16146 ;
    wire new_AGEMA_signal_16147 ;
    wire new_AGEMA_signal_16148 ;
    wire new_AGEMA_signal_16149 ;
    wire new_AGEMA_signal_16150 ;
    wire new_AGEMA_signal_16151 ;
    wire new_AGEMA_signal_16152 ;
    wire new_AGEMA_signal_16153 ;
    wire new_AGEMA_signal_16154 ;
    wire new_AGEMA_signal_16155 ;
    wire new_AGEMA_signal_16156 ;
    wire new_AGEMA_signal_16157 ;
    wire new_AGEMA_signal_16158 ;
    wire new_AGEMA_signal_16159 ;
    wire new_AGEMA_signal_16160 ;
    wire new_AGEMA_signal_16161 ;
    wire new_AGEMA_signal_16162 ;
    wire new_AGEMA_signal_16163 ;
    wire new_AGEMA_signal_16164 ;
    wire new_AGEMA_signal_16165 ;
    wire new_AGEMA_signal_16166 ;
    wire new_AGEMA_signal_16167 ;
    wire new_AGEMA_signal_16168 ;
    wire new_AGEMA_signal_16169 ;
    wire new_AGEMA_signal_16170 ;
    wire new_AGEMA_signal_16171 ;
    wire new_AGEMA_signal_16172 ;
    wire new_AGEMA_signal_16173 ;
    wire new_AGEMA_signal_16174 ;
    wire new_AGEMA_signal_16175 ;
    wire new_AGEMA_signal_16176 ;
    wire new_AGEMA_signal_16177 ;
    wire new_AGEMA_signal_16178 ;
    wire new_AGEMA_signal_16179 ;
    wire new_AGEMA_signal_16180 ;
    wire new_AGEMA_signal_16181 ;
    wire new_AGEMA_signal_16182 ;
    wire new_AGEMA_signal_16183 ;
    wire new_AGEMA_signal_16184 ;
    wire new_AGEMA_signal_16185 ;
    wire new_AGEMA_signal_16186 ;
    wire new_AGEMA_signal_16187 ;
    wire new_AGEMA_signal_16188 ;
    wire new_AGEMA_signal_16189 ;
    wire new_AGEMA_signal_16190 ;
    wire new_AGEMA_signal_16191 ;
    wire new_AGEMA_signal_16192 ;
    wire new_AGEMA_signal_16193 ;
    wire new_AGEMA_signal_16194 ;
    wire new_AGEMA_signal_16195 ;
    wire new_AGEMA_signal_16196 ;
    wire new_AGEMA_signal_16197 ;
    wire new_AGEMA_signal_16198 ;
    wire new_AGEMA_signal_16199 ;
    wire new_AGEMA_signal_16200 ;
    wire new_AGEMA_signal_16201 ;
    wire new_AGEMA_signal_16202 ;
    wire new_AGEMA_signal_16203 ;
    wire new_AGEMA_signal_16204 ;
    wire new_AGEMA_signal_16205 ;
    wire new_AGEMA_signal_16206 ;
    wire new_AGEMA_signal_16207 ;
    wire new_AGEMA_signal_16208 ;
    wire new_AGEMA_signal_16209 ;
    wire new_AGEMA_signal_16210 ;
    wire new_AGEMA_signal_16211 ;
    wire new_AGEMA_signal_16212 ;
    wire new_AGEMA_signal_16213 ;
    wire new_AGEMA_signal_16214 ;
    wire new_AGEMA_signal_16215 ;
    wire new_AGEMA_signal_16216 ;
    wire new_AGEMA_signal_16217 ;
    wire new_AGEMA_signal_16218 ;
    wire new_AGEMA_signal_16219 ;
    wire new_AGEMA_signal_16220 ;
    wire new_AGEMA_signal_16221 ;
    wire new_AGEMA_signal_16222 ;
    wire new_AGEMA_signal_16223 ;
    wire new_AGEMA_signal_16224 ;
    wire new_AGEMA_signal_16225 ;
    wire new_AGEMA_signal_16226 ;
    wire new_AGEMA_signal_16227 ;
    wire new_AGEMA_signal_16228 ;
    wire new_AGEMA_signal_16229 ;
    wire new_AGEMA_signal_16230 ;
    wire new_AGEMA_signal_16231 ;
    wire new_AGEMA_signal_16232 ;
    wire new_AGEMA_signal_16233 ;
    wire new_AGEMA_signal_16234 ;
    wire new_AGEMA_signal_16235 ;
    wire new_AGEMA_signal_16236 ;
    wire new_AGEMA_signal_16237 ;
    wire new_AGEMA_signal_16238 ;
    wire new_AGEMA_signal_16239 ;
    wire new_AGEMA_signal_16240 ;
    wire new_AGEMA_signal_16241 ;
    wire new_AGEMA_signal_16242 ;
    wire new_AGEMA_signal_16243 ;
    wire new_AGEMA_signal_16244 ;
    wire new_AGEMA_signal_16245 ;
    wire new_AGEMA_signal_16246 ;
    wire new_AGEMA_signal_16247 ;
    wire new_AGEMA_signal_16248 ;
    wire new_AGEMA_signal_16249 ;
    wire new_AGEMA_signal_16250 ;
    wire new_AGEMA_signal_16251 ;
    wire new_AGEMA_signal_16252 ;
    wire new_AGEMA_signal_16253 ;
    wire new_AGEMA_signal_16254 ;
    wire new_AGEMA_signal_16255 ;
    wire new_AGEMA_signal_16256 ;
    wire new_AGEMA_signal_16257 ;
    wire new_AGEMA_signal_16258 ;
    wire new_AGEMA_signal_16259 ;
    wire new_AGEMA_signal_16260 ;
    wire new_AGEMA_signal_16261 ;
    wire new_AGEMA_signal_16262 ;
    wire new_AGEMA_signal_16263 ;
    wire new_AGEMA_signal_16264 ;
    wire new_AGEMA_signal_16265 ;
    wire new_AGEMA_signal_16266 ;
    wire new_AGEMA_signal_16267 ;
    wire new_AGEMA_signal_16268 ;
    wire new_AGEMA_signal_16269 ;
    wire new_AGEMA_signal_16270 ;
    wire new_AGEMA_signal_16271 ;
    wire new_AGEMA_signal_16272 ;
    wire new_AGEMA_signal_16273 ;
    wire new_AGEMA_signal_16274 ;
    wire new_AGEMA_signal_16275 ;
    wire new_AGEMA_signal_16276 ;
    wire new_AGEMA_signal_16277 ;
    wire new_AGEMA_signal_16278 ;
    wire new_AGEMA_signal_16279 ;
    wire new_AGEMA_signal_16280 ;
    wire new_AGEMA_signal_16281 ;
    wire new_AGEMA_signal_16282 ;
    wire new_AGEMA_signal_16283 ;
    wire new_AGEMA_signal_16284 ;
    wire new_AGEMA_signal_16285 ;
    wire new_AGEMA_signal_16286 ;
    wire new_AGEMA_signal_16287 ;
    wire new_AGEMA_signal_16288 ;
    wire new_AGEMA_signal_16289 ;
    wire new_AGEMA_signal_16290 ;
    wire new_AGEMA_signal_16291 ;
    wire new_AGEMA_signal_16292 ;
    wire new_AGEMA_signal_16293 ;
    wire new_AGEMA_signal_16294 ;
    wire new_AGEMA_signal_16295 ;
    wire new_AGEMA_signal_16296 ;
    wire new_AGEMA_signal_16297 ;
    wire new_AGEMA_signal_16298 ;
    wire new_AGEMA_signal_16299 ;
    wire new_AGEMA_signal_16300 ;
    wire new_AGEMA_signal_16301 ;
    wire new_AGEMA_signal_16302 ;
    wire new_AGEMA_signal_16303 ;
    wire new_AGEMA_signal_16304 ;
    wire new_AGEMA_signal_16305 ;
    wire new_AGEMA_signal_16306 ;
    wire new_AGEMA_signal_16307 ;
    wire new_AGEMA_signal_16308 ;
    wire new_AGEMA_signal_16309 ;
    wire new_AGEMA_signal_16310 ;
    wire new_AGEMA_signal_16311 ;
    wire new_AGEMA_signal_16312 ;
    wire new_AGEMA_signal_16313 ;
    wire new_AGEMA_signal_16314 ;
    wire new_AGEMA_signal_16315 ;
    wire new_AGEMA_signal_16316 ;
    wire new_AGEMA_signal_16317 ;
    wire new_AGEMA_signal_16318 ;
    wire new_AGEMA_signal_16319 ;
    wire new_AGEMA_signal_16320 ;
    wire new_AGEMA_signal_16321 ;
    wire new_AGEMA_signal_16322 ;
    wire new_AGEMA_signal_16323 ;
    wire new_AGEMA_signal_16324 ;
    wire new_AGEMA_signal_16325 ;
    wire new_AGEMA_signal_16326 ;
    wire new_AGEMA_signal_16327 ;
    wire new_AGEMA_signal_16328 ;
    wire new_AGEMA_signal_16329 ;
    wire new_AGEMA_signal_16330 ;
    wire new_AGEMA_signal_16331 ;
    wire new_AGEMA_signal_16332 ;
    wire new_AGEMA_signal_16333 ;
    wire new_AGEMA_signal_16334 ;
    wire new_AGEMA_signal_16335 ;
    wire new_AGEMA_signal_16336 ;
    wire new_AGEMA_signal_16337 ;
    wire new_AGEMA_signal_16338 ;
    wire new_AGEMA_signal_16339 ;
    wire new_AGEMA_signal_16340 ;
    wire new_AGEMA_signal_16341 ;
    wire new_AGEMA_signal_16342 ;
    wire new_AGEMA_signal_16343 ;
    wire new_AGEMA_signal_16344 ;
    wire new_AGEMA_signal_16345 ;
    wire new_AGEMA_signal_16346 ;
    wire new_AGEMA_signal_16347 ;
    wire new_AGEMA_signal_16348 ;
    wire new_AGEMA_signal_16349 ;
    wire new_AGEMA_signal_16350 ;
    wire new_AGEMA_signal_16351 ;
    wire new_AGEMA_signal_16352 ;
    wire new_AGEMA_signal_16353 ;
    wire new_AGEMA_signal_16354 ;
    wire new_AGEMA_signal_16355 ;
    wire new_AGEMA_signal_16356 ;
    wire new_AGEMA_signal_16357 ;
    wire new_AGEMA_signal_16358 ;
    wire new_AGEMA_signal_16359 ;
    wire new_AGEMA_signal_16360 ;
    wire new_AGEMA_signal_16361 ;
    wire new_AGEMA_signal_16362 ;
    wire new_AGEMA_signal_16363 ;
    wire new_AGEMA_signal_16364 ;
    wire new_AGEMA_signal_16365 ;
    wire new_AGEMA_signal_16366 ;
    wire new_AGEMA_signal_16367 ;
    wire new_AGEMA_signal_16368 ;
    wire new_AGEMA_signal_16369 ;
    wire new_AGEMA_signal_16370 ;
    wire new_AGEMA_signal_16371 ;
    wire new_AGEMA_signal_16372 ;
    wire new_AGEMA_signal_16373 ;
    wire new_AGEMA_signal_16374 ;
    wire new_AGEMA_signal_16375 ;
    wire new_AGEMA_signal_16376 ;
    wire new_AGEMA_signal_16377 ;
    wire new_AGEMA_signal_16378 ;
    wire new_AGEMA_signal_16379 ;
    wire new_AGEMA_signal_16380 ;
    wire new_AGEMA_signal_16381 ;
    wire new_AGEMA_signal_16382 ;
    wire new_AGEMA_signal_16383 ;
    wire new_AGEMA_signal_16384 ;
    wire new_AGEMA_signal_16385 ;
    wire new_AGEMA_signal_16386 ;
    wire new_AGEMA_signal_16387 ;
    wire new_AGEMA_signal_16388 ;
    wire new_AGEMA_signal_16389 ;
    wire new_AGEMA_signal_16390 ;
    wire new_AGEMA_signal_16391 ;
    wire new_AGEMA_signal_16392 ;
    wire new_AGEMA_signal_16393 ;
    wire new_AGEMA_signal_16394 ;
    wire new_AGEMA_signal_16395 ;
    wire new_AGEMA_signal_16396 ;
    wire new_AGEMA_signal_16397 ;
    wire new_AGEMA_signal_16398 ;
    wire new_AGEMA_signal_16399 ;
    wire new_AGEMA_signal_16400 ;
    wire new_AGEMA_signal_16401 ;
    wire new_AGEMA_signal_16402 ;
    wire new_AGEMA_signal_16403 ;
    wire new_AGEMA_signal_16404 ;
    wire new_AGEMA_signal_16405 ;
    wire new_AGEMA_signal_16406 ;
    wire new_AGEMA_signal_16407 ;
    wire new_AGEMA_signal_16408 ;
    wire new_AGEMA_signal_16409 ;
    wire new_AGEMA_signal_16410 ;
    wire new_AGEMA_signal_16411 ;
    wire new_AGEMA_signal_16412 ;
    wire new_AGEMA_signal_16413 ;
    wire new_AGEMA_signal_16414 ;
    wire new_AGEMA_signal_16415 ;
    wire new_AGEMA_signal_16416 ;
    wire new_AGEMA_signal_16417 ;
    wire new_AGEMA_signal_16418 ;
    wire new_AGEMA_signal_16419 ;
    wire new_AGEMA_signal_16420 ;
    wire new_AGEMA_signal_16421 ;
    wire new_AGEMA_signal_16422 ;
    wire new_AGEMA_signal_16423 ;
    wire new_AGEMA_signal_16424 ;
    wire new_AGEMA_signal_16425 ;
    wire new_AGEMA_signal_16426 ;
    wire new_AGEMA_signal_16427 ;
    wire new_AGEMA_signal_16428 ;
    wire new_AGEMA_signal_16429 ;
    wire new_AGEMA_signal_16430 ;
    wire new_AGEMA_signal_16431 ;
    wire new_AGEMA_signal_16432 ;
    wire new_AGEMA_signal_16433 ;
    wire new_AGEMA_signal_16434 ;
    wire new_AGEMA_signal_16435 ;
    wire new_AGEMA_signal_16436 ;
    wire new_AGEMA_signal_16437 ;
    wire new_AGEMA_signal_16438 ;
    wire new_AGEMA_signal_16439 ;
    wire new_AGEMA_signal_16440 ;
    wire new_AGEMA_signal_16441 ;
    wire new_AGEMA_signal_16442 ;
    wire new_AGEMA_signal_16443 ;
    wire new_AGEMA_signal_16444 ;
    wire new_AGEMA_signal_16445 ;
    wire new_AGEMA_signal_16446 ;
    wire new_AGEMA_signal_16447 ;
    wire new_AGEMA_signal_16448 ;
    wire new_AGEMA_signal_16449 ;
    wire new_AGEMA_signal_16450 ;
    wire new_AGEMA_signal_16451 ;
    wire new_AGEMA_signal_16452 ;
    wire new_AGEMA_signal_16453 ;
    wire new_AGEMA_signal_16454 ;
    wire new_AGEMA_signal_16455 ;
    wire new_AGEMA_signal_16456 ;
    wire new_AGEMA_signal_16457 ;
    wire new_AGEMA_signal_16458 ;
    wire new_AGEMA_signal_16459 ;
    wire new_AGEMA_signal_16460 ;
    wire new_AGEMA_signal_16461 ;
    wire new_AGEMA_signal_16462 ;
    wire new_AGEMA_signal_16463 ;
    wire new_AGEMA_signal_16464 ;
    wire new_AGEMA_signal_16465 ;
    wire new_AGEMA_signal_16466 ;
    wire new_AGEMA_signal_16467 ;
    wire new_AGEMA_signal_16468 ;
    wire new_AGEMA_signal_16469 ;
    wire new_AGEMA_signal_16470 ;
    wire new_AGEMA_signal_16471 ;
    wire new_AGEMA_signal_16472 ;
    wire new_AGEMA_signal_16473 ;
    wire new_AGEMA_signal_16474 ;
    wire new_AGEMA_signal_16475 ;
    wire new_AGEMA_signal_16476 ;
    wire new_AGEMA_signal_16477 ;
    wire new_AGEMA_signal_16478 ;
    wire new_AGEMA_signal_16479 ;
    wire new_AGEMA_signal_16480 ;
    wire new_AGEMA_signal_16481 ;
    wire new_AGEMA_signal_16482 ;
    wire new_AGEMA_signal_16483 ;
    wire new_AGEMA_signal_16484 ;
    wire new_AGEMA_signal_16485 ;
    wire new_AGEMA_signal_16486 ;
    wire new_AGEMA_signal_16487 ;
    wire new_AGEMA_signal_16488 ;
    wire new_AGEMA_signal_16489 ;
    wire new_AGEMA_signal_16490 ;
    wire new_AGEMA_signal_16491 ;
    wire new_AGEMA_signal_16492 ;
    wire new_AGEMA_signal_16493 ;
    wire new_AGEMA_signal_16494 ;
    wire new_AGEMA_signal_16495 ;
    wire new_AGEMA_signal_16496 ;
    wire new_AGEMA_signal_16497 ;
    wire new_AGEMA_signal_16498 ;
    wire new_AGEMA_signal_16499 ;
    wire new_AGEMA_signal_16500 ;
    wire new_AGEMA_signal_16501 ;
    wire new_AGEMA_signal_16502 ;
    wire new_AGEMA_signal_16503 ;
    wire new_AGEMA_signal_16504 ;
    wire new_AGEMA_signal_16505 ;
    wire new_AGEMA_signal_16506 ;
    wire new_AGEMA_signal_16507 ;
    wire new_AGEMA_signal_16508 ;
    wire new_AGEMA_signal_16509 ;
    wire new_AGEMA_signal_16510 ;
    wire new_AGEMA_signal_16511 ;
    wire new_AGEMA_signal_16512 ;
    wire new_AGEMA_signal_16513 ;
    wire new_AGEMA_signal_16514 ;
    wire new_AGEMA_signal_16515 ;
    wire new_AGEMA_signal_16516 ;
    wire new_AGEMA_signal_16517 ;
    wire new_AGEMA_signal_16518 ;
    wire new_AGEMA_signal_16519 ;
    wire new_AGEMA_signal_16520 ;
    wire new_AGEMA_signal_16521 ;
    wire new_AGEMA_signal_16522 ;
    wire new_AGEMA_signal_16523 ;
    wire new_AGEMA_signal_16524 ;
    wire new_AGEMA_signal_16525 ;
    wire new_AGEMA_signal_16526 ;
    wire new_AGEMA_signal_16527 ;
    wire new_AGEMA_signal_16528 ;
    wire new_AGEMA_signal_16529 ;
    wire new_AGEMA_signal_16530 ;
    wire new_AGEMA_signal_16531 ;
    wire new_AGEMA_signal_16532 ;
    wire new_AGEMA_signal_16533 ;
    wire new_AGEMA_signal_16534 ;
    wire new_AGEMA_signal_16535 ;
    wire new_AGEMA_signal_16536 ;
    wire new_AGEMA_signal_16537 ;
    wire new_AGEMA_signal_16538 ;
    wire new_AGEMA_signal_16539 ;
    wire new_AGEMA_signal_16540 ;
    wire new_AGEMA_signal_16541 ;
    wire new_AGEMA_signal_16542 ;
    wire new_AGEMA_signal_16543 ;
    wire new_AGEMA_signal_16544 ;
    wire new_AGEMA_signal_16545 ;
    wire new_AGEMA_signal_16546 ;
    wire new_AGEMA_signal_16547 ;
    wire new_AGEMA_signal_16548 ;
    wire new_AGEMA_signal_16549 ;
    wire new_AGEMA_signal_16550 ;
    wire new_AGEMA_signal_16551 ;
    wire new_AGEMA_signal_16552 ;
    wire new_AGEMA_signal_16553 ;
    wire new_AGEMA_signal_16554 ;
    wire new_AGEMA_signal_16555 ;
    wire new_AGEMA_signal_16556 ;
    wire new_AGEMA_signal_16557 ;
    wire new_AGEMA_signal_16558 ;
    wire new_AGEMA_signal_16559 ;
    wire new_AGEMA_signal_16560 ;
    wire new_AGEMA_signal_16561 ;
    wire new_AGEMA_signal_16562 ;
    wire new_AGEMA_signal_16563 ;
    wire new_AGEMA_signal_16564 ;
    wire new_AGEMA_signal_16565 ;
    wire new_AGEMA_signal_16566 ;
    wire new_AGEMA_signal_16567 ;
    wire new_AGEMA_signal_16568 ;
    wire new_AGEMA_signal_16569 ;
    wire new_AGEMA_signal_16570 ;
    wire new_AGEMA_signal_16571 ;
    wire new_AGEMA_signal_16572 ;
    wire new_AGEMA_signal_16573 ;
    wire new_AGEMA_signal_16574 ;
    wire new_AGEMA_signal_16575 ;
    wire new_AGEMA_signal_16576 ;
    wire new_AGEMA_signal_16577 ;
    wire new_AGEMA_signal_16578 ;
    wire new_AGEMA_signal_16579 ;
    wire new_AGEMA_signal_16580 ;
    wire new_AGEMA_signal_16581 ;
    wire new_AGEMA_signal_16582 ;
    wire new_AGEMA_signal_16583 ;
    wire new_AGEMA_signal_16584 ;
    wire new_AGEMA_signal_16585 ;
    wire new_AGEMA_signal_16586 ;
    wire new_AGEMA_signal_16587 ;
    wire new_AGEMA_signal_16588 ;
    wire new_AGEMA_signal_16589 ;
    wire new_AGEMA_signal_16590 ;
    wire new_AGEMA_signal_16591 ;
    wire new_AGEMA_signal_16592 ;
    wire new_AGEMA_signal_16593 ;
    wire new_AGEMA_signal_16594 ;
    wire new_AGEMA_signal_16595 ;
    wire new_AGEMA_signal_16596 ;
    wire new_AGEMA_signal_16597 ;
    wire new_AGEMA_signal_16598 ;
    wire new_AGEMA_signal_16599 ;
    wire new_AGEMA_signal_16600 ;
    wire new_AGEMA_signal_16601 ;
    wire new_AGEMA_signal_16602 ;
    wire new_AGEMA_signal_16603 ;
    wire new_AGEMA_signal_16604 ;
    wire new_AGEMA_signal_16605 ;
    wire new_AGEMA_signal_16606 ;
    wire new_AGEMA_signal_16607 ;
    wire new_AGEMA_signal_16608 ;
    wire new_AGEMA_signal_16609 ;
    wire new_AGEMA_signal_16610 ;
    wire new_AGEMA_signal_16611 ;
    wire new_AGEMA_signal_16612 ;
    wire new_AGEMA_signal_16613 ;
    wire new_AGEMA_signal_16614 ;
    wire new_AGEMA_signal_16615 ;
    wire new_AGEMA_signal_16616 ;
    wire new_AGEMA_signal_16617 ;
    wire new_AGEMA_signal_16618 ;
    wire new_AGEMA_signal_16619 ;
    wire new_AGEMA_signal_16620 ;
    wire new_AGEMA_signal_16621 ;
    wire new_AGEMA_signal_16622 ;
    wire new_AGEMA_signal_16623 ;
    wire new_AGEMA_signal_16624 ;
    wire new_AGEMA_signal_16625 ;
    wire new_AGEMA_signal_16626 ;
    wire new_AGEMA_signal_16627 ;
    wire new_AGEMA_signal_16628 ;
    wire new_AGEMA_signal_16629 ;
    wire new_AGEMA_signal_16630 ;
    wire new_AGEMA_signal_16631 ;
    wire new_AGEMA_signal_16632 ;
    wire new_AGEMA_signal_16633 ;
    wire new_AGEMA_signal_16634 ;
    wire new_AGEMA_signal_16635 ;
    wire new_AGEMA_signal_16636 ;
    wire new_AGEMA_signal_16637 ;
    wire new_AGEMA_signal_16638 ;
    wire new_AGEMA_signal_16639 ;
    wire new_AGEMA_signal_16640 ;
    wire new_AGEMA_signal_16641 ;
    wire new_AGEMA_signal_16642 ;
    wire new_AGEMA_signal_16643 ;
    wire new_AGEMA_signal_16644 ;
    wire new_AGEMA_signal_16645 ;
    wire new_AGEMA_signal_16646 ;
    wire new_AGEMA_signal_16647 ;
    wire new_AGEMA_signal_16648 ;
    wire new_AGEMA_signal_16649 ;
    wire new_AGEMA_signal_16650 ;
    wire new_AGEMA_signal_16651 ;
    wire new_AGEMA_signal_16652 ;
    wire new_AGEMA_signal_16653 ;
    wire new_AGEMA_signal_16654 ;
    wire new_AGEMA_signal_16655 ;
    wire new_AGEMA_signal_16656 ;
    wire new_AGEMA_signal_16657 ;
    wire new_AGEMA_signal_16658 ;
    wire new_AGEMA_signal_16659 ;
    wire new_AGEMA_signal_16660 ;
    wire new_AGEMA_signal_16661 ;
    wire new_AGEMA_signal_16662 ;
    wire new_AGEMA_signal_16663 ;
    wire new_AGEMA_signal_16664 ;
    wire new_AGEMA_signal_16665 ;
    wire new_AGEMA_signal_16666 ;
    wire new_AGEMA_signal_16667 ;
    wire new_AGEMA_signal_16668 ;
    wire new_AGEMA_signal_16669 ;
    wire new_AGEMA_signal_16670 ;
    wire new_AGEMA_signal_16671 ;
    wire new_AGEMA_signal_16672 ;
    wire new_AGEMA_signal_16673 ;
    wire new_AGEMA_signal_16674 ;
    wire new_AGEMA_signal_16675 ;
    wire new_AGEMA_signal_16676 ;
    wire new_AGEMA_signal_16677 ;
    wire new_AGEMA_signal_16678 ;
    wire new_AGEMA_signal_16679 ;
    wire new_AGEMA_signal_16680 ;
    wire new_AGEMA_signal_16681 ;
    wire new_AGEMA_signal_16682 ;
    wire new_AGEMA_signal_16683 ;
    wire new_AGEMA_signal_16684 ;
    wire new_AGEMA_signal_16685 ;
    wire new_AGEMA_signal_16686 ;
    wire new_AGEMA_signal_16687 ;
    wire new_AGEMA_signal_16688 ;
    wire new_AGEMA_signal_16689 ;
    wire new_AGEMA_signal_16690 ;
    wire new_AGEMA_signal_16691 ;
    wire new_AGEMA_signal_16692 ;
    wire new_AGEMA_signal_16693 ;
    wire new_AGEMA_signal_16694 ;
    wire new_AGEMA_signal_16695 ;
    wire new_AGEMA_signal_16696 ;
    wire new_AGEMA_signal_16697 ;
    wire new_AGEMA_signal_16698 ;
    wire new_AGEMA_signal_16699 ;
    wire new_AGEMA_signal_16700 ;
    wire new_AGEMA_signal_16701 ;
    wire new_AGEMA_signal_16702 ;
    wire new_AGEMA_signal_16703 ;
    wire new_AGEMA_signal_16704 ;
    wire new_AGEMA_signal_16705 ;
    wire new_AGEMA_signal_16706 ;
    wire new_AGEMA_signal_16707 ;
    wire new_AGEMA_signal_16708 ;
    wire new_AGEMA_signal_16709 ;
    wire new_AGEMA_signal_16710 ;
    wire new_AGEMA_signal_16711 ;
    wire new_AGEMA_signal_16712 ;
    wire new_AGEMA_signal_16713 ;
    wire new_AGEMA_signal_16714 ;
    wire new_AGEMA_signal_16715 ;
    wire new_AGEMA_signal_16716 ;
    wire new_AGEMA_signal_16717 ;
    wire new_AGEMA_signal_16718 ;
    wire new_AGEMA_signal_16719 ;
    wire new_AGEMA_signal_16720 ;
    wire new_AGEMA_signal_16721 ;
    wire new_AGEMA_signal_16722 ;
    wire new_AGEMA_signal_16723 ;
    wire new_AGEMA_signal_16724 ;
    wire new_AGEMA_signal_16725 ;
    wire new_AGEMA_signal_16726 ;
    wire new_AGEMA_signal_16727 ;
    wire new_AGEMA_signal_16728 ;
    wire new_AGEMA_signal_16729 ;
    wire new_AGEMA_signal_16730 ;
    wire new_AGEMA_signal_16731 ;
    wire new_AGEMA_signal_16732 ;
    wire new_AGEMA_signal_16733 ;
    wire new_AGEMA_signal_16734 ;
    wire new_AGEMA_signal_16735 ;
    wire new_AGEMA_signal_16736 ;
    wire new_AGEMA_signal_16737 ;
    wire new_AGEMA_signal_16738 ;
    wire new_AGEMA_signal_16739 ;
    wire new_AGEMA_signal_16740 ;
    wire new_AGEMA_signal_16741 ;
    wire new_AGEMA_signal_16742 ;
    wire new_AGEMA_signal_16743 ;
    wire new_AGEMA_signal_16744 ;
    wire new_AGEMA_signal_16745 ;
    wire new_AGEMA_signal_16746 ;
    wire new_AGEMA_signal_16747 ;
    wire new_AGEMA_signal_16748 ;
    wire new_AGEMA_signal_16749 ;
    wire new_AGEMA_signal_16750 ;
    wire new_AGEMA_signal_16751 ;
    wire new_AGEMA_signal_16752 ;
    wire new_AGEMA_signal_16753 ;
    wire new_AGEMA_signal_16754 ;
    wire new_AGEMA_signal_16755 ;
    wire new_AGEMA_signal_16756 ;
    wire new_AGEMA_signal_16757 ;
    wire new_AGEMA_signal_16758 ;
    wire new_AGEMA_signal_16759 ;
    wire new_AGEMA_signal_16760 ;
    wire new_AGEMA_signal_16761 ;
    wire new_AGEMA_signal_16762 ;
    wire new_AGEMA_signal_16763 ;
    wire new_AGEMA_signal_16764 ;
    wire new_AGEMA_signal_16765 ;
    wire new_AGEMA_signal_16766 ;
    wire new_AGEMA_signal_16767 ;
    wire new_AGEMA_signal_16768 ;
    wire new_AGEMA_signal_16769 ;
    wire new_AGEMA_signal_16770 ;
    wire new_AGEMA_signal_16771 ;
    wire new_AGEMA_signal_16772 ;
    wire new_AGEMA_signal_16773 ;
    wire new_AGEMA_signal_16774 ;
    wire new_AGEMA_signal_16775 ;
    wire new_AGEMA_signal_16776 ;
    wire new_AGEMA_signal_16777 ;
    wire new_AGEMA_signal_16778 ;
    wire new_AGEMA_signal_16779 ;
    wire new_AGEMA_signal_16780 ;
    wire new_AGEMA_signal_16781 ;
    wire new_AGEMA_signal_16782 ;
    wire new_AGEMA_signal_16783 ;
    wire new_AGEMA_signal_16784 ;
    wire new_AGEMA_signal_16785 ;
    wire new_AGEMA_signal_16786 ;
    wire new_AGEMA_signal_16787 ;
    wire new_AGEMA_signal_16788 ;
    wire new_AGEMA_signal_16789 ;
    wire new_AGEMA_signal_16790 ;
    wire new_AGEMA_signal_16791 ;
    wire new_AGEMA_signal_16792 ;
    wire new_AGEMA_signal_16793 ;
    wire new_AGEMA_signal_16794 ;
    wire new_AGEMA_signal_16795 ;
    wire new_AGEMA_signal_16796 ;
    wire new_AGEMA_signal_16797 ;
    wire new_AGEMA_signal_16798 ;
    wire new_AGEMA_signal_16799 ;
    wire new_AGEMA_signal_16800 ;
    wire new_AGEMA_signal_16801 ;
    wire new_AGEMA_signal_16802 ;
    wire new_AGEMA_signal_16803 ;
    wire new_AGEMA_signal_16804 ;
    wire new_AGEMA_signal_16805 ;
    wire new_AGEMA_signal_16806 ;
    wire new_AGEMA_signal_16807 ;
    wire new_AGEMA_signal_16808 ;
    wire new_AGEMA_signal_16809 ;
    wire new_AGEMA_signal_16810 ;
    wire new_AGEMA_signal_16811 ;
    wire new_AGEMA_signal_16812 ;
    wire new_AGEMA_signal_16813 ;
    wire new_AGEMA_signal_16814 ;
    wire new_AGEMA_signal_16815 ;
    wire new_AGEMA_signal_16816 ;
    wire new_AGEMA_signal_16817 ;
    wire new_AGEMA_signal_16818 ;
    wire new_AGEMA_signal_16819 ;
    wire new_AGEMA_signal_16820 ;
    wire new_AGEMA_signal_16821 ;
    wire new_AGEMA_signal_16822 ;
    wire new_AGEMA_signal_16823 ;
    wire new_AGEMA_signal_16824 ;
    wire new_AGEMA_signal_16825 ;
    wire new_AGEMA_signal_16826 ;
    wire new_AGEMA_signal_16827 ;
    wire new_AGEMA_signal_16828 ;
    wire new_AGEMA_signal_16829 ;
    wire new_AGEMA_signal_16830 ;
    wire new_AGEMA_signal_16831 ;
    wire new_AGEMA_signal_16832 ;
    wire new_AGEMA_signal_16833 ;
    wire new_AGEMA_signal_16834 ;
    wire new_AGEMA_signal_16835 ;
    wire new_AGEMA_signal_16836 ;
    wire new_AGEMA_signal_16837 ;
    wire new_AGEMA_signal_16838 ;
    wire new_AGEMA_signal_16839 ;
    wire new_AGEMA_signal_16840 ;
    wire new_AGEMA_signal_16841 ;
    wire new_AGEMA_signal_16842 ;
    wire new_AGEMA_signal_16843 ;
    wire new_AGEMA_signal_16844 ;
    wire new_AGEMA_signal_16845 ;
    wire new_AGEMA_signal_16846 ;
    wire new_AGEMA_signal_16847 ;
    wire new_AGEMA_signal_16848 ;
    wire new_AGEMA_signal_16849 ;
    wire new_AGEMA_signal_16850 ;
    wire new_AGEMA_signal_16851 ;
    wire new_AGEMA_signal_16852 ;
    wire new_AGEMA_signal_16853 ;
    wire new_AGEMA_signal_16854 ;
    wire new_AGEMA_signal_16855 ;
    wire new_AGEMA_signal_16856 ;
    wire new_AGEMA_signal_16857 ;
    wire new_AGEMA_signal_16858 ;
    wire new_AGEMA_signal_16859 ;
    wire new_AGEMA_signal_16860 ;
    wire new_AGEMA_signal_16861 ;
    wire new_AGEMA_signal_16862 ;
    wire new_AGEMA_signal_16863 ;
    wire new_AGEMA_signal_16864 ;
    wire new_AGEMA_signal_16865 ;
    wire new_AGEMA_signal_16866 ;
    wire new_AGEMA_signal_16867 ;
    wire new_AGEMA_signal_16868 ;
    wire new_AGEMA_signal_16869 ;
    wire new_AGEMA_signal_16870 ;
    wire new_AGEMA_signal_16871 ;
    wire new_AGEMA_signal_16872 ;
    wire new_AGEMA_signal_16873 ;
    wire new_AGEMA_signal_16874 ;
    wire new_AGEMA_signal_16875 ;
    wire new_AGEMA_signal_16876 ;
    wire new_AGEMA_signal_16877 ;
    wire new_AGEMA_signal_16878 ;
    wire new_AGEMA_signal_16879 ;
    wire new_AGEMA_signal_16880 ;
    wire new_AGEMA_signal_16881 ;
    wire new_AGEMA_signal_16882 ;
    wire new_AGEMA_signal_16883 ;
    wire new_AGEMA_signal_16884 ;
    wire new_AGEMA_signal_16885 ;
    wire new_AGEMA_signal_16886 ;
    wire new_AGEMA_signal_16887 ;
    wire new_AGEMA_signal_16888 ;
    wire new_AGEMA_signal_16889 ;
    wire new_AGEMA_signal_16890 ;
    wire new_AGEMA_signal_16891 ;
    wire new_AGEMA_signal_16892 ;
    wire new_AGEMA_signal_16893 ;
    wire new_AGEMA_signal_16894 ;
    wire new_AGEMA_signal_16895 ;
    wire new_AGEMA_signal_16896 ;
    wire new_AGEMA_signal_16897 ;
    wire new_AGEMA_signal_16898 ;
    wire new_AGEMA_signal_16899 ;
    wire new_AGEMA_signal_16900 ;
    wire new_AGEMA_signal_16901 ;
    wire new_AGEMA_signal_16902 ;
    wire new_AGEMA_signal_16903 ;
    wire new_AGEMA_signal_16904 ;
    wire new_AGEMA_signal_16905 ;
    wire new_AGEMA_signal_16906 ;
    wire new_AGEMA_signal_16907 ;
    wire new_AGEMA_signal_16908 ;
    wire new_AGEMA_signal_16909 ;
    wire new_AGEMA_signal_16910 ;
    wire new_AGEMA_signal_16911 ;
    wire new_AGEMA_signal_16912 ;
    wire new_AGEMA_signal_16913 ;
    wire new_AGEMA_signal_16914 ;
    wire new_AGEMA_signal_16915 ;
    wire new_AGEMA_signal_16916 ;
    wire new_AGEMA_signal_16917 ;
    wire new_AGEMA_signal_16918 ;
    wire new_AGEMA_signal_16919 ;
    wire new_AGEMA_signal_16920 ;
    wire new_AGEMA_signal_16921 ;
    wire new_AGEMA_signal_16922 ;
    wire new_AGEMA_signal_16923 ;
    wire new_AGEMA_signal_16924 ;
    wire new_AGEMA_signal_16925 ;
    wire new_AGEMA_signal_16926 ;
    wire new_AGEMA_signal_16927 ;
    wire new_AGEMA_signal_16928 ;
    wire new_AGEMA_signal_16929 ;
    wire new_AGEMA_signal_16930 ;
    wire new_AGEMA_signal_16931 ;
    wire new_AGEMA_signal_16932 ;
    wire new_AGEMA_signal_16933 ;
    wire new_AGEMA_signal_16934 ;
    wire new_AGEMA_signal_16935 ;
    wire new_AGEMA_signal_16936 ;
    wire new_AGEMA_signal_16937 ;
    wire new_AGEMA_signal_16938 ;
    wire new_AGEMA_signal_16939 ;
    wire new_AGEMA_signal_16940 ;
    wire new_AGEMA_signal_16941 ;
    wire new_AGEMA_signal_16942 ;
    wire new_AGEMA_signal_16943 ;
    wire new_AGEMA_signal_16944 ;
    wire new_AGEMA_signal_16945 ;
    wire new_AGEMA_signal_16946 ;
    wire new_AGEMA_signal_16947 ;
    wire new_AGEMA_signal_16948 ;
    wire new_AGEMA_signal_16949 ;
    wire new_AGEMA_signal_16950 ;
    wire new_AGEMA_signal_16951 ;
    wire new_AGEMA_signal_16952 ;
    wire new_AGEMA_signal_16953 ;
    wire new_AGEMA_signal_16954 ;
    wire new_AGEMA_signal_16955 ;
    wire new_AGEMA_signal_16956 ;
    wire new_AGEMA_signal_16957 ;
    wire new_AGEMA_signal_16958 ;
    wire new_AGEMA_signal_16959 ;
    wire new_AGEMA_signal_16960 ;
    wire new_AGEMA_signal_16961 ;
    wire new_AGEMA_signal_16962 ;
    wire new_AGEMA_signal_16963 ;
    wire new_AGEMA_signal_16964 ;
    wire new_AGEMA_signal_16965 ;
    wire new_AGEMA_signal_16966 ;
    wire new_AGEMA_signal_16967 ;
    wire new_AGEMA_signal_16968 ;
    wire new_AGEMA_signal_16969 ;
    wire new_AGEMA_signal_16970 ;
    wire new_AGEMA_signal_16971 ;
    wire new_AGEMA_signal_16972 ;
    wire new_AGEMA_signal_16973 ;
    wire new_AGEMA_signal_16974 ;
    wire new_AGEMA_signal_16975 ;
    wire new_AGEMA_signal_16976 ;
    wire new_AGEMA_signal_16977 ;
    wire new_AGEMA_signal_16978 ;
    wire new_AGEMA_signal_16979 ;
    wire new_AGEMA_signal_16980 ;
    wire new_AGEMA_signal_16981 ;
    wire new_AGEMA_signal_16982 ;
    wire new_AGEMA_signal_16983 ;
    wire new_AGEMA_signal_16984 ;
    wire new_AGEMA_signal_16985 ;
    wire new_AGEMA_signal_16986 ;
    wire new_AGEMA_signal_16987 ;
    wire new_AGEMA_signal_16988 ;
    wire new_AGEMA_signal_16989 ;
    wire new_AGEMA_signal_16990 ;
    wire new_AGEMA_signal_16991 ;
    wire new_AGEMA_signal_16992 ;
    wire new_AGEMA_signal_16993 ;
    wire new_AGEMA_signal_16994 ;
    wire new_AGEMA_signal_16995 ;
    wire new_AGEMA_signal_16996 ;
    wire new_AGEMA_signal_16997 ;
    wire new_AGEMA_signal_16998 ;
    wire new_AGEMA_signal_16999 ;
    wire new_AGEMA_signal_17000 ;
    wire new_AGEMA_signal_17001 ;
    wire new_AGEMA_signal_17002 ;
    wire new_AGEMA_signal_17003 ;
    wire new_AGEMA_signal_17004 ;
    wire new_AGEMA_signal_17005 ;
    wire new_AGEMA_signal_17006 ;
    wire new_AGEMA_signal_17007 ;
    wire new_AGEMA_signal_17008 ;
    wire new_AGEMA_signal_17009 ;
    wire new_AGEMA_signal_17010 ;
    wire new_AGEMA_signal_17011 ;
    wire new_AGEMA_signal_17012 ;
    wire new_AGEMA_signal_17013 ;
    wire new_AGEMA_signal_17014 ;
    wire new_AGEMA_signal_17015 ;
    wire new_AGEMA_signal_17016 ;
    wire new_AGEMA_signal_17017 ;
    wire new_AGEMA_signal_17018 ;
    wire new_AGEMA_signal_17019 ;
    wire new_AGEMA_signal_17020 ;
    wire new_AGEMA_signal_17021 ;
    wire new_AGEMA_signal_17022 ;
    wire new_AGEMA_signal_17023 ;
    wire new_AGEMA_signal_17024 ;
    wire new_AGEMA_signal_17025 ;
    wire new_AGEMA_signal_17026 ;
    wire new_AGEMA_signal_17027 ;
    wire new_AGEMA_signal_17028 ;
    wire new_AGEMA_signal_17029 ;
    wire new_AGEMA_signal_17030 ;
    wire new_AGEMA_signal_17031 ;
    wire new_AGEMA_signal_17032 ;
    wire new_AGEMA_signal_17033 ;
    wire new_AGEMA_signal_17034 ;
    wire new_AGEMA_signal_17035 ;
    wire new_AGEMA_signal_17036 ;
    wire new_AGEMA_signal_17037 ;
    wire new_AGEMA_signal_17038 ;
    wire new_AGEMA_signal_17039 ;
    wire new_AGEMA_signal_17040 ;
    wire new_AGEMA_signal_17041 ;
    wire new_AGEMA_signal_17042 ;
    wire new_AGEMA_signal_17043 ;
    wire new_AGEMA_signal_17044 ;
    wire new_AGEMA_signal_17045 ;
    wire new_AGEMA_signal_17046 ;
    wire new_AGEMA_signal_17047 ;
    wire new_AGEMA_signal_17048 ;
    wire new_AGEMA_signal_17049 ;
    wire new_AGEMA_signal_17050 ;
    wire new_AGEMA_signal_17051 ;
    wire new_AGEMA_signal_17052 ;
    wire new_AGEMA_signal_17053 ;
    wire new_AGEMA_signal_17054 ;
    wire new_AGEMA_signal_17055 ;
    wire new_AGEMA_signal_17056 ;
    wire new_AGEMA_signal_17057 ;
    wire new_AGEMA_signal_17058 ;
    wire new_AGEMA_signal_17059 ;
    wire new_AGEMA_signal_17060 ;
    wire new_AGEMA_signal_17061 ;
    wire new_AGEMA_signal_17062 ;
    wire new_AGEMA_signal_17063 ;
    wire new_AGEMA_signal_17064 ;
    wire new_AGEMA_signal_17065 ;
    wire new_AGEMA_signal_17066 ;
    wire new_AGEMA_signal_17067 ;
    wire new_AGEMA_signal_17068 ;
    wire new_AGEMA_signal_17069 ;
    wire new_AGEMA_signal_17070 ;
    wire new_AGEMA_signal_17071 ;
    wire new_AGEMA_signal_17072 ;
    wire new_AGEMA_signal_17073 ;
    wire new_AGEMA_signal_17074 ;
    wire new_AGEMA_signal_17075 ;
    wire new_AGEMA_signal_17076 ;
    wire new_AGEMA_signal_17077 ;
    wire new_AGEMA_signal_17078 ;
    wire new_AGEMA_signal_17079 ;
    wire new_AGEMA_signal_17080 ;
    wire new_AGEMA_signal_17081 ;
    wire new_AGEMA_signal_17082 ;
    wire new_AGEMA_signal_17083 ;
    wire new_AGEMA_signal_17084 ;
    wire new_AGEMA_signal_17085 ;
    wire new_AGEMA_signal_17086 ;
    wire new_AGEMA_signal_17087 ;
    wire new_AGEMA_signal_17088 ;
    wire new_AGEMA_signal_17089 ;
    wire new_AGEMA_signal_17090 ;
    wire new_AGEMA_signal_17091 ;
    wire new_AGEMA_signal_17092 ;
    wire new_AGEMA_signal_17093 ;
    wire new_AGEMA_signal_17094 ;
    wire new_AGEMA_signal_17095 ;
    wire new_AGEMA_signal_17096 ;
    wire new_AGEMA_signal_17097 ;
    wire new_AGEMA_signal_17098 ;
    wire new_AGEMA_signal_17099 ;
    wire new_AGEMA_signal_17100 ;
    wire new_AGEMA_signal_17101 ;
    wire new_AGEMA_signal_17102 ;
    wire new_AGEMA_signal_17103 ;
    wire new_AGEMA_signal_17104 ;
    wire new_AGEMA_signal_17105 ;
    wire new_AGEMA_signal_17106 ;
    wire new_AGEMA_signal_17107 ;
    wire new_AGEMA_signal_17108 ;
    wire new_AGEMA_signal_17109 ;
    wire new_AGEMA_signal_17110 ;
    wire new_AGEMA_signal_17111 ;
    wire new_AGEMA_signal_17112 ;
    wire new_AGEMA_signal_17113 ;
    wire new_AGEMA_signal_17114 ;
    wire new_AGEMA_signal_17115 ;
    wire new_AGEMA_signal_17116 ;
    wire new_AGEMA_signal_17117 ;
    wire new_AGEMA_signal_17118 ;
    wire new_AGEMA_signal_17119 ;
    wire new_AGEMA_signal_17120 ;
    wire new_AGEMA_signal_17121 ;
    wire new_AGEMA_signal_17122 ;
    wire new_AGEMA_signal_17123 ;
    wire new_AGEMA_signal_17124 ;
    wire new_AGEMA_signal_17125 ;
    wire new_AGEMA_signal_17126 ;
    wire new_AGEMA_signal_17127 ;
    wire new_AGEMA_signal_17128 ;
    wire new_AGEMA_signal_17129 ;
    wire new_AGEMA_signal_17130 ;
    wire new_AGEMA_signal_17131 ;
    wire new_AGEMA_signal_17132 ;
    wire new_AGEMA_signal_17133 ;
    wire new_AGEMA_signal_17134 ;
    wire new_AGEMA_signal_17135 ;
    wire new_AGEMA_signal_17136 ;
    wire new_AGEMA_signal_17137 ;
    wire new_AGEMA_signal_17138 ;
    wire new_AGEMA_signal_17139 ;
    wire new_AGEMA_signal_17140 ;
    wire new_AGEMA_signal_17141 ;
    wire new_AGEMA_signal_17142 ;
    wire new_AGEMA_signal_17143 ;
    wire new_AGEMA_signal_17144 ;
    wire new_AGEMA_signal_17145 ;
    wire new_AGEMA_signal_17146 ;
    wire new_AGEMA_signal_17147 ;
    wire new_AGEMA_signal_17148 ;
    wire new_AGEMA_signal_17149 ;
    wire new_AGEMA_signal_17150 ;
    wire new_AGEMA_signal_17151 ;
    wire new_AGEMA_signal_17152 ;
    wire new_AGEMA_signal_17153 ;
    wire new_AGEMA_signal_17154 ;
    wire new_AGEMA_signal_17155 ;
    wire new_AGEMA_signal_17156 ;
    wire new_AGEMA_signal_17157 ;
    wire new_AGEMA_signal_17158 ;
    wire new_AGEMA_signal_17159 ;
    wire new_AGEMA_signal_17160 ;
    wire new_AGEMA_signal_17161 ;
    wire new_AGEMA_signal_17162 ;
    wire new_AGEMA_signal_17163 ;
    wire new_AGEMA_signal_17164 ;
    wire new_AGEMA_signal_17165 ;
    wire new_AGEMA_signal_17166 ;
    wire new_AGEMA_signal_17167 ;
    wire new_AGEMA_signal_17168 ;
    wire new_AGEMA_signal_17169 ;
    wire new_AGEMA_signal_17170 ;
    wire new_AGEMA_signal_17171 ;
    wire new_AGEMA_signal_17172 ;
    wire new_AGEMA_signal_17173 ;
    wire new_AGEMA_signal_17174 ;
    wire new_AGEMA_signal_17175 ;
    wire new_AGEMA_signal_17176 ;
    wire new_AGEMA_signal_17177 ;
    wire new_AGEMA_signal_17178 ;
    wire new_AGEMA_signal_17179 ;
    wire new_AGEMA_signal_17180 ;
    wire new_AGEMA_signal_17181 ;
    wire new_AGEMA_signal_17182 ;
    wire new_AGEMA_signal_17183 ;
    wire new_AGEMA_signal_17184 ;
    wire new_AGEMA_signal_17185 ;
    wire new_AGEMA_signal_17186 ;
    wire new_AGEMA_signal_17187 ;
    wire new_AGEMA_signal_17188 ;
    wire new_AGEMA_signal_17189 ;
    wire new_AGEMA_signal_17190 ;
    wire new_AGEMA_signal_17191 ;
    wire new_AGEMA_signal_17192 ;
    wire new_AGEMA_signal_17193 ;
    wire new_AGEMA_signal_17194 ;
    wire new_AGEMA_signal_17195 ;
    wire new_AGEMA_signal_17196 ;
    wire new_AGEMA_signal_17197 ;
    wire new_AGEMA_signal_17198 ;
    wire new_AGEMA_signal_17199 ;
    wire new_AGEMA_signal_17200 ;
    wire new_AGEMA_signal_17201 ;
    wire new_AGEMA_signal_17202 ;
    wire new_AGEMA_signal_17203 ;
    wire new_AGEMA_signal_17204 ;
    wire new_AGEMA_signal_17205 ;
    wire new_AGEMA_signal_17206 ;
    wire new_AGEMA_signal_17207 ;
    wire new_AGEMA_signal_17208 ;
    wire new_AGEMA_signal_17209 ;
    wire new_AGEMA_signal_17210 ;
    wire new_AGEMA_signal_17211 ;
    wire new_AGEMA_signal_17212 ;
    wire new_AGEMA_signal_17213 ;
    wire new_AGEMA_signal_17214 ;
    wire new_AGEMA_signal_17215 ;
    wire new_AGEMA_signal_17216 ;
    wire new_AGEMA_signal_17217 ;
    wire new_AGEMA_signal_17218 ;
    wire new_AGEMA_signal_17219 ;
    wire new_AGEMA_signal_17220 ;
    wire new_AGEMA_signal_17221 ;
    wire new_AGEMA_signal_17222 ;
    wire new_AGEMA_signal_17223 ;
    wire new_AGEMA_signal_17224 ;
    wire new_AGEMA_signal_17225 ;
    wire new_AGEMA_signal_17226 ;
    wire new_AGEMA_signal_17227 ;
    wire new_AGEMA_signal_17228 ;
    wire new_AGEMA_signal_17229 ;
    wire new_AGEMA_signal_17230 ;
    wire new_AGEMA_signal_17231 ;
    wire new_AGEMA_signal_17232 ;
    wire new_AGEMA_signal_17233 ;
    wire new_AGEMA_signal_17234 ;
    wire new_AGEMA_signal_17235 ;
    wire new_AGEMA_signal_17236 ;
    wire new_AGEMA_signal_17237 ;
    wire new_AGEMA_signal_17238 ;
    wire new_AGEMA_signal_17239 ;
    wire new_AGEMA_signal_17240 ;
    wire new_AGEMA_signal_17241 ;
    wire new_AGEMA_signal_17242 ;
    wire new_AGEMA_signal_17243 ;
    wire new_AGEMA_signal_17244 ;
    wire new_AGEMA_signal_17245 ;
    wire new_AGEMA_signal_17246 ;
    wire new_AGEMA_signal_17247 ;
    wire new_AGEMA_signal_17248 ;
    wire new_AGEMA_signal_17249 ;
    wire new_AGEMA_signal_17250 ;
    wire new_AGEMA_signal_17251 ;
    wire new_AGEMA_signal_17252 ;
    wire new_AGEMA_signal_17253 ;
    wire new_AGEMA_signal_17254 ;
    wire new_AGEMA_signal_17255 ;
    wire new_AGEMA_signal_17256 ;
    wire new_AGEMA_signal_17257 ;
    wire new_AGEMA_signal_17258 ;
    wire new_AGEMA_signal_17259 ;
    wire new_AGEMA_signal_17260 ;
    wire new_AGEMA_signal_17261 ;
    wire new_AGEMA_signal_17262 ;
    wire new_AGEMA_signal_17263 ;
    wire new_AGEMA_signal_17264 ;
    wire new_AGEMA_signal_17265 ;
    wire new_AGEMA_signal_17266 ;
    wire new_AGEMA_signal_17267 ;
    wire new_AGEMA_signal_17268 ;
    wire new_AGEMA_signal_17269 ;
    wire new_AGEMA_signal_17270 ;
    wire new_AGEMA_signal_17271 ;
    wire new_AGEMA_signal_17272 ;
    wire new_AGEMA_signal_17273 ;
    wire new_AGEMA_signal_17274 ;
    wire new_AGEMA_signal_17275 ;
    wire new_AGEMA_signal_17276 ;
    wire new_AGEMA_signal_17277 ;
    wire new_AGEMA_signal_17278 ;
    wire new_AGEMA_signal_17279 ;
    wire new_AGEMA_signal_17280 ;
    wire new_AGEMA_signal_17281 ;
    wire new_AGEMA_signal_17282 ;
    wire new_AGEMA_signal_17283 ;
    wire new_AGEMA_signal_17284 ;
    wire new_AGEMA_signal_17285 ;
    wire new_AGEMA_signal_17286 ;
    wire new_AGEMA_signal_17287 ;
    wire new_AGEMA_signal_17288 ;
    wire new_AGEMA_signal_17289 ;
    wire new_AGEMA_signal_17290 ;
    wire new_AGEMA_signal_17291 ;
    wire new_AGEMA_signal_17292 ;
    wire new_AGEMA_signal_17293 ;
    wire new_AGEMA_signal_17294 ;
    wire new_AGEMA_signal_17295 ;
    wire new_AGEMA_signal_17296 ;
    wire new_AGEMA_signal_17297 ;
    wire new_AGEMA_signal_17298 ;
    wire new_AGEMA_signal_17299 ;
    wire new_AGEMA_signal_17300 ;
    wire new_AGEMA_signal_17301 ;
    wire new_AGEMA_signal_17302 ;
    wire new_AGEMA_signal_17303 ;
    wire new_AGEMA_signal_17304 ;
    wire new_AGEMA_signal_17305 ;
    wire new_AGEMA_signal_17306 ;
    wire new_AGEMA_signal_17307 ;
    wire new_AGEMA_signal_17308 ;
    wire new_AGEMA_signal_17309 ;
    wire new_AGEMA_signal_17310 ;
    wire new_AGEMA_signal_17311 ;
    wire new_AGEMA_signal_17312 ;
    wire new_AGEMA_signal_17313 ;
    wire new_AGEMA_signal_17314 ;
    wire new_AGEMA_signal_17315 ;
    wire new_AGEMA_signal_17316 ;
    wire new_AGEMA_signal_17317 ;
    wire new_AGEMA_signal_17318 ;
    wire new_AGEMA_signal_17319 ;
    wire new_AGEMA_signal_17320 ;
    wire new_AGEMA_signal_17321 ;
    wire new_AGEMA_signal_17322 ;
    wire new_AGEMA_signal_17323 ;
    wire new_AGEMA_signal_17324 ;
    wire new_AGEMA_signal_17325 ;
    wire new_AGEMA_signal_17326 ;
    wire new_AGEMA_signal_17327 ;
    wire new_AGEMA_signal_17328 ;
    wire new_AGEMA_signal_17329 ;
    wire new_AGEMA_signal_17330 ;
    wire new_AGEMA_signal_17331 ;
    wire new_AGEMA_signal_17332 ;
    wire new_AGEMA_signal_17333 ;
    wire new_AGEMA_signal_17334 ;
    wire new_AGEMA_signal_17335 ;
    wire new_AGEMA_signal_17336 ;
    wire new_AGEMA_signal_17337 ;
    wire new_AGEMA_signal_17338 ;
    wire new_AGEMA_signal_17339 ;
    wire new_AGEMA_signal_17340 ;
    wire new_AGEMA_signal_17341 ;
    wire new_AGEMA_signal_17342 ;
    wire new_AGEMA_signal_17343 ;
    wire new_AGEMA_signal_17344 ;
    wire new_AGEMA_signal_17345 ;
    wire new_AGEMA_signal_17346 ;
    wire new_AGEMA_signal_17347 ;
    wire new_AGEMA_signal_17348 ;
    wire new_AGEMA_signal_17349 ;
    wire new_AGEMA_signal_17350 ;
    wire new_AGEMA_signal_17351 ;
    wire new_AGEMA_signal_17352 ;
    wire new_AGEMA_signal_17353 ;
    wire new_AGEMA_signal_17354 ;
    wire new_AGEMA_signal_17355 ;
    wire new_AGEMA_signal_17356 ;
    wire new_AGEMA_signal_17357 ;
    wire new_AGEMA_signal_17358 ;
    wire new_AGEMA_signal_17359 ;
    wire new_AGEMA_signal_17360 ;
    wire new_AGEMA_signal_17361 ;
    wire new_AGEMA_signal_17362 ;
    wire new_AGEMA_signal_17363 ;
    wire new_AGEMA_signal_17364 ;
    wire new_AGEMA_signal_17365 ;
    wire new_AGEMA_signal_17366 ;
    wire new_AGEMA_signal_17367 ;
    wire new_AGEMA_signal_17368 ;
    wire new_AGEMA_signal_17369 ;
    wire new_AGEMA_signal_17370 ;
    wire new_AGEMA_signal_17371 ;
    wire new_AGEMA_signal_17372 ;
    wire new_AGEMA_signal_17373 ;
    wire new_AGEMA_signal_17374 ;
    wire new_AGEMA_signal_17375 ;
    wire new_AGEMA_signal_17376 ;
    wire new_AGEMA_signal_17377 ;
    wire new_AGEMA_signal_17378 ;
    wire new_AGEMA_signal_17379 ;
    wire new_AGEMA_signal_17380 ;
    wire new_AGEMA_signal_17381 ;
    wire new_AGEMA_signal_17382 ;
    wire new_AGEMA_signal_17383 ;
    wire new_AGEMA_signal_17384 ;
    wire new_AGEMA_signal_17385 ;
    wire new_AGEMA_signal_17386 ;
    wire new_AGEMA_signal_17387 ;
    wire new_AGEMA_signal_17388 ;
    wire new_AGEMA_signal_17389 ;
    wire new_AGEMA_signal_17390 ;
    wire new_AGEMA_signal_17391 ;
    wire new_AGEMA_signal_17392 ;
    wire new_AGEMA_signal_17393 ;
    wire new_AGEMA_signal_17394 ;
    wire new_AGEMA_signal_17395 ;
    wire new_AGEMA_signal_17396 ;
    wire new_AGEMA_signal_17397 ;
    wire new_AGEMA_signal_17398 ;
    wire new_AGEMA_signal_17399 ;
    wire new_AGEMA_signal_17400 ;
    wire new_AGEMA_signal_17401 ;
    wire new_AGEMA_signal_17402 ;
    wire new_AGEMA_signal_17403 ;
    wire new_AGEMA_signal_17404 ;
    wire new_AGEMA_signal_17405 ;
    wire new_AGEMA_signal_17406 ;
    wire new_AGEMA_signal_17407 ;
    wire new_AGEMA_signal_17408 ;
    wire new_AGEMA_signal_17409 ;
    wire new_AGEMA_signal_17410 ;
    wire new_AGEMA_signal_17411 ;
    wire new_AGEMA_signal_17412 ;
    wire new_AGEMA_signal_17413 ;
    wire new_AGEMA_signal_17414 ;
    wire new_AGEMA_signal_17415 ;
    wire new_AGEMA_signal_17416 ;
    wire new_AGEMA_signal_17417 ;
    wire new_AGEMA_signal_17418 ;
    wire new_AGEMA_signal_17419 ;
    wire new_AGEMA_signal_17420 ;
    wire new_AGEMA_signal_17421 ;
    wire new_AGEMA_signal_17422 ;
    wire new_AGEMA_signal_17423 ;
    wire new_AGEMA_signal_17424 ;
    wire new_AGEMA_signal_17425 ;
    wire new_AGEMA_signal_17426 ;
    wire new_AGEMA_signal_17427 ;
    wire new_AGEMA_signal_17428 ;
    wire new_AGEMA_signal_17429 ;
    wire new_AGEMA_signal_17430 ;
    wire new_AGEMA_signal_17431 ;
    wire new_AGEMA_signal_17432 ;
    wire new_AGEMA_signal_17433 ;
    wire new_AGEMA_signal_17434 ;
    wire new_AGEMA_signal_17435 ;
    wire new_AGEMA_signal_17436 ;
    wire new_AGEMA_signal_17437 ;
    wire new_AGEMA_signal_17438 ;
    wire new_AGEMA_signal_17439 ;
    wire new_AGEMA_signal_17440 ;
    wire new_AGEMA_signal_17441 ;
    wire new_AGEMA_signal_17442 ;
    wire new_AGEMA_signal_17443 ;
    wire new_AGEMA_signal_17444 ;
    wire new_AGEMA_signal_17445 ;
    wire new_AGEMA_signal_17446 ;
    wire new_AGEMA_signal_17447 ;
    wire new_AGEMA_signal_17448 ;
    wire new_AGEMA_signal_17449 ;
    wire new_AGEMA_signal_17450 ;
    wire new_AGEMA_signal_17451 ;
    wire new_AGEMA_signal_17452 ;
    wire new_AGEMA_signal_17453 ;
    wire new_AGEMA_signal_17454 ;
    wire new_AGEMA_signal_17455 ;
    wire new_AGEMA_signal_17456 ;
    wire new_AGEMA_signal_17457 ;
    wire new_AGEMA_signal_17458 ;
    wire new_AGEMA_signal_17459 ;
    wire new_AGEMA_signal_17460 ;
    wire new_AGEMA_signal_17461 ;
    wire new_AGEMA_signal_17462 ;
    wire new_AGEMA_signal_17463 ;
    wire new_AGEMA_signal_17464 ;
    wire new_AGEMA_signal_17465 ;
    wire new_AGEMA_signal_17466 ;
    wire new_AGEMA_signal_17467 ;
    wire new_AGEMA_signal_17468 ;
    wire new_AGEMA_signal_17469 ;
    wire new_AGEMA_signal_17470 ;
    wire new_AGEMA_signal_17471 ;
    wire new_AGEMA_signal_17472 ;
    wire new_AGEMA_signal_17473 ;
    wire new_AGEMA_signal_17474 ;
    wire new_AGEMA_signal_17475 ;
    wire new_AGEMA_signal_17476 ;
    wire new_AGEMA_signal_17477 ;
    wire new_AGEMA_signal_17478 ;
    wire new_AGEMA_signal_17479 ;
    wire new_AGEMA_signal_17480 ;
    wire new_AGEMA_signal_17481 ;
    wire new_AGEMA_signal_17482 ;
    wire new_AGEMA_signal_17483 ;
    wire new_AGEMA_signal_17484 ;
    wire new_AGEMA_signal_17485 ;
    wire new_AGEMA_signal_17486 ;
    wire new_AGEMA_signal_17487 ;
    wire new_AGEMA_signal_17488 ;
    wire new_AGEMA_signal_17489 ;
    wire new_AGEMA_signal_17490 ;
    wire new_AGEMA_signal_17491 ;
    wire new_AGEMA_signal_17492 ;
    wire new_AGEMA_signal_17493 ;
    wire new_AGEMA_signal_17494 ;
    wire new_AGEMA_signal_17495 ;
    wire new_AGEMA_signal_17496 ;
    wire new_AGEMA_signal_17497 ;
    wire new_AGEMA_signal_17498 ;
    wire new_AGEMA_signal_17499 ;
    wire new_AGEMA_signal_17500 ;
    wire new_AGEMA_signal_17501 ;
    wire new_AGEMA_signal_17502 ;
    wire new_AGEMA_signal_17503 ;
    wire new_AGEMA_signal_17504 ;
    wire new_AGEMA_signal_17505 ;
    wire new_AGEMA_signal_17506 ;
    wire new_AGEMA_signal_17507 ;
    wire new_AGEMA_signal_17508 ;
    wire new_AGEMA_signal_17509 ;
    wire new_AGEMA_signal_17510 ;
    wire new_AGEMA_signal_17511 ;
    wire new_AGEMA_signal_17512 ;
    wire new_AGEMA_signal_17513 ;
    wire new_AGEMA_signal_17514 ;
    wire new_AGEMA_signal_17515 ;
    wire new_AGEMA_signal_17516 ;
    wire new_AGEMA_signal_17517 ;
    wire new_AGEMA_signal_17518 ;
    wire new_AGEMA_signal_17519 ;
    wire new_AGEMA_signal_17520 ;
    wire new_AGEMA_signal_17521 ;
    wire new_AGEMA_signal_17522 ;
    wire new_AGEMA_signal_17523 ;
    wire new_AGEMA_signal_17524 ;
    wire new_AGEMA_signal_17525 ;
    wire new_AGEMA_signal_17526 ;
    wire new_AGEMA_signal_17527 ;
    wire new_AGEMA_signal_17528 ;
    wire new_AGEMA_signal_17529 ;
    wire new_AGEMA_signal_17530 ;
    wire new_AGEMA_signal_17531 ;
    wire new_AGEMA_signal_17532 ;
    wire new_AGEMA_signal_17533 ;
    wire new_AGEMA_signal_17534 ;
    wire new_AGEMA_signal_17535 ;
    wire new_AGEMA_signal_17536 ;
    wire new_AGEMA_signal_17537 ;
    wire new_AGEMA_signal_17538 ;
    wire new_AGEMA_signal_17539 ;
    wire new_AGEMA_signal_17540 ;
    wire new_AGEMA_signal_17541 ;
    wire new_AGEMA_signal_17542 ;
    wire new_AGEMA_signal_17543 ;
    wire new_AGEMA_signal_17544 ;
    wire new_AGEMA_signal_17545 ;
    wire new_AGEMA_signal_17546 ;
    wire new_AGEMA_signal_17547 ;
    wire new_AGEMA_signal_17548 ;
    wire new_AGEMA_signal_17549 ;
    wire new_AGEMA_signal_17550 ;
    wire new_AGEMA_signal_17551 ;
    wire new_AGEMA_signal_17552 ;
    wire new_AGEMA_signal_17553 ;
    wire new_AGEMA_signal_17554 ;
    wire new_AGEMA_signal_17555 ;
    wire new_AGEMA_signal_17556 ;
    wire new_AGEMA_signal_17557 ;
    wire new_AGEMA_signal_17558 ;
    wire new_AGEMA_signal_17559 ;
    wire new_AGEMA_signal_17560 ;
    wire new_AGEMA_signal_17561 ;
    wire new_AGEMA_signal_17562 ;
    wire new_AGEMA_signal_17563 ;
    wire new_AGEMA_signal_17564 ;
    wire new_AGEMA_signal_17565 ;
    wire new_AGEMA_signal_17566 ;
    wire new_AGEMA_signal_17567 ;
    wire new_AGEMA_signal_17568 ;
    wire new_AGEMA_signal_17569 ;
    wire new_AGEMA_signal_17570 ;
    wire new_AGEMA_signal_17571 ;
    wire new_AGEMA_signal_17572 ;
    wire new_AGEMA_signal_17573 ;
    wire new_AGEMA_signal_17574 ;
    wire new_AGEMA_signal_17575 ;
    wire new_AGEMA_signal_17576 ;
    wire new_AGEMA_signal_17577 ;
    wire new_AGEMA_signal_17578 ;
    wire new_AGEMA_signal_17579 ;
    wire new_AGEMA_signal_17580 ;
    wire new_AGEMA_signal_17581 ;
    wire new_AGEMA_signal_17582 ;
    wire new_AGEMA_signal_17583 ;
    wire new_AGEMA_signal_17584 ;
    wire new_AGEMA_signal_17585 ;
    wire new_AGEMA_signal_17586 ;
    wire new_AGEMA_signal_17587 ;
    wire new_AGEMA_signal_17588 ;
    wire new_AGEMA_signal_17589 ;
    wire new_AGEMA_signal_17590 ;
    wire new_AGEMA_signal_17591 ;
    wire new_AGEMA_signal_17592 ;
    wire new_AGEMA_signal_17593 ;
    wire new_AGEMA_signal_17594 ;
    wire new_AGEMA_signal_17595 ;
    wire new_AGEMA_signal_17596 ;
    wire new_AGEMA_signal_17597 ;
    wire new_AGEMA_signal_17598 ;
    wire new_AGEMA_signal_17599 ;
    wire new_AGEMA_signal_17600 ;
    wire new_AGEMA_signal_17601 ;
    wire new_AGEMA_signal_17602 ;
    wire new_AGEMA_signal_17603 ;
    wire new_AGEMA_signal_17604 ;
    wire new_AGEMA_signal_17605 ;
    wire new_AGEMA_signal_17606 ;
    wire new_AGEMA_signal_17607 ;
    wire new_AGEMA_signal_17608 ;
    wire new_AGEMA_signal_17609 ;
    wire new_AGEMA_signal_17610 ;
    wire new_AGEMA_signal_17611 ;
    wire new_AGEMA_signal_17612 ;
    wire new_AGEMA_signal_17613 ;
    wire new_AGEMA_signal_17614 ;
    wire new_AGEMA_signal_17615 ;
    wire new_AGEMA_signal_17616 ;
    wire new_AGEMA_signal_17617 ;
    wire new_AGEMA_signal_17618 ;
    wire new_AGEMA_signal_17619 ;
    wire new_AGEMA_signal_17620 ;
    wire new_AGEMA_signal_17621 ;
    wire new_AGEMA_signal_17622 ;
    wire new_AGEMA_signal_17623 ;
    wire new_AGEMA_signal_17624 ;
    wire new_AGEMA_signal_17625 ;
    wire new_AGEMA_signal_17626 ;
    wire new_AGEMA_signal_17627 ;
    wire new_AGEMA_signal_17628 ;
    wire new_AGEMA_signal_17629 ;
    wire new_AGEMA_signal_17630 ;
    wire new_AGEMA_signal_17631 ;
    wire new_AGEMA_signal_17632 ;
    wire new_AGEMA_signal_17633 ;
    wire new_AGEMA_signal_17634 ;
    wire new_AGEMA_signal_17635 ;
    wire new_AGEMA_signal_17636 ;
    wire new_AGEMA_signal_17637 ;
    wire new_AGEMA_signal_17638 ;
    wire new_AGEMA_signal_17639 ;
    wire new_AGEMA_signal_17640 ;
    wire new_AGEMA_signal_17641 ;
    wire new_AGEMA_signal_17642 ;
    wire new_AGEMA_signal_17643 ;
    wire new_AGEMA_signal_17644 ;
    wire new_AGEMA_signal_17645 ;
    wire new_AGEMA_signal_17646 ;
    wire new_AGEMA_signal_17647 ;
    wire new_AGEMA_signal_17648 ;
    wire new_AGEMA_signal_17649 ;
    wire new_AGEMA_signal_17650 ;
    wire new_AGEMA_signal_17651 ;
    wire new_AGEMA_signal_17652 ;
    wire new_AGEMA_signal_17653 ;
    wire new_AGEMA_signal_17654 ;
    wire new_AGEMA_signal_17655 ;
    wire new_AGEMA_signal_17656 ;
    wire new_AGEMA_signal_17657 ;
    wire new_AGEMA_signal_17658 ;
    wire new_AGEMA_signal_17659 ;
    wire new_AGEMA_signal_17660 ;
    wire new_AGEMA_signal_17661 ;
    wire new_AGEMA_signal_17662 ;
    wire new_AGEMA_signal_17663 ;
    wire new_AGEMA_signal_17664 ;
    wire new_AGEMA_signal_17665 ;
    wire new_AGEMA_signal_17666 ;
    wire new_AGEMA_signal_17667 ;
    wire new_AGEMA_signal_17668 ;
    wire new_AGEMA_signal_17669 ;
    wire new_AGEMA_signal_17670 ;
    wire new_AGEMA_signal_17671 ;
    wire new_AGEMA_signal_17672 ;
    wire new_AGEMA_signal_17673 ;
    wire new_AGEMA_signal_17674 ;
    wire new_AGEMA_signal_17675 ;
    wire new_AGEMA_signal_17676 ;
    wire new_AGEMA_signal_17677 ;
    wire new_AGEMA_signal_17678 ;
    wire new_AGEMA_signal_17679 ;
    wire new_AGEMA_signal_17680 ;
    wire new_AGEMA_signal_17681 ;
    wire new_AGEMA_signal_17682 ;
    wire new_AGEMA_signal_17683 ;
    wire new_AGEMA_signal_17684 ;
    wire new_AGEMA_signal_17685 ;
    wire new_AGEMA_signal_17686 ;
    wire new_AGEMA_signal_17687 ;
    wire new_AGEMA_signal_17688 ;
    wire new_AGEMA_signal_17689 ;
    wire new_AGEMA_signal_17690 ;
    wire new_AGEMA_signal_17691 ;
    wire new_AGEMA_signal_17692 ;
    wire new_AGEMA_signal_17693 ;
    wire new_AGEMA_signal_17694 ;
    wire new_AGEMA_signal_17695 ;
    wire new_AGEMA_signal_17696 ;
    wire new_AGEMA_signal_17697 ;
    wire new_AGEMA_signal_17698 ;
    wire new_AGEMA_signal_17699 ;
    wire new_AGEMA_signal_17700 ;
    wire new_AGEMA_signal_17701 ;
    wire new_AGEMA_signal_17702 ;
    wire new_AGEMA_signal_17703 ;
    wire new_AGEMA_signal_17704 ;
    wire new_AGEMA_signal_17705 ;
    wire new_AGEMA_signal_17706 ;
    wire new_AGEMA_signal_17707 ;
    wire new_AGEMA_signal_17708 ;
    wire new_AGEMA_signal_17709 ;
    wire new_AGEMA_signal_17710 ;
    wire new_AGEMA_signal_17711 ;
    wire new_AGEMA_signal_17712 ;
    wire new_AGEMA_signal_17713 ;
    wire new_AGEMA_signal_17714 ;
    wire new_AGEMA_signal_17715 ;
    wire new_AGEMA_signal_17716 ;
    wire new_AGEMA_signal_17717 ;
    wire new_AGEMA_signal_17718 ;
    wire new_AGEMA_signal_17719 ;
    wire new_AGEMA_signal_17720 ;
    wire new_AGEMA_signal_17721 ;
    wire new_AGEMA_signal_17722 ;
    wire new_AGEMA_signal_17723 ;
    wire new_AGEMA_signal_17724 ;
    wire new_AGEMA_signal_17725 ;
    wire new_AGEMA_signal_17726 ;
    wire new_AGEMA_signal_17727 ;
    wire new_AGEMA_signal_17728 ;
    wire new_AGEMA_signal_17729 ;

    /* cells in depth 0 */
    AND2_X1 U323 ( .A1 (n45), .A2 (n44), .ZN (AKSRnotDone) ) ;
    NOR2_X1 U324 ( .A1 (n60), .A2 (n49), .ZN (LastRoundorDone) ) ;
    AND2_X1 U325 ( .A1 (RoundCounter[0]), .A2 (LastRoundorDone), .ZN (done) ) ;
    INV_X1 U326 ( .A (RoundCounter[3]), .ZN (n60) ) ;
    NOR2_X1 U327 ( .A1 (InRoundCounter[0]), .A2 (InRoundCounter[1]), .ZN (n45) ) ;
    INV_X1 U328 ( .A (RoundCounter[2]), .ZN (n46) ) ;
    NAND2_X1 U329 ( .A1 (RoundCounter[1]), .A2 (n46), .ZN (n49) ) ;
    NOR2_X1 U330 ( .A1 (done), .A2 (InRoundCounter[2]), .ZN (n44) ) ;
    INV_X1 U331 ( .A (RoundCounter[1]), .ZN (n55) ) ;
    NAND2_X1 U332 ( .A1 (n55), .A2 (n46), .ZN (n47) ) ;
    NOR2_X1 U333 ( .A1 (RoundCounter[0]), .A2 (n47), .ZN (Rcon[0]) ) ;
    NOR2_X1 U334 ( .A1 (RoundCounter[0]), .A2 (RoundCounter[3]), .ZN (n58) ) ;
    NOR2_X1 U335 ( .A1 (n58), .A2 (n47), .ZN (Rcon[1]) ) ;
    NOR2_X1 U336 ( .A1 (RoundCounter[3]), .A2 (n49), .ZN (n48) ) ;
    NOR2_X1 U337 ( .A1 (n60), .A2 (n47), .ZN (n54) ) ;
    MUX2_X1 U338 ( .S (RoundCounter[0]), .A (n48), .B (n54), .Z (Rcon[2]) ) ;
    INV_X1 U339 ( .A (RoundCounter[0]), .ZN (n50) ) ;
    NOR2_X1 U340 ( .A1 (n50), .A2 (n49), .ZN (n51) ) ;
    MUX2_X1 U341 ( .S (RoundCounter[3]), .A (n51), .B (Rcon[0]), .Z (Rcon[3]) ) ;
    NAND2_X1 U342 ( .A1 (RoundCounter[2]), .A2 (n58), .ZN (n52) ) ;
    NOR2_X1 U343 ( .A1 (RoundCounter[1]), .A2 (n52), .ZN (n53) ) ;
    OR2_X1 U344 ( .A1 (n54), .A2 (n53), .ZN (Rcon[4]) ) ;
    XNOR2_X1 U345 ( .A (RoundCounter[2]), .B (RoundCounter[3]), .ZN (n57) ) ;
    NAND2_X1 U346 ( .A1 (RoundCounter[0]), .A2 (n55), .ZN (n56) ) ;
    NOR2_X1 U347 ( .A1 (n57), .A2 (n56), .ZN (Rcon[5]) ) ;
    INV_X1 U348 ( .A (n58), .ZN (n59) ) ;
    NAND2_X1 U349 ( .A1 (RoundCounter[1]), .A2 (RoundCounter[2]), .ZN (n61) ) ;
    NOR2_X1 U350 ( .A1 (n59), .A2 (n61), .ZN (Rcon[6]) ) ;
    NAND2_X1 U351 ( .A1 (RoundCounter[0]), .A2 (n60), .ZN (n62) ) ;
    NOR2_X1 U352 ( .A1 (n62), .A2 (n61), .ZN (Rcon[7]) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U353 ( .a ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, new_AGEMA_signal_2341, KSSubBytesInput[16]}), .c ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, new_AGEMA_signal_2344, ShiftRowsOutput[96]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U354 ( .a ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({new_AGEMA_signal_2352, new_AGEMA_signal_2351, new_AGEMA_signal_2350, RoundKey[100]}), .c ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, new_AGEMA_signal_2353, ShiftRowsOutput[68]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U355 ( .a ({ciphertext_s3[5], ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .b ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, new_AGEMA_signal_2359, RoundKey[101]}), .c ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, new_AGEMA_signal_2362, ShiftRowsOutput[69]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U356 ( .a ({ciphertext_s3[6], ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, new_AGEMA_signal_2368, RoundKey[102]}), .c ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, new_AGEMA_signal_2371, ShiftRowsOutput[70]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U357 ( .a ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, new_AGEMA_signal_2377, RoundKey[103]}), .c ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, new_AGEMA_signal_2380, ShiftRowsOutput[71]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U358 ( .a ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, new_AGEMA_signal_2386, RoundKey[104]}), .c ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, new_AGEMA_signal_2389, ShiftRowsOutput[40]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U359 ( .a ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .b ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, new_AGEMA_signal_2395, RoundKey[105]}), .c ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, new_AGEMA_signal_2398, ShiftRowsOutput[41]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U360 ( .a ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, new_AGEMA_signal_2404, RoundKey[106]}), .c ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, new_AGEMA_signal_2407, ShiftRowsOutput[42]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U361 ( .a ({ciphertext_s3[43], ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .b ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, new_AGEMA_signal_2413, RoundKey[107]}), .c ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, new_AGEMA_signal_2416, ShiftRowsOutput[43]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U362 ( .a ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, new_AGEMA_signal_2422, RoundKey[108]}), .c ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, new_AGEMA_signal_2425, ShiftRowsOutput[44]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U363 ( .a ({ciphertext_s3[45], ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .b ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, new_AGEMA_signal_2431, RoundKey[109]}), .c ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, new_AGEMA_signal_2434, ShiftRowsOutput[45]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U364 ( .a ({ciphertext_s3[74], ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .b ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, new_AGEMA_signal_2440, KSSubBytesInput[10]}), .c ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, new_AGEMA_signal_2443, ShiftRowsOutput[74]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U365 ( .a ({ciphertext_s3[46], ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, new_AGEMA_signal_2449, RoundKey[110]}), .c ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, new_AGEMA_signal_2452, ShiftRowsOutput[46]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U366 ( .a ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, new_AGEMA_signal_2458, RoundKey[111]}), .c ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, new_AGEMA_signal_2461, ShiftRowsOutput[47]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U367 ( .a ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, new_AGEMA_signal_2467, RoundKey[112]}), .c ({new_AGEMA_signal_2472, new_AGEMA_signal_2471, new_AGEMA_signal_2470, ShiftRowsOutput[16]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U368 ( .a ({ciphertext_s3[81], ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .b ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, new_AGEMA_signal_2476, RoundKey[113]}), .c ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, new_AGEMA_signal_2479, ShiftRowsOutput[17]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U369 ( .a ({ciphertext_s3[82], ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .b ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, new_AGEMA_signal_2485, RoundKey[114]}), .c ({new_AGEMA_signal_2490, new_AGEMA_signal_2489, new_AGEMA_signal_2488, ShiftRowsOutput[18]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U370 ( .a ({ciphertext_s3[83], ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}), .b ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, new_AGEMA_signal_2494, RoundKey[115]}), .c ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, new_AGEMA_signal_2497, ShiftRowsOutput[19]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U371 ( .a ({ciphertext_s3[84], ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .b ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, new_AGEMA_signal_2503, RoundKey[116]}), .c ({new_AGEMA_signal_2508, new_AGEMA_signal_2507, new_AGEMA_signal_2506, ShiftRowsOutput[20]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U372 ( .a ({ciphertext_s3[85], ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}), .b ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, new_AGEMA_signal_2512, RoundKey[117]}), .c ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, new_AGEMA_signal_2515, ShiftRowsOutput[21]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U373 ( .a ({ciphertext_s3[86], ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}), .b ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, new_AGEMA_signal_2521, RoundKey[118]}), .c ({new_AGEMA_signal_2526, new_AGEMA_signal_2525, new_AGEMA_signal_2524, ShiftRowsOutput[22]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U374 ( .a ({ciphertext_s3[87], ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .b ({new_AGEMA_signal_2532, new_AGEMA_signal_2531, new_AGEMA_signal_2530, RoundKey[119]}), .c ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, new_AGEMA_signal_2533, ShiftRowsOutput[23]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U375 ( .a ({ciphertext_s3[75], ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}), .b ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, new_AGEMA_signal_2539, KSSubBytesInput[11]}), .c ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, new_AGEMA_signal_2542, ShiftRowsOutput[75]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U376 ( .a ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_2550, new_AGEMA_signal_2549, new_AGEMA_signal_2548, RoundKey[120]}), .c ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, new_AGEMA_signal_2551, ShiftRowsOutput[120]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U377 ( .a ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, new_AGEMA_signal_2557, RoundKey[121]}), .c ({new_AGEMA_signal_2562, new_AGEMA_signal_2561, new_AGEMA_signal_2560, ShiftRowsOutput[121]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U378 ( .a ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .b ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, new_AGEMA_signal_2566, RoundKey[122]}), .c ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, new_AGEMA_signal_2569, ShiftRowsOutput[122]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U379 ( .a ({ciphertext_s3[123], ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .b ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, new_AGEMA_signal_2575, RoundKey[123]}), .c ({new_AGEMA_signal_2580, new_AGEMA_signal_2579, new_AGEMA_signal_2578, ShiftRowsOutput[123]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U380 ( .a ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, new_AGEMA_signal_2584, RoundKey[124]}), .c ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, new_AGEMA_signal_2587, ShiftRowsOutput[124]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U381 ( .a ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .b ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, new_AGEMA_signal_2593, RoundKey[125]}), .c ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, new_AGEMA_signal_2596, ShiftRowsOutput[125]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U382 ( .a ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .b ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, new_AGEMA_signal_2602, RoundKey[126]}), .c ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, new_AGEMA_signal_2605, ShiftRowsOutput[126]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U383 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, new_AGEMA_signal_2611, RoundKey[127]}), .c ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, new_AGEMA_signal_2614, ShiftRowsOutput[127]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U384 ( .a ({ciphertext_s3[76], ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .b ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, new_AGEMA_signal_2620, KSSubBytesInput[12]}), .c ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, new_AGEMA_signal_2623, ShiftRowsOutput[76]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U385 ( .a ({ciphertext_s3[77], ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}), .b ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, new_AGEMA_signal_2629, KSSubBytesInput[13]}), .c ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, new_AGEMA_signal_2632, ShiftRowsOutput[77]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U386 ( .a ({ciphertext_s3[78], ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}), .b ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, new_AGEMA_signal_2638, KSSubBytesInput[14]}), .c ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, new_AGEMA_signal_2641, ShiftRowsOutput[78]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U387 ( .a ({ciphertext_s3[79], ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .b ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, new_AGEMA_signal_2647, KSSubBytesInput[15]}), .c ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, new_AGEMA_signal_2650, ShiftRowsOutput[79]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U388 ( .a ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, new_AGEMA_signal_2656, KSSubBytesInput[0]}), .c ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, new_AGEMA_signal_2659, ShiftRowsOutput[48]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U389 ( .a ({ciphertext_s3[113], ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .b ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, new_AGEMA_signal_2665, KSSubBytesInput[1]}), .c ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, new_AGEMA_signal_2668, ShiftRowsOutput[49]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U390 ( .a ({ciphertext_s3[114], ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .b ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, new_AGEMA_signal_2674, KSSubBytesInput[2]}), .c ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, new_AGEMA_signal_2677, ShiftRowsOutput[50]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U391 ( .a ({ciphertext_s3[115], ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}), .b ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, new_AGEMA_signal_2683, KSSubBytesInput[3]}), .c ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, new_AGEMA_signal_2686, ShiftRowsOutput[51]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U392 ( .a ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .b ({new_AGEMA_signal_2694, new_AGEMA_signal_2693, new_AGEMA_signal_2692, KSSubBytesInput[17]}), .c ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, new_AGEMA_signal_2695, ShiftRowsOutput[97]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U393 ( .a ({ciphertext_s3[116], ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .b ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, new_AGEMA_signal_2701, KSSubBytesInput[4]}), .c ({new_AGEMA_signal_2706, new_AGEMA_signal_2705, new_AGEMA_signal_2704, ShiftRowsOutput[52]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U394 ( .a ({ciphertext_s3[117], ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}), .b ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, new_AGEMA_signal_2710, KSSubBytesInput[5]}), .c ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, new_AGEMA_signal_2713, ShiftRowsOutput[53]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U395 ( .a ({ciphertext_s3[118], ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}), .b ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, new_AGEMA_signal_2719, KSSubBytesInput[6]}), .c ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, new_AGEMA_signal_2722, ShiftRowsOutput[54]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U396 ( .a ({ciphertext_s3[119], ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .b ({new_AGEMA_signal_2730, new_AGEMA_signal_2729, new_AGEMA_signal_2728, KSSubBytesInput[7]}), .c ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, new_AGEMA_signal_2731, ShiftRowsOutput[55]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U397 ( .a ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, new_AGEMA_signal_2737, KSSubBytesInput[24]}), .c ({new_AGEMA_signal_2742, new_AGEMA_signal_2741, new_AGEMA_signal_2740, ShiftRowsOutput[24]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U398 ( .a ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, new_AGEMA_signal_2746, KSSubBytesInput[25]}), .c ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, new_AGEMA_signal_2749, ShiftRowsOutput[25]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U399 ( .a ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, new_AGEMA_signal_2755, KSSubBytesInput[26]}), .c ({new_AGEMA_signal_2760, new_AGEMA_signal_2759, new_AGEMA_signal_2758, ShiftRowsOutput[26]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U400 ( .a ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_2766, new_AGEMA_signal_2765, new_AGEMA_signal_2764, KSSubBytesInput[27]}), .c ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, new_AGEMA_signal_2767, ShiftRowsOutput[27]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U401 ( .a ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, new_AGEMA_signal_2773, KSSubBytesInput[28]}), .c ({new_AGEMA_signal_2778, new_AGEMA_signal_2777, new_AGEMA_signal_2776, ShiftRowsOutput[28]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U402 ( .a ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .b ({new_AGEMA_signal_2784, new_AGEMA_signal_2783, new_AGEMA_signal_2782, KSSubBytesInput[29]}), .c ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, new_AGEMA_signal_2785, ShiftRowsOutput[29]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U403 ( .a ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, new_AGEMA_signal_2791, KSSubBytesInput[18]}), .c ({new_AGEMA_signal_2796, new_AGEMA_signal_2795, new_AGEMA_signal_2794, ShiftRowsOutput[98]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U404 ( .a ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_2802, new_AGEMA_signal_2801, new_AGEMA_signal_2800, KSSubBytesInput[30]}), .c ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, new_AGEMA_signal_2803, ShiftRowsOutput[30]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U405 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, new_AGEMA_signal_2809, KSSubBytesInput[31]}), .c ({new_AGEMA_signal_2814, new_AGEMA_signal_2813, new_AGEMA_signal_2812, ShiftRowsOutput[31]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U406 ( .a ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_2820, new_AGEMA_signal_2819, new_AGEMA_signal_2818, RoundKey[32]}), .c ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, new_AGEMA_signal_2821, ShiftRowsOutput[0]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U407 ( .a ({ciphertext_s3[65], ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .b ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, new_AGEMA_signal_2827, RoundKey[33]}), .c ({new_AGEMA_signal_2832, new_AGEMA_signal_2831, new_AGEMA_signal_2830, ShiftRowsOutput[1]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U408 ( .a ({ciphertext_s3[66], ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .b ({new_AGEMA_signal_2838, new_AGEMA_signal_2837, new_AGEMA_signal_2836, RoundKey[34]}), .c ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, new_AGEMA_signal_2839, ShiftRowsOutput[2]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U409 ( .a ({ciphertext_s3[67], ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}), .b ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, new_AGEMA_signal_2845, RoundKey[35]}), .c ({new_AGEMA_signal_2850, new_AGEMA_signal_2849, new_AGEMA_signal_2848, ShiftRowsOutput[3]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U410 ( .a ({ciphertext_s3[68], ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .b ({new_AGEMA_signal_2856, new_AGEMA_signal_2855, new_AGEMA_signal_2854, RoundKey[36]}), .c ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, new_AGEMA_signal_2857, ShiftRowsOutput[4]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U411 ( .a ({ciphertext_s3[69], ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, new_AGEMA_signal_2863, RoundKey[37]}), .c ({new_AGEMA_signal_2868, new_AGEMA_signal_2867, new_AGEMA_signal_2866, ShiftRowsOutput[5]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U412 ( .a ({ciphertext_s3[70], ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}), .b ({new_AGEMA_signal_2874, new_AGEMA_signal_2873, new_AGEMA_signal_2872, RoundKey[38]}), .c ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, new_AGEMA_signal_2875, ShiftRowsOutput[6]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U413 ( .a ({ciphertext_s3[71], ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, new_AGEMA_signal_2881, RoundKey[39]}), .c ({new_AGEMA_signal_2886, new_AGEMA_signal_2885, new_AGEMA_signal_2884, ShiftRowsOutput[7]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U414 ( .a ({ciphertext_s3[35], ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .b ({new_AGEMA_signal_2892, new_AGEMA_signal_2891, new_AGEMA_signal_2890, KSSubBytesInput[19]}), .c ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, new_AGEMA_signal_2893, ShiftRowsOutput[99]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U415 ( .a ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, new_AGEMA_signal_2899, RoundKey[40]}), .c ({new_AGEMA_signal_2904, new_AGEMA_signal_2903, new_AGEMA_signal_2902, ShiftRowsOutput[104]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U416 ( .a ({ciphertext_s3[105], ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .b ({new_AGEMA_signal_2910, new_AGEMA_signal_2909, new_AGEMA_signal_2908, RoundKey[41]}), .c ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, new_AGEMA_signal_2911, ShiftRowsOutput[105]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U417 ( .a ({ciphertext_s3[106], ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .b ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, new_AGEMA_signal_2917, RoundKey[42]}), .c ({new_AGEMA_signal_2922, new_AGEMA_signal_2921, new_AGEMA_signal_2920, ShiftRowsOutput[106]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U418 ( .a ({ciphertext_s3[107], ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}), .b ({new_AGEMA_signal_2928, new_AGEMA_signal_2927, new_AGEMA_signal_2926, RoundKey[43]}), .c ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, new_AGEMA_signal_2929, ShiftRowsOutput[107]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U419 ( .a ({ciphertext_s3[108], ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .b ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, new_AGEMA_signal_2935, RoundKey[44]}), .c ({new_AGEMA_signal_2940, new_AGEMA_signal_2939, new_AGEMA_signal_2938, ShiftRowsOutput[108]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U420 ( .a ({ciphertext_s3[109], ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}), .b ({new_AGEMA_signal_2946, new_AGEMA_signal_2945, new_AGEMA_signal_2944, RoundKey[45]}), .c ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, new_AGEMA_signal_2947, ShiftRowsOutput[109]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U421 ( .a ({ciphertext_s3[110], ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}), .b ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, new_AGEMA_signal_2953, RoundKey[46]}), .c ({new_AGEMA_signal_2958, new_AGEMA_signal_2957, new_AGEMA_signal_2956, ShiftRowsOutput[110]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U422 ( .a ({ciphertext_s3[111], ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .b ({new_AGEMA_signal_2964, new_AGEMA_signal_2963, new_AGEMA_signal_2962, RoundKey[47]}), .c ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, new_AGEMA_signal_2965, ShiftRowsOutput[111]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U423 ( .a ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, new_AGEMA_signal_2971, RoundKey[48]}), .c ({new_AGEMA_signal_2976, new_AGEMA_signal_2975, new_AGEMA_signal_2974, ShiftRowsOutput[80]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U424 ( .a ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .b ({new_AGEMA_signal_2982, new_AGEMA_signal_2981, new_AGEMA_signal_2980, RoundKey[49]}), .c ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, new_AGEMA_signal_2983, ShiftRowsOutput[81]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U425 ( .a ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, new_AGEMA_signal_2989, KSSubBytesInput[20]}), .c ({new_AGEMA_signal_2994, new_AGEMA_signal_2993, new_AGEMA_signal_2992, ShiftRowsOutput[100]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U426 ( .a ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_3000, new_AGEMA_signal_2999, new_AGEMA_signal_2998, RoundKey[50]}), .c ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, new_AGEMA_signal_3001, ShiftRowsOutput[82]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U427 ( .a ({ciphertext_s3[19], ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .b ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, new_AGEMA_signal_3007, RoundKey[51]}), .c ({new_AGEMA_signal_3012, new_AGEMA_signal_3011, new_AGEMA_signal_3010, ShiftRowsOutput[83]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U428 ( .a ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({new_AGEMA_signal_3018, new_AGEMA_signal_3017, new_AGEMA_signal_3016, RoundKey[52]}), .c ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, new_AGEMA_signal_3019, ShiftRowsOutput[84]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U429 ( .a ({ciphertext_s3[21], ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .b ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, new_AGEMA_signal_3025, RoundKey[53]}), .c ({new_AGEMA_signal_3030, new_AGEMA_signal_3029, new_AGEMA_signal_3028, ShiftRowsOutput[85]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U430 ( .a ({ciphertext_s3[22], ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_3036, new_AGEMA_signal_3035, new_AGEMA_signal_3034, RoundKey[54]}), .c ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, new_AGEMA_signal_3037, ShiftRowsOutput[86]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U431 ( .a ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, new_AGEMA_signal_3043, RoundKey[55]}), .c ({new_AGEMA_signal_3048, new_AGEMA_signal_3047, new_AGEMA_signal_3046, ShiftRowsOutput[87]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U432 ( .a ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_3054, new_AGEMA_signal_3053, new_AGEMA_signal_3052, RoundKey[56]}), .c ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, new_AGEMA_signal_3055, ShiftRowsOutput[56]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U433 ( .a ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, new_AGEMA_signal_3061, RoundKey[57]}), .c ({new_AGEMA_signal_3066, new_AGEMA_signal_3065, new_AGEMA_signal_3064, ShiftRowsOutput[57]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U434 ( .a ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_3072, new_AGEMA_signal_3071, new_AGEMA_signal_3070, RoundKey[58]}), .c ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, new_AGEMA_signal_3073, ShiftRowsOutput[58]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U435 ( .a ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, new_AGEMA_signal_3079, RoundKey[59]}), .c ({new_AGEMA_signal_3084, new_AGEMA_signal_3083, new_AGEMA_signal_3082, ShiftRowsOutput[59]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U436 ( .a ({ciphertext_s3[37], ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .b ({new_AGEMA_signal_3090, new_AGEMA_signal_3089, new_AGEMA_signal_3088, KSSubBytesInput[21]}), .c ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, new_AGEMA_signal_3091, ShiftRowsOutput[101]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U437 ( .a ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, new_AGEMA_signal_3097, RoundKey[60]}), .c ({new_AGEMA_signal_3102, new_AGEMA_signal_3101, new_AGEMA_signal_3100, ShiftRowsOutput[60]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U438 ( .a ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .b ({new_AGEMA_signal_3108, new_AGEMA_signal_3107, new_AGEMA_signal_3106, RoundKey[61]}), .c ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, new_AGEMA_signal_3109, ShiftRowsOutput[61]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U439 ( .a ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, new_AGEMA_signal_3115, RoundKey[62]}), .c ({new_AGEMA_signal_3120, new_AGEMA_signal_3119, new_AGEMA_signal_3118, ShiftRowsOutput[62]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U440 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_3126, new_AGEMA_signal_3125, new_AGEMA_signal_3124, RoundKey[63]}), .c ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, new_AGEMA_signal_3127, ShiftRowsOutput[63]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U441 ( .a ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, new_AGEMA_signal_3133, RoundKey[64]}), .c ({new_AGEMA_signal_3138, new_AGEMA_signal_3137, new_AGEMA_signal_3136, ShiftRowsOutput[32]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U442 ( .a ({ciphertext_s3[97], ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .b ({new_AGEMA_signal_3144, new_AGEMA_signal_3143, new_AGEMA_signal_3142, RoundKey[65]}), .c ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, new_AGEMA_signal_3145, ShiftRowsOutput[33]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U443 ( .a ({ciphertext_s3[98], ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .b ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, new_AGEMA_signal_3151, RoundKey[66]}), .c ({new_AGEMA_signal_3156, new_AGEMA_signal_3155, new_AGEMA_signal_3154, ShiftRowsOutput[34]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U444 ( .a ({ciphertext_s3[99], ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}), .b ({new_AGEMA_signal_3162, new_AGEMA_signal_3161, new_AGEMA_signal_3160, RoundKey[67]}), .c ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, new_AGEMA_signal_3163, ShiftRowsOutput[35]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U445 ( .a ({ciphertext_s3[100], ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .b ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, new_AGEMA_signal_3169, RoundKey[68]}), .c ({new_AGEMA_signal_3174, new_AGEMA_signal_3173, new_AGEMA_signal_3172, ShiftRowsOutput[36]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U446 ( .a ({ciphertext_s3[101], ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}), .b ({new_AGEMA_signal_3180, new_AGEMA_signal_3179, new_AGEMA_signal_3178, RoundKey[69]}), .c ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, new_AGEMA_signal_3181, ShiftRowsOutput[37]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U447 ( .a ({ciphertext_s3[38], ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, new_AGEMA_signal_3187, KSSubBytesInput[22]}), .c ({new_AGEMA_signal_3192, new_AGEMA_signal_3191, new_AGEMA_signal_3190, ShiftRowsOutput[102]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U448 ( .a ({ciphertext_s3[102], ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}), .b ({new_AGEMA_signal_3198, new_AGEMA_signal_3197, new_AGEMA_signal_3196, RoundKey[70]}), .c ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, new_AGEMA_signal_3199, ShiftRowsOutput[38]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U449 ( .a ({ciphertext_s3[103], ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .b ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, new_AGEMA_signal_3205, RoundKey[71]}), .c ({new_AGEMA_signal_3210, new_AGEMA_signal_3209, new_AGEMA_signal_3208, ShiftRowsOutput[39]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U450 ( .a ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_3216, new_AGEMA_signal_3215, new_AGEMA_signal_3214, RoundKey[72]}), .c ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, new_AGEMA_signal_3217, ShiftRowsOutput[8]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U451 ( .a ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .b ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, new_AGEMA_signal_3223, RoundKey[73]}), .c ({new_AGEMA_signal_3228, new_AGEMA_signal_3227, new_AGEMA_signal_3226, ShiftRowsOutput[9]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U452 ( .a ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_3234, new_AGEMA_signal_3233, new_AGEMA_signal_3232, RoundKey[74]}), .c ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, new_AGEMA_signal_3235, ShiftRowsOutput[10]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U453 ( .a ({ciphertext_s3[11], ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .b ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, new_AGEMA_signal_3241, RoundKey[75]}), .c ({new_AGEMA_signal_3246, new_AGEMA_signal_3245, new_AGEMA_signal_3244, ShiftRowsOutput[11]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U454 ( .a ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({new_AGEMA_signal_3252, new_AGEMA_signal_3251, new_AGEMA_signal_3250, RoundKey[76]}), .c ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, new_AGEMA_signal_3253, ShiftRowsOutput[12]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U455 ( .a ({ciphertext_s3[13], ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .b ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, new_AGEMA_signal_3259, RoundKey[77]}), .c ({new_AGEMA_signal_3264, new_AGEMA_signal_3263, new_AGEMA_signal_3262, ShiftRowsOutput[13]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U456 ( .a ({ciphertext_s3[14], ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_3270, new_AGEMA_signal_3269, new_AGEMA_signal_3268, RoundKey[78]}), .c ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, new_AGEMA_signal_3271, ShiftRowsOutput[14]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U457 ( .a ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, new_AGEMA_signal_3277, RoundKey[79]}), .c ({new_AGEMA_signal_3282, new_AGEMA_signal_3281, new_AGEMA_signal_3280, ShiftRowsOutput[15]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U458 ( .a ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({new_AGEMA_signal_3288, new_AGEMA_signal_3287, new_AGEMA_signal_3286, KSSubBytesInput[23]}), .c ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, new_AGEMA_signal_3289, ShiftRowsOutput[103]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U459 ( .a ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, new_AGEMA_signal_3295, RoundKey[80]}), .c ({new_AGEMA_signal_3300, new_AGEMA_signal_3299, new_AGEMA_signal_3298, ShiftRowsOutput[112]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U460 ( .a ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .b ({new_AGEMA_signal_3306, new_AGEMA_signal_3305, new_AGEMA_signal_3304, RoundKey[81]}), .c ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, new_AGEMA_signal_3307, ShiftRowsOutput[113]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U461 ( .a ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, new_AGEMA_signal_3313, RoundKey[82]}), .c ({new_AGEMA_signal_3318, new_AGEMA_signal_3317, new_AGEMA_signal_3316, ShiftRowsOutput[114]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U462 ( .a ({ciphertext_s3[51], ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .b ({new_AGEMA_signal_3324, new_AGEMA_signal_3323, new_AGEMA_signal_3322, RoundKey[83]}), .c ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, new_AGEMA_signal_3325, ShiftRowsOutput[115]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U463 ( .a ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, new_AGEMA_signal_3331, RoundKey[84]}), .c ({new_AGEMA_signal_3336, new_AGEMA_signal_3335, new_AGEMA_signal_3334, ShiftRowsOutput[116]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U464 ( .a ({ciphertext_s3[53], ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .b ({new_AGEMA_signal_3342, new_AGEMA_signal_3341, new_AGEMA_signal_3340, RoundKey[85]}), .c ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, new_AGEMA_signal_3343, ShiftRowsOutput[117]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U465 ( .a ({ciphertext_s3[54], ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, new_AGEMA_signal_3349, RoundKey[86]}), .c ({new_AGEMA_signal_3354, new_AGEMA_signal_3353, new_AGEMA_signal_3352, ShiftRowsOutput[118]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U466 ( .a ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({new_AGEMA_signal_3360, new_AGEMA_signal_3359, new_AGEMA_signal_3358, RoundKey[87]}), .c ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, new_AGEMA_signal_3361, ShiftRowsOutput[119]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U467 ( .a ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, new_AGEMA_signal_3367, RoundKey[88]}), .c ({new_AGEMA_signal_3372, new_AGEMA_signal_3371, new_AGEMA_signal_3370, ShiftRowsOutput[88]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U468 ( .a ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .b ({new_AGEMA_signal_3378, new_AGEMA_signal_3377, new_AGEMA_signal_3376, RoundKey[89]}), .c ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, new_AGEMA_signal_3379, ShiftRowsOutput[89]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U469 ( .a ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, new_AGEMA_signal_3385, KSSubBytesInput[8]}), .c ({new_AGEMA_signal_3390, new_AGEMA_signal_3389, new_AGEMA_signal_3388, ShiftRowsOutput[72]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U470 ( .a ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .b ({new_AGEMA_signal_3396, new_AGEMA_signal_3395, new_AGEMA_signal_3394, RoundKey[90]}), .c ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, new_AGEMA_signal_3397, ShiftRowsOutput[90]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U471 ( .a ({ciphertext_s3[91], ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .b ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, new_AGEMA_signal_3403, RoundKey[91]}), .c ({new_AGEMA_signal_3408, new_AGEMA_signal_3407, new_AGEMA_signal_3406, ShiftRowsOutput[91]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U472 ( .a ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .b ({new_AGEMA_signal_3414, new_AGEMA_signal_3413, new_AGEMA_signal_3412, RoundKey[92]}), .c ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, new_AGEMA_signal_3415, ShiftRowsOutput[92]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U473 ( .a ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .b ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, new_AGEMA_signal_3421, RoundKey[93]}), .c ({new_AGEMA_signal_3426, new_AGEMA_signal_3425, new_AGEMA_signal_3424, ShiftRowsOutput[93]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U474 ( .a ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .b ({new_AGEMA_signal_3432, new_AGEMA_signal_3431, new_AGEMA_signal_3430, RoundKey[94]}), .c ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, new_AGEMA_signal_3433, ShiftRowsOutput[94]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U475 ( .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, new_AGEMA_signal_3439, RoundKey[95]}), .c ({new_AGEMA_signal_3444, new_AGEMA_signal_3443, new_AGEMA_signal_3442, ShiftRowsOutput[95]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U476 ( .a ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_3450, new_AGEMA_signal_3449, new_AGEMA_signal_3448, RoundKey[96]}), .c ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, new_AGEMA_signal_3451, ShiftRowsOutput[64]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U477 ( .a ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .b ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, new_AGEMA_signal_3457, RoundKey[97]}), .c ({new_AGEMA_signal_3462, new_AGEMA_signal_3461, new_AGEMA_signal_3460, ShiftRowsOutput[65]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U478 ( .a ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_3468, new_AGEMA_signal_3467, new_AGEMA_signal_3466, RoundKey[98]}), .c ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, new_AGEMA_signal_3469, ShiftRowsOutput[66]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U479 ( .a ({ciphertext_s3[3], ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .b ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, new_AGEMA_signal_3475, RoundKey[99]}), .c ({new_AGEMA_signal_3480, new_AGEMA_signal_3479, new_AGEMA_signal_3478, ShiftRowsOutput[67]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) U480 ( .a ({ciphertext_s3[73], ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .b ({new_AGEMA_signal_3486, new_AGEMA_signal_3485, new_AGEMA_signal_3484, KSSubBytesInput[9]}), .c ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, new_AGEMA_signal_3487, ShiftRowsOutput[73]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3588, new_AGEMA_signal_3587, new_AGEMA_signal_3586, RoundOutput[32]}), .a ({plaintext_s3[32], plaintext_s2[32], plaintext_s1[32], plaintext_s0[32]}), .c ({new_AGEMA_signal_3879, new_AGEMA_signal_3878, new_AGEMA_signal_3877, RoundReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, new_AGEMA_signal_3589, RoundOutput[33]}), .a ({plaintext_s3[33], plaintext_s2[33], plaintext_s1[33], plaintext_s0[33]}), .c ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, new_AGEMA_signal_3883, RoundReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3594, new_AGEMA_signal_3593, new_AGEMA_signal_3592, RoundOutput[34]}), .a ({plaintext_s3[34], plaintext_s2[34], plaintext_s1[34], plaintext_s0[34]}), .c ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, new_AGEMA_signal_3889, RoundReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, new_AGEMA_signal_3595, RoundOutput[35]}), .a ({plaintext_s3[35], plaintext_s2[35], plaintext_s1[35], plaintext_s0[35]}), .c ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, new_AGEMA_signal_3895, RoundReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3600, new_AGEMA_signal_3599, new_AGEMA_signal_3598, RoundOutput[36]}), .a ({plaintext_s3[36], plaintext_s2[36], plaintext_s1[36], plaintext_s0[36]}), .c ({new_AGEMA_signal_3903, new_AGEMA_signal_3902, new_AGEMA_signal_3901, RoundReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, new_AGEMA_signal_3601, RoundOutput[37]}), .a ({plaintext_s3[37], plaintext_s2[37], plaintext_s1[37], plaintext_s0[37]}), .c ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, new_AGEMA_signal_3907, RoundReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3606, new_AGEMA_signal_3605, new_AGEMA_signal_3604, RoundOutput[38]}), .a ({plaintext_s3[38], plaintext_s2[38], plaintext_s1[38], plaintext_s0[38]}), .c ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, new_AGEMA_signal_3913, RoundReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, new_AGEMA_signal_3607, RoundOutput[39]}), .a ({plaintext_s3[39], plaintext_s2[39], plaintext_s1[39], plaintext_s0[39]}), .c ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, new_AGEMA_signal_3919, RoundReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3612, new_AGEMA_signal_3611, new_AGEMA_signal_3610, RoundOutput[40]}), .a ({plaintext_s3[40], plaintext_s2[40], plaintext_s1[40], plaintext_s0[40]}), .c ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, new_AGEMA_signal_3925, RoundReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, new_AGEMA_signal_3613, RoundOutput[41]}), .a ({plaintext_s3[41], plaintext_s2[41], plaintext_s1[41], plaintext_s0[41]}), .c ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, new_AGEMA_signal_3931, RoundReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3618, new_AGEMA_signal_3617, new_AGEMA_signal_3616, RoundOutput[42]}), .a ({plaintext_s3[42], plaintext_s2[42], plaintext_s1[42], plaintext_s0[42]}), .c ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, new_AGEMA_signal_3937, RoundReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, new_AGEMA_signal_3619, RoundOutput[43]}), .a ({plaintext_s3[43], plaintext_s2[43], plaintext_s1[43], plaintext_s0[43]}), .c ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, new_AGEMA_signal_3943, RoundReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3624, new_AGEMA_signal_3623, new_AGEMA_signal_3622, RoundOutput[44]}), .a ({plaintext_s3[44], plaintext_s2[44], plaintext_s1[44], plaintext_s0[44]}), .c ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, new_AGEMA_signal_3949, RoundReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, new_AGEMA_signal_3625, RoundOutput[45]}), .a ({plaintext_s3[45], plaintext_s2[45], plaintext_s1[45], plaintext_s0[45]}), .c ({new_AGEMA_signal_3957, new_AGEMA_signal_3956, new_AGEMA_signal_3955, RoundReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3630, new_AGEMA_signal_3629, new_AGEMA_signal_3628, RoundOutput[46]}), .a ({plaintext_s3[46], plaintext_s2[46], plaintext_s1[46], plaintext_s0[46]}), .c ({new_AGEMA_signal_3963, new_AGEMA_signal_3962, new_AGEMA_signal_3961, RoundReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, new_AGEMA_signal_3631, RoundOutput[47]}), .a ({plaintext_s3[47], plaintext_s2[47], plaintext_s1[47], plaintext_s0[47]}), .c ({new_AGEMA_signal_3969, new_AGEMA_signal_3968, new_AGEMA_signal_3967, RoundReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3636, new_AGEMA_signal_3635, new_AGEMA_signal_3634, RoundOutput[48]}), .a ({plaintext_s3[48], plaintext_s2[48], plaintext_s1[48], plaintext_s0[48]}), .c ({new_AGEMA_signal_3975, new_AGEMA_signal_3974, new_AGEMA_signal_3973, RoundReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, new_AGEMA_signal_3637, RoundOutput[49]}), .a ({plaintext_s3[49], plaintext_s2[49], plaintext_s1[49], plaintext_s0[49]}), .c ({new_AGEMA_signal_3981, new_AGEMA_signal_3980, new_AGEMA_signal_3979, RoundReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3642, new_AGEMA_signal_3641, new_AGEMA_signal_3640, RoundOutput[50]}), .a ({plaintext_s3[50], plaintext_s2[50], plaintext_s1[50], plaintext_s0[50]}), .c ({new_AGEMA_signal_3987, new_AGEMA_signal_3986, new_AGEMA_signal_3985, RoundReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, new_AGEMA_signal_3643, RoundOutput[51]}), .a ({plaintext_s3[51], plaintext_s2[51], plaintext_s1[51], plaintext_s0[51]}), .c ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, new_AGEMA_signal_3991, RoundReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3648, new_AGEMA_signal_3647, new_AGEMA_signal_3646, RoundOutput[52]}), .a ({plaintext_s3[52], plaintext_s2[52], plaintext_s1[52], plaintext_s0[52]}), .c ({new_AGEMA_signal_3999, new_AGEMA_signal_3998, new_AGEMA_signal_3997, RoundReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, new_AGEMA_signal_3649, RoundOutput[53]}), .a ({plaintext_s3[53], plaintext_s2[53], plaintext_s1[53], plaintext_s0[53]}), .c ({new_AGEMA_signal_4005, new_AGEMA_signal_4004, new_AGEMA_signal_4003, RoundReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3654, new_AGEMA_signal_3653, new_AGEMA_signal_3652, RoundOutput[54]}), .a ({plaintext_s3[54], plaintext_s2[54], plaintext_s1[54], plaintext_s0[54]}), .c ({new_AGEMA_signal_4011, new_AGEMA_signal_4010, new_AGEMA_signal_4009, RoundReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, new_AGEMA_signal_3655, RoundOutput[55]}), .a ({plaintext_s3[55], plaintext_s2[55], plaintext_s1[55], plaintext_s0[55]}), .c ({new_AGEMA_signal_4017, new_AGEMA_signal_4016, new_AGEMA_signal_4015, RoundReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3660, new_AGEMA_signal_3659, new_AGEMA_signal_3658, RoundOutput[56]}), .a ({plaintext_s3[56], plaintext_s2[56], plaintext_s1[56], plaintext_s0[56]}), .c ({new_AGEMA_signal_4023, new_AGEMA_signal_4022, new_AGEMA_signal_4021, RoundReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, new_AGEMA_signal_3661, RoundOutput[57]}), .a ({plaintext_s3[57], plaintext_s2[57], plaintext_s1[57], plaintext_s0[57]}), .c ({new_AGEMA_signal_4029, new_AGEMA_signal_4028, new_AGEMA_signal_4027, RoundReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3666, new_AGEMA_signal_3665, new_AGEMA_signal_3664, RoundOutput[58]}), .a ({plaintext_s3[58], plaintext_s2[58], plaintext_s1[58], plaintext_s0[58]}), .c ({new_AGEMA_signal_4035, new_AGEMA_signal_4034, new_AGEMA_signal_4033, RoundReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, new_AGEMA_signal_3667, RoundOutput[59]}), .a ({plaintext_s3[59], plaintext_s2[59], plaintext_s1[59], plaintext_s0[59]}), .c ({new_AGEMA_signal_4041, new_AGEMA_signal_4040, new_AGEMA_signal_4039, RoundReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3672, new_AGEMA_signal_3671, new_AGEMA_signal_3670, RoundOutput[60]}), .a ({plaintext_s3[60], plaintext_s2[60], plaintext_s1[60], plaintext_s0[60]}), .c ({new_AGEMA_signal_4047, new_AGEMA_signal_4046, new_AGEMA_signal_4045, RoundReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, new_AGEMA_signal_3673, RoundOutput[61]}), .a ({plaintext_s3[61], plaintext_s2[61], plaintext_s1[61], plaintext_s0[61]}), .c ({new_AGEMA_signal_4053, new_AGEMA_signal_4052, new_AGEMA_signal_4051, RoundReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3678, new_AGEMA_signal_3677, new_AGEMA_signal_3676, RoundOutput[62]}), .a ({plaintext_s3[62], plaintext_s2[62], plaintext_s1[62], plaintext_s0[62]}), .c ({new_AGEMA_signal_4059, new_AGEMA_signal_4058, new_AGEMA_signal_4057, RoundReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, new_AGEMA_signal_3679, RoundOutput[63]}), .a ({plaintext_s3[63], plaintext_s2[63], plaintext_s1[63], plaintext_s0[63]}), .c ({new_AGEMA_signal_4065, new_AGEMA_signal_4064, new_AGEMA_signal_4063, RoundReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3684, new_AGEMA_signal_3683, new_AGEMA_signal_3682, RoundOutput[64]}), .a ({plaintext_s3[64], plaintext_s2[64], plaintext_s1[64], plaintext_s0[64]}), .c ({new_AGEMA_signal_4071, new_AGEMA_signal_4070, new_AGEMA_signal_4069, RoundReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, new_AGEMA_signal_3685, RoundOutput[65]}), .a ({plaintext_s3[65], plaintext_s2[65], plaintext_s1[65], plaintext_s0[65]}), .c ({new_AGEMA_signal_4077, new_AGEMA_signal_4076, new_AGEMA_signal_4075, RoundReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3690, new_AGEMA_signal_3689, new_AGEMA_signal_3688, RoundOutput[66]}), .a ({plaintext_s3[66], plaintext_s2[66], plaintext_s1[66], plaintext_s0[66]}), .c ({new_AGEMA_signal_4083, new_AGEMA_signal_4082, new_AGEMA_signal_4081, RoundReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, new_AGEMA_signal_3691, RoundOutput[67]}), .a ({plaintext_s3[67], plaintext_s2[67], plaintext_s1[67], plaintext_s0[67]}), .c ({new_AGEMA_signal_4089, new_AGEMA_signal_4088, new_AGEMA_signal_4087, RoundReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3696, new_AGEMA_signal_3695, new_AGEMA_signal_3694, RoundOutput[68]}), .a ({plaintext_s3[68], plaintext_s2[68], plaintext_s1[68], plaintext_s0[68]}), .c ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, new_AGEMA_signal_4093, RoundReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, new_AGEMA_signal_3697, RoundOutput[69]}), .a ({plaintext_s3[69], plaintext_s2[69], plaintext_s1[69], plaintext_s0[69]}), .c ({new_AGEMA_signal_4101, new_AGEMA_signal_4100, new_AGEMA_signal_4099, RoundReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3702, new_AGEMA_signal_3701, new_AGEMA_signal_3700, RoundOutput[70]}), .a ({plaintext_s3[70], plaintext_s2[70], plaintext_s1[70], plaintext_s0[70]}), .c ({new_AGEMA_signal_4107, new_AGEMA_signal_4106, new_AGEMA_signal_4105, RoundReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, new_AGEMA_signal_3703, RoundOutput[71]}), .a ({plaintext_s3[71], plaintext_s2[71], plaintext_s1[71], plaintext_s0[71]}), .c ({new_AGEMA_signal_4113, new_AGEMA_signal_4112, new_AGEMA_signal_4111, RoundReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3708, new_AGEMA_signal_3707, new_AGEMA_signal_3706, RoundOutput[72]}), .a ({plaintext_s3[72], plaintext_s2[72], plaintext_s1[72], plaintext_s0[72]}), .c ({new_AGEMA_signal_4119, new_AGEMA_signal_4118, new_AGEMA_signal_4117, RoundReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, new_AGEMA_signal_3709, RoundOutput[73]}), .a ({plaintext_s3[73], plaintext_s2[73], plaintext_s1[73], plaintext_s0[73]}), .c ({new_AGEMA_signal_4125, new_AGEMA_signal_4124, new_AGEMA_signal_4123, RoundReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3714, new_AGEMA_signal_3713, new_AGEMA_signal_3712, RoundOutput[74]}), .a ({plaintext_s3[74], plaintext_s2[74], plaintext_s1[74], plaintext_s0[74]}), .c ({new_AGEMA_signal_4131, new_AGEMA_signal_4130, new_AGEMA_signal_4129, RoundReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, new_AGEMA_signal_3715, RoundOutput[75]}), .a ({plaintext_s3[75], plaintext_s2[75], plaintext_s1[75], plaintext_s0[75]}), .c ({new_AGEMA_signal_4137, new_AGEMA_signal_4136, new_AGEMA_signal_4135, RoundReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3720, new_AGEMA_signal_3719, new_AGEMA_signal_3718, RoundOutput[76]}), .a ({plaintext_s3[76], plaintext_s2[76], plaintext_s1[76], plaintext_s0[76]}), .c ({new_AGEMA_signal_4143, new_AGEMA_signal_4142, new_AGEMA_signal_4141, RoundReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3723, new_AGEMA_signal_3722, new_AGEMA_signal_3721, RoundOutput[77]}), .a ({plaintext_s3[77], plaintext_s2[77], plaintext_s1[77], plaintext_s0[77]}), .c ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, new_AGEMA_signal_4147, RoundReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3726, new_AGEMA_signal_3725, new_AGEMA_signal_3724, RoundOutput[78]}), .a ({plaintext_s3[78], plaintext_s2[78], plaintext_s1[78], plaintext_s0[78]}), .c ({new_AGEMA_signal_4155, new_AGEMA_signal_4154, new_AGEMA_signal_4153, RoundReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3729, new_AGEMA_signal_3728, new_AGEMA_signal_3727, RoundOutput[79]}), .a ({plaintext_s3[79], plaintext_s2[79], plaintext_s1[79], plaintext_s0[79]}), .c ({new_AGEMA_signal_4161, new_AGEMA_signal_4160, new_AGEMA_signal_4159, RoundReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3732, new_AGEMA_signal_3731, new_AGEMA_signal_3730, RoundOutput[80]}), .a ({plaintext_s3[80], plaintext_s2[80], plaintext_s1[80], plaintext_s0[80]}), .c ({new_AGEMA_signal_4167, new_AGEMA_signal_4166, new_AGEMA_signal_4165, RoundReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3735, new_AGEMA_signal_3734, new_AGEMA_signal_3733, RoundOutput[81]}), .a ({plaintext_s3[81], plaintext_s2[81], plaintext_s1[81], plaintext_s0[81]}), .c ({new_AGEMA_signal_4173, new_AGEMA_signal_4172, new_AGEMA_signal_4171, RoundReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3738, new_AGEMA_signal_3737, new_AGEMA_signal_3736, RoundOutput[82]}), .a ({plaintext_s3[82], plaintext_s2[82], plaintext_s1[82], plaintext_s0[82]}), .c ({new_AGEMA_signal_4179, new_AGEMA_signal_4178, new_AGEMA_signal_4177, RoundReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3741, new_AGEMA_signal_3740, new_AGEMA_signal_3739, RoundOutput[83]}), .a ({plaintext_s3[83], plaintext_s2[83], plaintext_s1[83], plaintext_s0[83]}), .c ({new_AGEMA_signal_4185, new_AGEMA_signal_4184, new_AGEMA_signal_4183, RoundReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3744, new_AGEMA_signal_3743, new_AGEMA_signal_3742, RoundOutput[84]}), .a ({plaintext_s3[84], plaintext_s2[84], plaintext_s1[84], plaintext_s0[84]}), .c ({new_AGEMA_signal_4191, new_AGEMA_signal_4190, new_AGEMA_signal_4189, RoundReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, new_AGEMA_signal_3745, RoundOutput[85]}), .a ({plaintext_s3[85], plaintext_s2[85], plaintext_s1[85], plaintext_s0[85]}), .c ({new_AGEMA_signal_4197, new_AGEMA_signal_4196, new_AGEMA_signal_4195, RoundReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3750, new_AGEMA_signal_3749, new_AGEMA_signal_3748, RoundOutput[86]}), .a ({plaintext_s3[86], plaintext_s2[86], plaintext_s1[86], plaintext_s0[86]}), .c ({new_AGEMA_signal_4203, new_AGEMA_signal_4202, new_AGEMA_signal_4201, RoundReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, new_AGEMA_signal_3751, RoundOutput[87]}), .a ({plaintext_s3[87], plaintext_s2[87], plaintext_s1[87], plaintext_s0[87]}), .c ({new_AGEMA_signal_4209, new_AGEMA_signal_4208, new_AGEMA_signal_4207, RoundReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3756, new_AGEMA_signal_3755, new_AGEMA_signal_3754, RoundOutput[88]}), .a ({plaintext_s3[88], plaintext_s2[88], plaintext_s1[88], plaintext_s0[88]}), .c ({new_AGEMA_signal_4215, new_AGEMA_signal_4214, new_AGEMA_signal_4213, RoundReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, new_AGEMA_signal_3757, RoundOutput[89]}), .a ({plaintext_s3[89], plaintext_s2[89], plaintext_s1[89], plaintext_s0[89]}), .c ({new_AGEMA_signal_4221, new_AGEMA_signal_4220, new_AGEMA_signal_4219, RoundReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3762, new_AGEMA_signal_3761, new_AGEMA_signal_3760, RoundOutput[90]}), .a ({plaintext_s3[90], plaintext_s2[90], plaintext_s1[90], plaintext_s0[90]}), .c ({new_AGEMA_signal_4227, new_AGEMA_signal_4226, new_AGEMA_signal_4225, RoundReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, new_AGEMA_signal_3763, RoundOutput[91]}), .a ({plaintext_s3[91], plaintext_s2[91], plaintext_s1[91], plaintext_s0[91]}), .c ({new_AGEMA_signal_4233, new_AGEMA_signal_4232, new_AGEMA_signal_4231, RoundReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3768, new_AGEMA_signal_3767, new_AGEMA_signal_3766, RoundOutput[92]}), .a ({plaintext_s3[92], plaintext_s2[92], plaintext_s1[92], plaintext_s0[92]}), .c ({new_AGEMA_signal_4239, new_AGEMA_signal_4238, new_AGEMA_signal_4237, RoundReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, new_AGEMA_signal_3769, RoundOutput[93]}), .a ({plaintext_s3[93], plaintext_s2[93], plaintext_s1[93], plaintext_s0[93]}), .c ({new_AGEMA_signal_4245, new_AGEMA_signal_4244, new_AGEMA_signal_4243, RoundReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3774, new_AGEMA_signal_3773, new_AGEMA_signal_3772, RoundOutput[94]}), .a ({plaintext_s3[94], plaintext_s2[94], plaintext_s1[94], plaintext_s0[94]}), .c ({new_AGEMA_signal_4251, new_AGEMA_signal_4250, new_AGEMA_signal_4249, RoundReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, new_AGEMA_signal_3775, RoundOutput[95]}), .a ({plaintext_s3[95], plaintext_s2[95], plaintext_s1[95], plaintext_s0[95]}), .c ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, new_AGEMA_signal_4255, RoundReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3780, new_AGEMA_signal_3779, new_AGEMA_signal_3778, RoundOutput[96]}), .a ({plaintext_s3[96], plaintext_s2[96], plaintext_s1[96], plaintext_s0[96]}), .c ({new_AGEMA_signal_4263, new_AGEMA_signal_4262, new_AGEMA_signal_4261, RoundReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, new_AGEMA_signal_3781, RoundOutput[97]}), .a ({plaintext_s3[97], plaintext_s2[97], plaintext_s1[97], plaintext_s0[97]}), .c ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, new_AGEMA_signal_4267, RoundReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3786, new_AGEMA_signal_3785, new_AGEMA_signal_3784, RoundOutput[98]}), .a ({plaintext_s3[98], plaintext_s2[98], plaintext_s1[98], plaintext_s0[98]}), .c ({new_AGEMA_signal_4275, new_AGEMA_signal_4274, new_AGEMA_signal_4273, RoundReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, new_AGEMA_signal_3787, RoundOutput[99]}), .a ({plaintext_s3[99], plaintext_s2[99], plaintext_s1[99], plaintext_s0[99]}), .c ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, new_AGEMA_signal_4279, RoundReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3792, new_AGEMA_signal_3791, new_AGEMA_signal_3790, RoundOutput[100]}), .a ({plaintext_s3[100], plaintext_s2[100], plaintext_s1[100], plaintext_s0[100]}), .c ({new_AGEMA_signal_4287, new_AGEMA_signal_4286, new_AGEMA_signal_4285, RoundReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, new_AGEMA_signal_3793, RoundOutput[101]}), .a ({plaintext_s3[101], plaintext_s2[101], plaintext_s1[101], plaintext_s0[101]}), .c ({new_AGEMA_signal_4293, new_AGEMA_signal_4292, new_AGEMA_signal_4291, RoundReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3798, new_AGEMA_signal_3797, new_AGEMA_signal_3796, RoundOutput[102]}), .a ({plaintext_s3[102], plaintext_s2[102], plaintext_s1[102], plaintext_s0[102]}), .c ({new_AGEMA_signal_4299, new_AGEMA_signal_4298, new_AGEMA_signal_4297, RoundReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, new_AGEMA_signal_3799, RoundOutput[103]}), .a ({plaintext_s3[103], plaintext_s2[103], plaintext_s1[103], plaintext_s0[103]}), .c ({new_AGEMA_signal_4305, new_AGEMA_signal_4304, new_AGEMA_signal_4303, RoundReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3804, new_AGEMA_signal_3803, new_AGEMA_signal_3802, RoundOutput[104]}), .a ({plaintext_s3[104], plaintext_s2[104], plaintext_s1[104], plaintext_s0[104]}), .c ({new_AGEMA_signal_4311, new_AGEMA_signal_4310, new_AGEMA_signal_4309, RoundReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, new_AGEMA_signal_3805, RoundOutput[105]}), .a ({plaintext_s3[105], plaintext_s2[105], plaintext_s1[105], plaintext_s0[105]}), .c ({new_AGEMA_signal_4317, new_AGEMA_signal_4316, new_AGEMA_signal_4315, RoundReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3810, new_AGEMA_signal_3809, new_AGEMA_signal_3808, RoundOutput[106]}), .a ({plaintext_s3[106], plaintext_s2[106], plaintext_s1[106], plaintext_s0[106]}), .c ({new_AGEMA_signal_4323, new_AGEMA_signal_4322, new_AGEMA_signal_4321, RoundReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, new_AGEMA_signal_3811, RoundOutput[107]}), .a ({plaintext_s3[107], plaintext_s2[107], plaintext_s1[107], plaintext_s0[107]}), .c ({new_AGEMA_signal_4329, new_AGEMA_signal_4328, new_AGEMA_signal_4327, RoundReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3816, new_AGEMA_signal_3815, new_AGEMA_signal_3814, RoundOutput[108]}), .a ({plaintext_s3[108], plaintext_s2[108], plaintext_s1[108], plaintext_s0[108]}), .c ({new_AGEMA_signal_4335, new_AGEMA_signal_4334, new_AGEMA_signal_4333, RoundReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, new_AGEMA_signal_3817, RoundOutput[109]}), .a ({plaintext_s3[109], plaintext_s2[109], plaintext_s1[109], plaintext_s0[109]}), .c ({new_AGEMA_signal_4341, new_AGEMA_signal_4340, new_AGEMA_signal_4339, RoundReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3822, new_AGEMA_signal_3821, new_AGEMA_signal_3820, RoundOutput[110]}), .a ({plaintext_s3[110], plaintext_s2[110], plaintext_s1[110], plaintext_s0[110]}), .c ({new_AGEMA_signal_4347, new_AGEMA_signal_4346, new_AGEMA_signal_4345, RoundReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, new_AGEMA_signal_3823, RoundOutput[111]}), .a ({plaintext_s3[111], plaintext_s2[111], plaintext_s1[111], plaintext_s0[111]}), .c ({new_AGEMA_signal_4353, new_AGEMA_signal_4352, new_AGEMA_signal_4351, RoundReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3828, new_AGEMA_signal_3827, new_AGEMA_signal_3826, RoundOutput[112]}), .a ({plaintext_s3[112], plaintext_s2[112], plaintext_s1[112], plaintext_s0[112]}), .c ({new_AGEMA_signal_4359, new_AGEMA_signal_4358, new_AGEMA_signal_4357, RoundReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, new_AGEMA_signal_3829, RoundOutput[113]}), .a ({plaintext_s3[113], plaintext_s2[113], plaintext_s1[113], plaintext_s0[113]}), .c ({new_AGEMA_signal_4365, new_AGEMA_signal_4364, new_AGEMA_signal_4363, RoundReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3834, new_AGEMA_signal_3833, new_AGEMA_signal_3832, RoundOutput[114]}), .a ({plaintext_s3[114], plaintext_s2[114], plaintext_s1[114], plaintext_s0[114]}), .c ({new_AGEMA_signal_4371, new_AGEMA_signal_4370, new_AGEMA_signal_4369, RoundReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, new_AGEMA_signal_3835, RoundOutput[115]}), .a ({plaintext_s3[115], plaintext_s2[115], plaintext_s1[115], plaintext_s0[115]}), .c ({new_AGEMA_signal_4377, new_AGEMA_signal_4376, new_AGEMA_signal_4375, RoundReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3840, new_AGEMA_signal_3839, new_AGEMA_signal_3838, RoundOutput[116]}), .a ({plaintext_s3[116], plaintext_s2[116], plaintext_s1[116], plaintext_s0[116]}), .c ({new_AGEMA_signal_4383, new_AGEMA_signal_4382, new_AGEMA_signal_4381, RoundReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, new_AGEMA_signal_3841, RoundOutput[117]}), .a ({plaintext_s3[117], plaintext_s2[117], plaintext_s1[117], plaintext_s0[117]}), .c ({new_AGEMA_signal_4389, new_AGEMA_signal_4388, new_AGEMA_signal_4387, RoundReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3846, new_AGEMA_signal_3845, new_AGEMA_signal_3844, RoundOutput[118]}), .a ({plaintext_s3[118], plaintext_s2[118], plaintext_s1[118], plaintext_s0[118]}), .c ({new_AGEMA_signal_4395, new_AGEMA_signal_4394, new_AGEMA_signal_4393, RoundReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, new_AGEMA_signal_3847, RoundOutput[119]}), .a ({plaintext_s3[119], plaintext_s2[119], plaintext_s1[119], plaintext_s0[119]}), .c ({new_AGEMA_signal_4401, new_AGEMA_signal_4400, new_AGEMA_signal_4399, RoundReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3852, new_AGEMA_signal_3851, new_AGEMA_signal_3850, RoundOutput[120]}), .a ({plaintext_s3[120], plaintext_s2[120], plaintext_s1[120], plaintext_s0[120]}), .c ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, new_AGEMA_signal_4405, RoundReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, new_AGEMA_signal_3853, RoundOutput[121]}), .a ({plaintext_s3[121], plaintext_s2[121], plaintext_s1[121], plaintext_s0[121]}), .c ({new_AGEMA_signal_4413, new_AGEMA_signal_4412, new_AGEMA_signal_4411, RoundReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3858, new_AGEMA_signal_3857, new_AGEMA_signal_3856, RoundOutput[122]}), .a ({plaintext_s3[122], plaintext_s2[122], plaintext_s1[122], plaintext_s0[122]}), .c ({new_AGEMA_signal_4419, new_AGEMA_signal_4418, new_AGEMA_signal_4417, RoundReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, new_AGEMA_signal_3859, RoundOutput[123]}), .a ({plaintext_s3[123], plaintext_s2[123], plaintext_s1[123], plaintext_s0[123]}), .c ({new_AGEMA_signal_4425, new_AGEMA_signal_4424, new_AGEMA_signal_4423, RoundReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3864, new_AGEMA_signal_3863, new_AGEMA_signal_3862, RoundOutput[124]}), .a ({plaintext_s3[124], plaintext_s2[124], plaintext_s1[124], plaintext_s0[124]}), .c ({new_AGEMA_signal_4431, new_AGEMA_signal_4430, new_AGEMA_signal_4429, RoundReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, new_AGEMA_signal_3865, RoundOutput[125]}), .a ({plaintext_s3[125], plaintext_s2[125], plaintext_s1[125], plaintext_s0[125]}), .c ({new_AGEMA_signal_4437, new_AGEMA_signal_4436, new_AGEMA_signal_4435, RoundReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3870, new_AGEMA_signal_3869, new_AGEMA_signal_3868, RoundOutput[126]}), .a ({plaintext_s3[126], plaintext_s2[126], plaintext_s1[126], plaintext_s0[126]}), .c ({new_AGEMA_signal_4443, new_AGEMA_signal_4442, new_AGEMA_signal_4441, RoundReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, new_AGEMA_signal_3871, RoundOutput[127]}), .a ({plaintext_s3[127], plaintext_s2[127], plaintext_s1[127], plaintext_s0[127]}), .c ({new_AGEMA_signal_4449, new_AGEMA_signal_4448, new_AGEMA_signal_4447, RoundReg_Inst_ff_SDE_127_next_state}) ) ;
    INV_X1 MuxSboxIn_U3 ( .A (AKSRnotDone), .ZN (MuxSboxIn_n7) ) ;
    INV_X1 MuxSboxIn_U2 ( .A (MuxSboxIn_n7), .ZN (MuxSboxIn_n5) ) ;
    INV_X1 MuxSboxIn_U1 ( .A (MuxSboxIn_n7), .ZN (MuxSboxIn_n6) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_0_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .a ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, new_AGEMA_signal_2656, KSSubBytesInput[0]}), .c ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, new_AGEMA_signal_3493, SubBytesInput[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_1_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .a ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, new_AGEMA_signal_2665, KSSubBytesInput[1]}), .c ({new_AGEMA_signal_3498, new_AGEMA_signal_3497, new_AGEMA_signal_3496, SubBytesInput[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_2_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .a ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, new_AGEMA_signal_2674, KSSubBytesInput[2]}), .c ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, new_AGEMA_signal_3499, SubBytesInput[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_3_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s3[3], ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .a ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, new_AGEMA_signal_2683, KSSubBytesInput[3]}), .c ({new_AGEMA_signal_3504, new_AGEMA_signal_3503, new_AGEMA_signal_3502, SubBytesInput[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_4_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .a ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, new_AGEMA_signal_2701, KSSubBytesInput[4]}), .c ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, new_AGEMA_signal_3505, SubBytesInput[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_5_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s3[5], ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .a ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, new_AGEMA_signal_2710, KSSubBytesInput[5]}), .c ({new_AGEMA_signal_3510, new_AGEMA_signal_3509, new_AGEMA_signal_3508, SubBytesInput[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_6_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s3[6], ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .a ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, new_AGEMA_signal_2719, KSSubBytesInput[6]}), .c ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, new_AGEMA_signal_3511, SubBytesInput[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_7_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .a ({new_AGEMA_signal_2730, new_AGEMA_signal_2729, new_AGEMA_signal_2728, KSSubBytesInput[7]}), .c ({new_AGEMA_signal_3516, new_AGEMA_signal_3515, new_AGEMA_signal_3514, SubBytesInput[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_8_U1 ( .s (AKSRnotDone), .b ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .a ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, new_AGEMA_signal_3385, KSSubBytesInput[8]}), .c ({new_AGEMA_signal_3492, new_AGEMA_signal_3491, new_AGEMA_signal_3490, SubBytesInput[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_9_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .a ({new_AGEMA_signal_3486, new_AGEMA_signal_3485, new_AGEMA_signal_3484, KSSubBytesInput[9]}), .c ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, new_AGEMA_signal_3517, SubBytesInput[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_10_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .a ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, new_AGEMA_signal_2440, KSSubBytesInput[10]}), .c ({new_AGEMA_signal_3522, new_AGEMA_signal_3521, new_AGEMA_signal_3520, SubBytesInput[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_11_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[43], ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .a ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, new_AGEMA_signal_2539, KSSubBytesInput[11]}), .c ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, new_AGEMA_signal_3523, SubBytesInput[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_12_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .a ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, new_AGEMA_signal_2620, KSSubBytesInput[12]}), .c ({new_AGEMA_signal_3528, new_AGEMA_signal_3527, new_AGEMA_signal_3526, SubBytesInput[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_13_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s3[45], ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .a ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, new_AGEMA_signal_2629, KSSubBytesInput[13]}), .c ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, new_AGEMA_signal_3529, SubBytesInput[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_14_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s3[46], ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .a ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, new_AGEMA_signal_2638, KSSubBytesInput[14]}), .c ({new_AGEMA_signal_3534, new_AGEMA_signal_3533, new_AGEMA_signal_3532, SubBytesInput[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_15_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .a ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, new_AGEMA_signal_2647, KSSubBytesInput[15]}), .c ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, new_AGEMA_signal_3535, SubBytesInput[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_16_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .a ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, new_AGEMA_signal_2341, KSSubBytesInput[16]}), .c ({new_AGEMA_signal_3540, new_AGEMA_signal_3539, new_AGEMA_signal_3538, SubBytesInput[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_17_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[81], ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .a ({new_AGEMA_signal_2694, new_AGEMA_signal_2693, new_AGEMA_signal_2692, KSSubBytesInput[17]}), .c ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, new_AGEMA_signal_3541, SubBytesInput[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_18_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[82], ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .a ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, new_AGEMA_signal_2791, KSSubBytesInput[18]}), .c ({new_AGEMA_signal_3546, new_AGEMA_signal_3545, new_AGEMA_signal_3544, SubBytesInput[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_19_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[83], ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}), .a ({new_AGEMA_signal_2892, new_AGEMA_signal_2891, new_AGEMA_signal_2890, KSSubBytesInput[19]}), .c ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, new_AGEMA_signal_3547, SubBytesInput[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_20_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[84], ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .a ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, new_AGEMA_signal_2989, KSSubBytesInput[20]}), .c ({new_AGEMA_signal_3552, new_AGEMA_signal_3551, new_AGEMA_signal_3550, SubBytesInput[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_21_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[85], ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}), .a ({new_AGEMA_signal_3090, new_AGEMA_signal_3089, new_AGEMA_signal_3088, KSSubBytesInput[21]}), .c ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, new_AGEMA_signal_3553, SubBytesInput[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_22_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[86], ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}), .a ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, new_AGEMA_signal_3187, KSSubBytesInput[22]}), .c ({new_AGEMA_signal_3558, new_AGEMA_signal_3557, new_AGEMA_signal_3556, SubBytesInput[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_23_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[87], ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .a ({new_AGEMA_signal_3288, new_AGEMA_signal_3287, new_AGEMA_signal_3286, KSSubBytesInput[23]}), .c ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, new_AGEMA_signal_3559, SubBytesInput[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_24_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .a ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, new_AGEMA_signal_2737, KSSubBytesInput[24]}), .c ({new_AGEMA_signal_3564, new_AGEMA_signal_3563, new_AGEMA_signal_3562, SubBytesInput[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_25_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .a ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, new_AGEMA_signal_2746, KSSubBytesInput[25]}), .c ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, new_AGEMA_signal_3565, SubBytesInput[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_26_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .a ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, new_AGEMA_signal_2755, KSSubBytesInput[26]}), .c ({new_AGEMA_signal_3570, new_AGEMA_signal_3569, new_AGEMA_signal_3568, SubBytesInput[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_27_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[123], ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .a ({new_AGEMA_signal_2766, new_AGEMA_signal_2765, new_AGEMA_signal_2764, KSSubBytesInput[27]}), .c ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, new_AGEMA_signal_3571, SubBytesInput[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_28_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .a ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, new_AGEMA_signal_2773, KSSubBytesInput[28]}), .c ({new_AGEMA_signal_3576, new_AGEMA_signal_3575, new_AGEMA_signal_3574, SubBytesInput[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_29_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .a ({new_AGEMA_signal_2784, new_AGEMA_signal_2783, new_AGEMA_signal_2782, KSSubBytesInput[29]}), .c ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, new_AGEMA_signal_3577, SubBytesInput[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_30_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .a ({new_AGEMA_signal_2802, new_AGEMA_signal_2801, new_AGEMA_signal_2800, KSSubBytesInput[30]}), .c ({new_AGEMA_signal_3582, new_AGEMA_signal_3581, new_AGEMA_signal_3580, SubBytesInput[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxSboxIn_mux_inst_31_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .a ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, new_AGEMA_signal_2809, KSSubBytesInput[31]}), .c ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, new_AGEMA_signal_3583, SubBytesInput[31]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T1_U1 ( .a ({new_AGEMA_signal_3516, new_AGEMA_signal_3515, new_AGEMA_signal_3514, SubBytesInput[7]}), .b ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, new_AGEMA_signal_3505, SubBytesInput[4]}), .c ({new_AGEMA_signal_4452, new_AGEMA_signal_4451, new_AGEMA_signal_4450, SubBytesIns_Inst_Sbox_0_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T2_U1 ( .a ({new_AGEMA_signal_3516, new_AGEMA_signal_3515, new_AGEMA_signal_3514, SubBytesInput[7]}), .b ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, new_AGEMA_signal_3499, SubBytesInput[2]}), .c ({new_AGEMA_signal_4455, new_AGEMA_signal_4454, new_AGEMA_signal_4453, SubBytesIns_Inst_Sbox_0_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T3_U1 ( .a ({new_AGEMA_signal_3516, new_AGEMA_signal_3515, new_AGEMA_signal_3514, SubBytesInput[7]}), .b ({new_AGEMA_signal_3498, new_AGEMA_signal_3497, new_AGEMA_signal_3496, SubBytesInput[1]}), .c ({new_AGEMA_signal_4458, new_AGEMA_signal_4457, new_AGEMA_signal_4456, SubBytesIns_Inst_Sbox_0_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T4_U1 ( .a ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, new_AGEMA_signal_3505, SubBytesInput[4]}), .b ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, new_AGEMA_signal_3499, SubBytesInput[2]}), .c ({new_AGEMA_signal_4461, new_AGEMA_signal_4460, new_AGEMA_signal_4459, SubBytesIns_Inst_Sbox_0_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T5_U1 ( .a ({new_AGEMA_signal_3504, new_AGEMA_signal_3503, new_AGEMA_signal_3502, SubBytesInput[3]}), .b ({new_AGEMA_signal_3498, new_AGEMA_signal_3497, new_AGEMA_signal_3496, SubBytesInput[1]}), .c ({new_AGEMA_signal_4464, new_AGEMA_signal_4463, new_AGEMA_signal_4462, SubBytesIns_Inst_Sbox_0_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_4452, new_AGEMA_signal_4451, new_AGEMA_signal_4450, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_4464, new_AGEMA_signal_4463, new_AGEMA_signal_4462, SubBytesIns_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_4572, new_AGEMA_signal_4571, new_AGEMA_signal_4570, SubBytesIns_Inst_Sbox_0_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T7_U1 ( .a ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, new_AGEMA_signal_3511, SubBytesInput[6]}), .b ({new_AGEMA_signal_3510, new_AGEMA_signal_3509, new_AGEMA_signal_3508, SubBytesInput[5]}), .c ({new_AGEMA_signal_4467, new_AGEMA_signal_4466, new_AGEMA_signal_4465, SubBytesIns_Inst_Sbox_0_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T8_U1 ( .a ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, new_AGEMA_signal_3493, SubBytesInput[0]}), .b ({new_AGEMA_signal_4572, new_AGEMA_signal_4571, new_AGEMA_signal_4570, SubBytesIns_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_4668, new_AGEMA_signal_4667, new_AGEMA_signal_4666, SubBytesIns_Inst_Sbox_0_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T9_U1 ( .a ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, new_AGEMA_signal_3493, SubBytesInput[0]}), .b ({new_AGEMA_signal_4467, new_AGEMA_signal_4466, new_AGEMA_signal_4465, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, new_AGEMA_signal_4573, SubBytesIns_Inst_Sbox_0_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_4572, new_AGEMA_signal_4571, new_AGEMA_signal_4570, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_4467, new_AGEMA_signal_4466, new_AGEMA_signal_4465, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, new_AGEMA_signal_4669, SubBytesIns_Inst_Sbox_0_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T11_U1 ( .a ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, new_AGEMA_signal_3511, SubBytesInput[6]}), .b ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, new_AGEMA_signal_3499, SubBytesInput[2]}), .c ({new_AGEMA_signal_4470, new_AGEMA_signal_4469, new_AGEMA_signal_4468, SubBytesIns_Inst_Sbox_0_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T12_U1 ( .a ({new_AGEMA_signal_3510, new_AGEMA_signal_3509, new_AGEMA_signal_3508, SubBytesInput[5]}), .b ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, new_AGEMA_signal_3499, SubBytesInput[2]}), .c ({new_AGEMA_signal_4473, new_AGEMA_signal_4472, new_AGEMA_signal_4471, SubBytesIns_Inst_Sbox_0_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_4458, new_AGEMA_signal_4457, new_AGEMA_signal_4456, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_4461, new_AGEMA_signal_4460, new_AGEMA_signal_4459, SubBytesIns_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_4578, new_AGEMA_signal_4577, new_AGEMA_signal_4576, SubBytesIns_Inst_Sbox_0_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_4572, new_AGEMA_signal_4571, new_AGEMA_signal_4570, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_4470, new_AGEMA_signal_4469, new_AGEMA_signal_4468, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_4674, new_AGEMA_signal_4673, new_AGEMA_signal_4672, SubBytesIns_Inst_Sbox_0_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_4464, new_AGEMA_signal_4463, new_AGEMA_signal_4462, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_4470, new_AGEMA_signal_4469, new_AGEMA_signal_4468, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, new_AGEMA_signal_4579, SubBytesIns_Inst_Sbox_0_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_4464, new_AGEMA_signal_4463, new_AGEMA_signal_4462, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_4473, new_AGEMA_signal_4472, new_AGEMA_signal_4471, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_4584, new_AGEMA_signal_4583, new_AGEMA_signal_4582, SubBytesIns_Inst_Sbox_0_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, new_AGEMA_signal_4573, SubBytesIns_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_4584, new_AGEMA_signal_4583, new_AGEMA_signal_4582, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_4677, new_AGEMA_signal_4676, new_AGEMA_signal_4675, SubBytesIns_Inst_Sbox_0_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T18_U1 ( .a ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, new_AGEMA_signal_3505, SubBytesInput[4]}), .b ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, new_AGEMA_signal_3493, SubBytesInput[0]}), .c ({new_AGEMA_signal_4476, new_AGEMA_signal_4475, new_AGEMA_signal_4474, SubBytesIns_Inst_Sbox_0_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_4467, new_AGEMA_signal_4466, new_AGEMA_signal_4465, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_4476, new_AGEMA_signal_4475, new_AGEMA_signal_4474, SubBytesIns_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_4587, new_AGEMA_signal_4586, new_AGEMA_signal_4585, SubBytesIns_Inst_Sbox_0_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_4452, new_AGEMA_signal_4451, new_AGEMA_signal_4450, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_4587, new_AGEMA_signal_4586, new_AGEMA_signal_4585, SubBytesIns_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_4680, new_AGEMA_signal_4679, new_AGEMA_signal_4678, SubBytesIns_Inst_Sbox_0_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T21_U1 ( .a ({new_AGEMA_signal_3498, new_AGEMA_signal_3497, new_AGEMA_signal_3496, SubBytesInput[1]}), .b ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, new_AGEMA_signal_3493, SubBytesInput[0]}), .c ({new_AGEMA_signal_4479, new_AGEMA_signal_4478, new_AGEMA_signal_4477, SubBytesIns_Inst_Sbox_0_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_4467, new_AGEMA_signal_4466, new_AGEMA_signal_4465, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_4479, new_AGEMA_signal_4478, new_AGEMA_signal_4477, SubBytesIns_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_4590, new_AGEMA_signal_4589, new_AGEMA_signal_4588, SubBytesIns_Inst_Sbox_0_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_4455, new_AGEMA_signal_4454, new_AGEMA_signal_4453, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_4590, new_AGEMA_signal_4589, new_AGEMA_signal_4588, SubBytesIns_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_4683, new_AGEMA_signal_4682, new_AGEMA_signal_4681, SubBytesIns_Inst_Sbox_0_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_4455, new_AGEMA_signal_4454, new_AGEMA_signal_4453, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, new_AGEMA_signal_4669, SubBytesIns_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_4824, new_AGEMA_signal_4823, new_AGEMA_signal_4822, SubBytesIns_Inst_Sbox_0_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_4680, new_AGEMA_signal_4679, new_AGEMA_signal_4678, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_4677, new_AGEMA_signal_4676, new_AGEMA_signal_4675, SubBytesIns_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_4827, new_AGEMA_signal_4826, new_AGEMA_signal_4825, SubBytesIns_Inst_Sbox_0_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_4458, new_AGEMA_signal_4457, new_AGEMA_signal_4456, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_4584, new_AGEMA_signal_4583, new_AGEMA_signal_4582, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_4686, new_AGEMA_signal_4685, new_AGEMA_signal_4684, SubBytesIns_Inst_Sbox_0_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_4452, new_AGEMA_signal_4451, new_AGEMA_signal_4450, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_4473, new_AGEMA_signal_4472, new_AGEMA_signal_4471, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, new_AGEMA_signal_4591, SubBytesIns_Inst_Sbox_0_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T1_U1 ( .a ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, new_AGEMA_signal_3535, SubBytesInput[15]}), .b ({new_AGEMA_signal_3528, new_AGEMA_signal_3527, new_AGEMA_signal_3526, SubBytesInput[12]}), .c ({new_AGEMA_signal_4482, new_AGEMA_signal_4481, new_AGEMA_signal_4480, SubBytesIns_Inst_Sbox_1_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T2_U1 ( .a ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, new_AGEMA_signal_3535, SubBytesInput[15]}), .b ({new_AGEMA_signal_3522, new_AGEMA_signal_3521, new_AGEMA_signal_3520, SubBytesInput[10]}), .c ({new_AGEMA_signal_4485, new_AGEMA_signal_4484, new_AGEMA_signal_4483, SubBytesIns_Inst_Sbox_1_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T3_U1 ( .a ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, new_AGEMA_signal_3535, SubBytesInput[15]}), .b ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, new_AGEMA_signal_3517, SubBytesInput[9]}), .c ({new_AGEMA_signal_4488, new_AGEMA_signal_4487, new_AGEMA_signal_4486, SubBytesIns_Inst_Sbox_1_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T4_U1 ( .a ({new_AGEMA_signal_3528, new_AGEMA_signal_3527, new_AGEMA_signal_3526, SubBytesInput[12]}), .b ({new_AGEMA_signal_3522, new_AGEMA_signal_3521, new_AGEMA_signal_3520, SubBytesInput[10]}), .c ({new_AGEMA_signal_4491, new_AGEMA_signal_4490, new_AGEMA_signal_4489, SubBytesIns_Inst_Sbox_1_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T5_U1 ( .a ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, new_AGEMA_signal_3523, SubBytesInput[11]}), .b ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, new_AGEMA_signal_3517, SubBytesInput[9]}), .c ({new_AGEMA_signal_4494, new_AGEMA_signal_4493, new_AGEMA_signal_4492, SubBytesIns_Inst_Sbox_1_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_4482, new_AGEMA_signal_4481, new_AGEMA_signal_4480, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_4494, new_AGEMA_signal_4493, new_AGEMA_signal_4492, SubBytesIns_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_4596, new_AGEMA_signal_4595, new_AGEMA_signal_4594, SubBytesIns_Inst_Sbox_1_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T7_U1 ( .a ({new_AGEMA_signal_3534, new_AGEMA_signal_3533, new_AGEMA_signal_3532, SubBytesInput[14]}), .b ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, new_AGEMA_signal_3529, SubBytesInput[13]}), .c ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, new_AGEMA_signal_4495, SubBytesIns_Inst_Sbox_1_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T8_U1 ( .a ({new_AGEMA_signal_3492, new_AGEMA_signal_3491, new_AGEMA_signal_3490, SubBytesInput[8]}), .b ({new_AGEMA_signal_4596, new_AGEMA_signal_4595, new_AGEMA_signal_4594, SubBytesIns_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_4707, new_AGEMA_signal_4706, new_AGEMA_signal_4705, SubBytesIns_Inst_Sbox_1_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T9_U1 ( .a ({new_AGEMA_signal_3492, new_AGEMA_signal_3491, new_AGEMA_signal_3490, SubBytesInput[8]}), .b ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, new_AGEMA_signal_4495, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, new_AGEMA_signal_4597, SubBytesIns_Inst_Sbox_1_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_4596, new_AGEMA_signal_4595, new_AGEMA_signal_4594, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, new_AGEMA_signal_4495, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_4710, new_AGEMA_signal_4709, new_AGEMA_signal_4708, SubBytesIns_Inst_Sbox_1_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T11_U1 ( .a ({new_AGEMA_signal_3534, new_AGEMA_signal_3533, new_AGEMA_signal_3532, SubBytesInput[14]}), .b ({new_AGEMA_signal_3522, new_AGEMA_signal_3521, new_AGEMA_signal_3520, SubBytesInput[10]}), .c ({new_AGEMA_signal_4500, new_AGEMA_signal_4499, new_AGEMA_signal_4498, SubBytesIns_Inst_Sbox_1_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T12_U1 ( .a ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, new_AGEMA_signal_3529, SubBytesInput[13]}), .b ({new_AGEMA_signal_3522, new_AGEMA_signal_3521, new_AGEMA_signal_3520, SubBytesInput[10]}), .c ({new_AGEMA_signal_4503, new_AGEMA_signal_4502, new_AGEMA_signal_4501, SubBytesIns_Inst_Sbox_1_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_4488, new_AGEMA_signal_4487, new_AGEMA_signal_4486, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_4491, new_AGEMA_signal_4490, new_AGEMA_signal_4489, SubBytesIns_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_4602, new_AGEMA_signal_4601, new_AGEMA_signal_4600, SubBytesIns_Inst_Sbox_1_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_4596, new_AGEMA_signal_4595, new_AGEMA_signal_4594, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_4500, new_AGEMA_signal_4499, new_AGEMA_signal_4498, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, new_AGEMA_signal_4711, SubBytesIns_Inst_Sbox_1_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_4494, new_AGEMA_signal_4493, new_AGEMA_signal_4492, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_4500, new_AGEMA_signal_4499, new_AGEMA_signal_4498, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_4605, new_AGEMA_signal_4604, new_AGEMA_signal_4603, SubBytesIns_Inst_Sbox_1_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_4494, new_AGEMA_signal_4493, new_AGEMA_signal_4492, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_4503, new_AGEMA_signal_4502, new_AGEMA_signal_4501, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_4608, new_AGEMA_signal_4607, new_AGEMA_signal_4606, SubBytesIns_Inst_Sbox_1_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, new_AGEMA_signal_4597, SubBytesIns_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_4608, new_AGEMA_signal_4607, new_AGEMA_signal_4606, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_4716, new_AGEMA_signal_4715, new_AGEMA_signal_4714, SubBytesIns_Inst_Sbox_1_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T18_U1 ( .a ({new_AGEMA_signal_3528, new_AGEMA_signal_3527, new_AGEMA_signal_3526, SubBytesInput[12]}), .b ({new_AGEMA_signal_3492, new_AGEMA_signal_3491, new_AGEMA_signal_3490, SubBytesInput[8]}), .c ({new_AGEMA_signal_4506, new_AGEMA_signal_4505, new_AGEMA_signal_4504, SubBytesIns_Inst_Sbox_1_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, new_AGEMA_signal_4495, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_4506, new_AGEMA_signal_4505, new_AGEMA_signal_4504, SubBytesIns_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_4611, new_AGEMA_signal_4610, new_AGEMA_signal_4609, SubBytesIns_Inst_Sbox_1_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_4482, new_AGEMA_signal_4481, new_AGEMA_signal_4480, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_4611, new_AGEMA_signal_4610, new_AGEMA_signal_4609, SubBytesIns_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, new_AGEMA_signal_4717, SubBytesIns_Inst_Sbox_1_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T21_U1 ( .a ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, new_AGEMA_signal_3517, SubBytesInput[9]}), .b ({new_AGEMA_signal_3492, new_AGEMA_signal_3491, new_AGEMA_signal_3490, SubBytesInput[8]}), .c ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, new_AGEMA_signal_4507, SubBytesIns_Inst_Sbox_1_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, new_AGEMA_signal_4495, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, new_AGEMA_signal_4507, SubBytesIns_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_4614, new_AGEMA_signal_4613, new_AGEMA_signal_4612, SubBytesIns_Inst_Sbox_1_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_4485, new_AGEMA_signal_4484, new_AGEMA_signal_4483, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_4614, new_AGEMA_signal_4613, new_AGEMA_signal_4612, SubBytesIns_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_4722, new_AGEMA_signal_4721, new_AGEMA_signal_4720, SubBytesIns_Inst_Sbox_1_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_4485, new_AGEMA_signal_4484, new_AGEMA_signal_4483, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_4710, new_AGEMA_signal_4709, new_AGEMA_signal_4708, SubBytesIns_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, new_AGEMA_signal_4849, SubBytesIns_Inst_Sbox_1_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, new_AGEMA_signal_4717, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_4716, new_AGEMA_signal_4715, new_AGEMA_signal_4714, SubBytesIns_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_4854, new_AGEMA_signal_4853, new_AGEMA_signal_4852, SubBytesIns_Inst_Sbox_1_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_4488, new_AGEMA_signal_4487, new_AGEMA_signal_4486, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_4608, new_AGEMA_signal_4607, new_AGEMA_signal_4606, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, new_AGEMA_signal_4723, SubBytesIns_Inst_Sbox_1_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_4482, new_AGEMA_signal_4481, new_AGEMA_signal_4480, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_4503, new_AGEMA_signal_4502, new_AGEMA_signal_4501, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, new_AGEMA_signal_4615, SubBytesIns_Inst_Sbox_1_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T1_U1 ( .a ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, new_AGEMA_signal_3559, SubBytesInput[23]}), .b ({new_AGEMA_signal_3552, new_AGEMA_signal_3551, new_AGEMA_signal_3550, SubBytesInput[20]}), .c ({new_AGEMA_signal_4512, new_AGEMA_signal_4511, new_AGEMA_signal_4510, SubBytesIns_Inst_Sbox_2_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T2_U1 ( .a ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, new_AGEMA_signal_3559, SubBytesInput[23]}), .b ({new_AGEMA_signal_3546, new_AGEMA_signal_3545, new_AGEMA_signal_3544, SubBytesInput[18]}), .c ({new_AGEMA_signal_4515, new_AGEMA_signal_4514, new_AGEMA_signal_4513, SubBytesIns_Inst_Sbox_2_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T3_U1 ( .a ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, new_AGEMA_signal_3559, SubBytesInput[23]}), .b ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, new_AGEMA_signal_3541, SubBytesInput[17]}), .c ({new_AGEMA_signal_4518, new_AGEMA_signal_4517, new_AGEMA_signal_4516, SubBytesIns_Inst_Sbox_2_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T4_U1 ( .a ({new_AGEMA_signal_3552, new_AGEMA_signal_3551, new_AGEMA_signal_3550, SubBytesInput[20]}), .b ({new_AGEMA_signal_3546, new_AGEMA_signal_3545, new_AGEMA_signal_3544, SubBytesInput[18]}), .c ({new_AGEMA_signal_4521, new_AGEMA_signal_4520, new_AGEMA_signal_4519, SubBytesIns_Inst_Sbox_2_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T5_U1 ( .a ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, new_AGEMA_signal_3547, SubBytesInput[19]}), .b ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, new_AGEMA_signal_3541, SubBytesInput[17]}), .c ({new_AGEMA_signal_4524, new_AGEMA_signal_4523, new_AGEMA_signal_4522, SubBytesIns_Inst_Sbox_2_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_4512, new_AGEMA_signal_4511, new_AGEMA_signal_4510, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_4524, new_AGEMA_signal_4523, new_AGEMA_signal_4522, SubBytesIns_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_4620, new_AGEMA_signal_4619, new_AGEMA_signal_4618, SubBytesIns_Inst_Sbox_2_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T7_U1 ( .a ({new_AGEMA_signal_3558, new_AGEMA_signal_3557, new_AGEMA_signal_3556, SubBytesInput[22]}), .b ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, new_AGEMA_signal_3553, SubBytesInput[21]}), .c ({new_AGEMA_signal_4527, new_AGEMA_signal_4526, new_AGEMA_signal_4525, SubBytesIns_Inst_Sbox_2_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T8_U1 ( .a ({new_AGEMA_signal_3540, new_AGEMA_signal_3539, new_AGEMA_signal_3538, SubBytesInput[16]}), .b ({new_AGEMA_signal_4620, new_AGEMA_signal_4619, new_AGEMA_signal_4618, SubBytesIns_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_4746, new_AGEMA_signal_4745, new_AGEMA_signal_4744, SubBytesIns_Inst_Sbox_2_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T9_U1 ( .a ({new_AGEMA_signal_3540, new_AGEMA_signal_3539, new_AGEMA_signal_3538, SubBytesInput[16]}), .b ({new_AGEMA_signal_4527, new_AGEMA_signal_4526, new_AGEMA_signal_4525, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_4623, new_AGEMA_signal_4622, new_AGEMA_signal_4621, SubBytesIns_Inst_Sbox_2_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_4620, new_AGEMA_signal_4619, new_AGEMA_signal_4618, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_4527, new_AGEMA_signal_4526, new_AGEMA_signal_4525, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, new_AGEMA_signal_4747, SubBytesIns_Inst_Sbox_2_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T11_U1 ( .a ({new_AGEMA_signal_3558, new_AGEMA_signal_3557, new_AGEMA_signal_3556, SubBytesInput[22]}), .b ({new_AGEMA_signal_3546, new_AGEMA_signal_3545, new_AGEMA_signal_3544, SubBytesInput[18]}), .c ({new_AGEMA_signal_4530, new_AGEMA_signal_4529, new_AGEMA_signal_4528, SubBytesIns_Inst_Sbox_2_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T12_U1 ( .a ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, new_AGEMA_signal_3553, SubBytesInput[21]}), .b ({new_AGEMA_signal_3546, new_AGEMA_signal_3545, new_AGEMA_signal_3544, SubBytesInput[18]}), .c ({new_AGEMA_signal_4533, new_AGEMA_signal_4532, new_AGEMA_signal_4531, SubBytesIns_Inst_Sbox_2_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_4518, new_AGEMA_signal_4517, new_AGEMA_signal_4516, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_4521, new_AGEMA_signal_4520, new_AGEMA_signal_4519, SubBytesIns_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_4626, new_AGEMA_signal_4625, new_AGEMA_signal_4624, SubBytesIns_Inst_Sbox_2_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_4620, new_AGEMA_signal_4619, new_AGEMA_signal_4618, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_4530, new_AGEMA_signal_4529, new_AGEMA_signal_4528, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_4752, new_AGEMA_signal_4751, new_AGEMA_signal_4750, SubBytesIns_Inst_Sbox_2_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_4524, new_AGEMA_signal_4523, new_AGEMA_signal_4522, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_4530, new_AGEMA_signal_4529, new_AGEMA_signal_4528, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_4629, new_AGEMA_signal_4628, new_AGEMA_signal_4627, SubBytesIns_Inst_Sbox_2_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_4524, new_AGEMA_signal_4523, new_AGEMA_signal_4522, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_4533, new_AGEMA_signal_4532, new_AGEMA_signal_4531, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_4632, new_AGEMA_signal_4631, new_AGEMA_signal_4630, SubBytesIns_Inst_Sbox_2_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_4623, new_AGEMA_signal_4622, new_AGEMA_signal_4621, SubBytesIns_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_4632, new_AGEMA_signal_4631, new_AGEMA_signal_4630, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, new_AGEMA_signal_4753, SubBytesIns_Inst_Sbox_2_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T18_U1 ( .a ({new_AGEMA_signal_3552, new_AGEMA_signal_3551, new_AGEMA_signal_3550, SubBytesInput[20]}), .b ({new_AGEMA_signal_3540, new_AGEMA_signal_3539, new_AGEMA_signal_3538, SubBytesInput[16]}), .c ({new_AGEMA_signal_4536, new_AGEMA_signal_4535, new_AGEMA_signal_4534, SubBytesIns_Inst_Sbox_2_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_4527, new_AGEMA_signal_4526, new_AGEMA_signal_4525, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_4536, new_AGEMA_signal_4535, new_AGEMA_signal_4534, SubBytesIns_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_4635, new_AGEMA_signal_4634, new_AGEMA_signal_4633, SubBytesIns_Inst_Sbox_2_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_4512, new_AGEMA_signal_4511, new_AGEMA_signal_4510, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_4635, new_AGEMA_signal_4634, new_AGEMA_signal_4633, SubBytesIns_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_4758, new_AGEMA_signal_4757, new_AGEMA_signal_4756, SubBytesIns_Inst_Sbox_2_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T21_U1 ( .a ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, new_AGEMA_signal_3541, SubBytesInput[17]}), .b ({new_AGEMA_signal_3540, new_AGEMA_signal_3539, new_AGEMA_signal_3538, SubBytesInput[16]}), .c ({new_AGEMA_signal_4539, new_AGEMA_signal_4538, new_AGEMA_signal_4537, SubBytesIns_Inst_Sbox_2_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_4527, new_AGEMA_signal_4526, new_AGEMA_signal_4525, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_4539, new_AGEMA_signal_4538, new_AGEMA_signal_4537, SubBytesIns_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_4638, new_AGEMA_signal_4637, new_AGEMA_signal_4636, SubBytesIns_Inst_Sbox_2_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_4515, new_AGEMA_signal_4514, new_AGEMA_signal_4513, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_4638, new_AGEMA_signal_4637, new_AGEMA_signal_4636, SubBytesIns_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, new_AGEMA_signal_4759, SubBytesIns_Inst_Sbox_2_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_4515, new_AGEMA_signal_4514, new_AGEMA_signal_4513, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, new_AGEMA_signal_4747, SubBytesIns_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_4878, new_AGEMA_signal_4877, new_AGEMA_signal_4876, SubBytesIns_Inst_Sbox_2_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_4758, new_AGEMA_signal_4757, new_AGEMA_signal_4756, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, new_AGEMA_signal_4753, SubBytesIns_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_4881, new_AGEMA_signal_4880, new_AGEMA_signal_4879, SubBytesIns_Inst_Sbox_2_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_4518, new_AGEMA_signal_4517, new_AGEMA_signal_4516, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_4632, new_AGEMA_signal_4631, new_AGEMA_signal_4630, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_4764, new_AGEMA_signal_4763, new_AGEMA_signal_4762, SubBytesIns_Inst_Sbox_2_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_4512, new_AGEMA_signal_4511, new_AGEMA_signal_4510, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_4533, new_AGEMA_signal_4532, new_AGEMA_signal_4531, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_4641, new_AGEMA_signal_4640, new_AGEMA_signal_4639, SubBytesIns_Inst_Sbox_2_T27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T1_U1 ( .a ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, new_AGEMA_signal_3583, SubBytesInput[31]}), .b ({new_AGEMA_signal_3576, new_AGEMA_signal_3575, new_AGEMA_signal_3574, SubBytesInput[28]}), .c ({new_AGEMA_signal_4542, new_AGEMA_signal_4541, new_AGEMA_signal_4540, SubBytesIns_Inst_Sbox_3_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T2_U1 ( .a ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, new_AGEMA_signal_3583, SubBytesInput[31]}), .b ({new_AGEMA_signal_3570, new_AGEMA_signal_3569, new_AGEMA_signal_3568, SubBytesInput[26]}), .c ({new_AGEMA_signal_4545, new_AGEMA_signal_4544, new_AGEMA_signal_4543, SubBytesIns_Inst_Sbox_3_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T3_U1 ( .a ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, new_AGEMA_signal_3583, SubBytesInput[31]}), .b ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, new_AGEMA_signal_3565, SubBytesInput[25]}), .c ({new_AGEMA_signal_4548, new_AGEMA_signal_4547, new_AGEMA_signal_4546, SubBytesIns_Inst_Sbox_3_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T4_U1 ( .a ({new_AGEMA_signal_3576, new_AGEMA_signal_3575, new_AGEMA_signal_3574, SubBytesInput[28]}), .b ({new_AGEMA_signal_3570, new_AGEMA_signal_3569, new_AGEMA_signal_3568, SubBytesInput[26]}), .c ({new_AGEMA_signal_4551, new_AGEMA_signal_4550, new_AGEMA_signal_4549, SubBytesIns_Inst_Sbox_3_T4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T5_U1 ( .a ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, new_AGEMA_signal_3571, SubBytesInput[27]}), .b ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, new_AGEMA_signal_3565, SubBytesInput[25]}), .c ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, SubBytesIns_Inst_Sbox_3_T5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_4542, new_AGEMA_signal_4541, new_AGEMA_signal_4540, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, SubBytesIns_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_4644, new_AGEMA_signal_4643, new_AGEMA_signal_4642, SubBytesIns_Inst_Sbox_3_T6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T7_U1 ( .a ({new_AGEMA_signal_3582, new_AGEMA_signal_3581, new_AGEMA_signal_3580, SubBytesInput[30]}), .b ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, new_AGEMA_signal_3577, SubBytesInput[29]}), .c ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, new_AGEMA_signal_4555, SubBytesIns_Inst_Sbox_3_T7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T8_U1 ( .a ({new_AGEMA_signal_3564, new_AGEMA_signal_3563, new_AGEMA_signal_3562, SubBytesInput[24]}), .b ({new_AGEMA_signal_4644, new_AGEMA_signal_4643, new_AGEMA_signal_4642, SubBytesIns_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_4785, new_AGEMA_signal_4784, new_AGEMA_signal_4783, SubBytesIns_Inst_Sbox_3_T8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T9_U1 ( .a ({new_AGEMA_signal_3564, new_AGEMA_signal_3563, new_AGEMA_signal_3562, SubBytesInput[24]}), .b ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, new_AGEMA_signal_4555, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, new_AGEMA_signal_4645, SubBytesIns_Inst_Sbox_3_T9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_4644, new_AGEMA_signal_4643, new_AGEMA_signal_4642, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, new_AGEMA_signal_4555, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_4788, new_AGEMA_signal_4787, new_AGEMA_signal_4786, SubBytesIns_Inst_Sbox_3_T10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T11_U1 ( .a ({new_AGEMA_signal_3582, new_AGEMA_signal_3581, new_AGEMA_signal_3580, SubBytesInput[30]}), .b ({new_AGEMA_signal_3570, new_AGEMA_signal_3569, new_AGEMA_signal_3568, SubBytesInput[26]}), .c ({new_AGEMA_signal_4560, new_AGEMA_signal_4559, new_AGEMA_signal_4558, SubBytesIns_Inst_Sbox_3_T11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T12_U1 ( .a ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, new_AGEMA_signal_3577, SubBytesInput[29]}), .b ({new_AGEMA_signal_3570, new_AGEMA_signal_3569, new_AGEMA_signal_3568, SubBytesInput[26]}), .c ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, new_AGEMA_signal_4561, SubBytesIns_Inst_Sbox_3_T12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_4548, new_AGEMA_signal_4547, new_AGEMA_signal_4546, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_4551, new_AGEMA_signal_4550, new_AGEMA_signal_4549, SubBytesIns_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_4650, new_AGEMA_signal_4649, new_AGEMA_signal_4648, SubBytesIns_Inst_Sbox_3_T13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_4644, new_AGEMA_signal_4643, new_AGEMA_signal_4642, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_4560, new_AGEMA_signal_4559, new_AGEMA_signal_4558, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_4791, new_AGEMA_signal_4790, new_AGEMA_signal_4789, SubBytesIns_Inst_Sbox_3_T14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_4560, new_AGEMA_signal_4559, new_AGEMA_signal_4558, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, SubBytesIns_Inst_Sbox_3_T15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, new_AGEMA_signal_4561, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_4656, new_AGEMA_signal_4655, new_AGEMA_signal_4654, SubBytesIns_Inst_Sbox_3_T16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, new_AGEMA_signal_4645, SubBytesIns_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_4656, new_AGEMA_signal_4655, new_AGEMA_signal_4654, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_4794, new_AGEMA_signal_4793, new_AGEMA_signal_4792, SubBytesIns_Inst_Sbox_3_T17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T18_U1 ( .a ({new_AGEMA_signal_3576, new_AGEMA_signal_3575, new_AGEMA_signal_3574, SubBytesInput[28]}), .b ({new_AGEMA_signal_3564, new_AGEMA_signal_3563, new_AGEMA_signal_3562, SubBytesInput[24]}), .c ({new_AGEMA_signal_4566, new_AGEMA_signal_4565, new_AGEMA_signal_4564, SubBytesIns_Inst_Sbox_3_T18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, new_AGEMA_signal_4555, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_4566, new_AGEMA_signal_4565, new_AGEMA_signal_4564, SubBytesIns_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_4659, new_AGEMA_signal_4658, new_AGEMA_signal_4657, SubBytesIns_Inst_Sbox_3_T19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_4542, new_AGEMA_signal_4541, new_AGEMA_signal_4540, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_4659, new_AGEMA_signal_4658, new_AGEMA_signal_4657, SubBytesIns_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, new_AGEMA_signal_4795, SubBytesIns_Inst_Sbox_3_T20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T21_U1 ( .a ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, new_AGEMA_signal_3565, SubBytesInput[25]}), .b ({new_AGEMA_signal_3564, new_AGEMA_signal_3563, new_AGEMA_signal_3562, SubBytesInput[24]}), .c ({new_AGEMA_signal_4569, new_AGEMA_signal_4568, new_AGEMA_signal_4567, SubBytesIns_Inst_Sbox_3_T21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, new_AGEMA_signal_4555, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_4569, new_AGEMA_signal_4568, new_AGEMA_signal_4567, SubBytesIns_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_4662, new_AGEMA_signal_4661, new_AGEMA_signal_4660, SubBytesIns_Inst_Sbox_3_T22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_4545, new_AGEMA_signal_4544, new_AGEMA_signal_4543, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_4662, new_AGEMA_signal_4661, new_AGEMA_signal_4660, SubBytesIns_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_4800, new_AGEMA_signal_4799, new_AGEMA_signal_4798, SubBytesIns_Inst_Sbox_3_T23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_4545, new_AGEMA_signal_4544, new_AGEMA_signal_4543, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_4788, new_AGEMA_signal_4787, new_AGEMA_signal_4786, SubBytesIns_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, new_AGEMA_signal_4903, SubBytesIns_Inst_Sbox_3_T24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, new_AGEMA_signal_4795, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_4794, new_AGEMA_signal_4793, new_AGEMA_signal_4792, SubBytesIns_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_4908, new_AGEMA_signal_4907, new_AGEMA_signal_4906, SubBytesIns_Inst_Sbox_3_T25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_4548, new_AGEMA_signal_4547, new_AGEMA_signal_4546, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_4656, new_AGEMA_signal_4655, new_AGEMA_signal_4654, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_4803, new_AGEMA_signal_4802, new_AGEMA_signal_4801, SubBytesIns_Inst_Sbox_3_T26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_4542, new_AGEMA_signal_4541, new_AGEMA_signal_4540, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, new_AGEMA_signal_4561, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_4665, new_AGEMA_signal_4664, new_AGEMA_signal_4663, SubBytesIns_Inst_Sbox_3_T27}) ) ;
    INV_X1 MuxMCOut_U3 ( .A (LastRoundorDone), .ZN (MuxMCOut_n6) ) ;
    INV_X1 MuxMCOut_U2 ( .A (MuxMCOut_n6), .ZN (MuxMCOut_n5) ) ;
    INV_X1 MuxMCOut_U1 ( .A (MuxMCOut_n6), .ZN (MuxMCOut_n4) ) ;
    INV_X1 MuxRound_U7 ( .A (AKSRnotDone), .ZN (MuxRound_n19) ) ;
    INV_X1 MuxRound_U6 ( .A (MuxRound_n19), .ZN (MuxRound_n16) ) ;
    INV_X1 MuxRound_U5 ( .A (MuxRound_n19), .ZN (MuxRound_n14) ) ;
    INV_X1 MuxRound_U4 ( .A (MuxRound_n19), .ZN (MuxRound_n13) ) ;
    INV_X1 MuxRound_U3 ( .A (MuxRound_n19), .ZN (MuxRound_n15) ) ;
    INV_X1 MuxRound_U2 ( .A (MuxRound_n19), .ZN (MuxRound_n18) ) ;
    INV_X1 MuxRound_U1 ( .A (MuxRound_n19), .ZN (MuxRound_n17) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_32_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .a ({new_AGEMA_signal_3138, new_AGEMA_signal_3137, new_AGEMA_signal_3136, ShiftRowsOutput[32]}), .c ({new_AGEMA_signal_3588, new_AGEMA_signal_3587, new_AGEMA_signal_3586, RoundOutput[32]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_33_U1 ( .s (MuxRound_n17), .b ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .a ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, new_AGEMA_signal_3145, ShiftRowsOutput[33]}), .c ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, new_AGEMA_signal_3589, RoundOutput[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_34_U1 ( .s (MuxRound_n13), .b ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .a ({new_AGEMA_signal_3156, new_AGEMA_signal_3155, new_AGEMA_signal_3154, ShiftRowsOutput[34]}), .c ({new_AGEMA_signal_3594, new_AGEMA_signal_3593, new_AGEMA_signal_3592, RoundOutput[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_35_U1 ( .s (MuxRound_n14), .b ({ciphertext_s3[35], ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .a ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, new_AGEMA_signal_3163, ShiftRowsOutput[35]}), .c ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, new_AGEMA_signal_3595, RoundOutput[35]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_36_U1 ( .s (MuxRound_n15), .b ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .a ({new_AGEMA_signal_3174, new_AGEMA_signal_3173, new_AGEMA_signal_3172, ShiftRowsOutput[36]}), .c ({new_AGEMA_signal_3600, new_AGEMA_signal_3599, new_AGEMA_signal_3598, RoundOutput[36]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_37_U1 ( .s (MuxRound_n16), .b ({ciphertext_s3[37], ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .a ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, new_AGEMA_signal_3181, ShiftRowsOutput[37]}), .c ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, new_AGEMA_signal_3601, RoundOutput[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_38_U1 ( .s (MuxRound_n17), .b ({ciphertext_s3[38], ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .a ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, new_AGEMA_signal_3199, ShiftRowsOutput[38]}), .c ({new_AGEMA_signal_3606, new_AGEMA_signal_3605, new_AGEMA_signal_3604, RoundOutput[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_39_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .a ({new_AGEMA_signal_3210, new_AGEMA_signal_3209, new_AGEMA_signal_3208, ShiftRowsOutput[39]}), .c ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, new_AGEMA_signal_3607, RoundOutput[39]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_40_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .a ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, new_AGEMA_signal_2389, ShiftRowsOutput[40]}), .c ({new_AGEMA_signal_3612, new_AGEMA_signal_3611, new_AGEMA_signal_3610, RoundOutput[40]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_41_U1 ( .s (MuxRound_n13), .b ({ciphertext_s3[73], ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .a ({new_AGEMA_signal_2400, new_AGEMA_signal_2399, new_AGEMA_signal_2398, ShiftRowsOutput[41]}), .c ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, new_AGEMA_signal_3613, RoundOutput[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_42_U1 ( .s (MuxRound_n14), .b ({ciphertext_s3[74], ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .a ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, new_AGEMA_signal_2407, ShiftRowsOutput[42]}), .c ({new_AGEMA_signal_3618, new_AGEMA_signal_3617, new_AGEMA_signal_3616, RoundOutput[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_43_U1 ( .s (MuxRound_n15), .b ({ciphertext_s3[75], ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}), .a ({new_AGEMA_signal_2418, new_AGEMA_signal_2417, new_AGEMA_signal_2416, ShiftRowsOutput[43]}), .c ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, new_AGEMA_signal_3619, RoundOutput[43]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_44_U1 ( .s (MuxRound_n13), .b ({ciphertext_s3[76], ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .a ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, new_AGEMA_signal_2425, ShiftRowsOutput[44]}), .c ({new_AGEMA_signal_3624, new_AGEMA_signal_3623, new_AGEMA_signal_3622, RoundOutput[44]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_45_U1 ( .s (MuxRound_n14), .b ({ciphertext_s3[77], ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}), .a ({new_AGEMA_signal_2436, new_AGEMA_signal_2435, new_AGEMA_signal_2434, ShiftRowsOutput[45]}), .c ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, new_AGEMA_signal_3625, RoundOutput[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_46_U1 ( .s (MuxRound_n15), .b ({ciphertext_s3[78], ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}), .a ({new_AGEMA_signal_2454, new_AGEMA_signal_2453, new_AGEMA_signal_2452, ShiftRowsOutput[46]}), .c ({new_AGEMA_signal_3630, new_AGEMA_signal_3629, new_AGEMA_signal_3628, RoundOutput[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_47_U1 ( .s (MuxRound_n16), .b ({ciphertext_s3[79], ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .a ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, new_AGEMA_signal_2461, ShiftRowsOutput[47]}), .c ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, new_AGEMA_signal_3631, RoundOutput[47]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_48_U1 ( .s (MuxRound_n17), .b ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .a ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, new_AGEMA_signal_2659, ShiftRowsOutput[48]}), .c ({new_AGEMA_signal_3636, new_AGEMA_signal_3635, new_AGEMA_signal_3634, RoundOutput[48]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_49_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[113], ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .a ({new_AGEMA_signal_2670, new_AGEMA_signal_2669, new_AGEMA_signal_2668, ShiftRowsOutput[49]}), .c ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, new_AGEMA_signal_3637, RoundOutput[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_50_U1 ( .s (MuxRound_n13), .b ({ciphertext_s3[114], ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .a ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, new_AGEMA_signal_2677, ShiftRowsOutput[50]}), .c ({new_AGEMA_signal_3642, new_AGEMA_signal_3641, new_AGEMA_signal_3640, RoundOutput[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_51_U1 ( .s (MuxRound_n14), .b ({ciphertext_s3[115], ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}), .a ({new_AGEMA_signal_2688, new_AGEMA_signal_2687, new_AGEMA_signal_2686, ShiftRowsOutput[51]}), .c ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, new_AGEMA_signal_3643, RoundOutput[51]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_52_U1 ( .s (MuxRound_n15), .b ({ciphertext_s3[116], ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .a ({new_AGEMA_signal_2706, new_AGEMA_signal_2705, new_AGEMA_signal_2704, ShiftRowsOutput[52]}), .c ({new_AGEMA_signal_3648, new_AGEMA_signal_3647, new_AGEMA_signal_3646, RoundOutput[52]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_53_U1 ( .s (MuxRound_n16), .b ({ciphertext_s3[117], ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}), .a ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, new_AGEMA_signal_2713, ShiftRowsOutput[53]}), .c ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, new_AGEMA_signal_3649, RoundOutput[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_54_U1 ( .s (MuxRound_n17), .b ({ciphertext_s3[118], ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}), .a ({new_AGEMA_signal_2724, new_AGEMA_signal_2723, new_AGEMA_signal_2722, ShiftRowsOutput[54]}), .c ({new_AGEMA_signal_3654, new_AGEMA_signal_3653, new_AGEMA_signal_3652, RoundOutput[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_55_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[119], ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .a ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, new_AGEMA_signal_2731, ShiftRowsOutput[55]}), .c ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, new_AGEMA_signal_3655, RoundOutput[55]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_56_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .a ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, new_AGEMA_signal_3055, ShiftRowsOutput[56]}), .c ({new_AGEMA_signal_3660, new_AGEMA_signal_3659, new_AGEMA_signal_3658, RoundOutput[56]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_57_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .a ({new_AGEMA_signal_3066, new_AGEMA_signal_3065, new_AGEMA_signal_3064, ShiftRowsOutput[57]}), .c ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, new_AGEMA_signal_3661, RoundOutput[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_58_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .a ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, new_AGEMA_signal_3073, ShiftRowsOutput[58]}), .c ({new_AGEMA_signal_3666, new_AGEMA_signal_3665, new_AGEMA_signal_3664, RoundOutput[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_59_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .a ({new_AGEMA_signal_3084, new_AGEMA_signal_3083, new_AGEMA_signal_3082, ShiftRowsOutput[59]}), .c ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, new_AGEMA_signal_3667, RoundOutput[59]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_60_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .a ({new_AGEMA_signal_3102, new_AGEMA_signal_3101, new_AGEMA_signal_3100, ShiftRowsOutput[60]}), .c ({new_AGEMA_signal_3672, new_AGEMA_signal_3671, new_AGEMA_signal_3670, RoundOutput[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_61_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .a ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, new_AGEMA_signal_3109, ShiftRowsOutput[61]}), .c ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, new_AGEMA_signal_3673, RoundOutput[61]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_62_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .a ({new_AGEMA_signal_3120, new_AGEMA_signal_3119, new_AGEMA_signal_3118, ShiftRowsOutput[62]}), .c ({new_AGEMA_signal_3678, new_AGEMA_signal_3677, new_AGEMA_signal_3676, RoundOutput[62]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_63_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .a ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, new_AGEMA_signal_3127, ShiftRowsOutput[63]}), .c ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, new_AGEMA_signal_3679, RoundOutput[63]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_64_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .a ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, new_AGEMA_signal_3451, ShiftRowsOutput[64]}), .c ({new_AGEMA_signal_3684, new_AGEMA_signal_3683, new_AGEMA_signal_3682, RoundOutput[64]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_65_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[65], ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .a ({new_AGEMA_signal_3462, new_AGEMA_signal_3461, new_AGEMA_signal_3460, ShiftRowsOutput[65]}), .c ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, new_AGEMA_signal_3685, RoundOutput[65]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_66_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[66], ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .a ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, new_AGEMA_signal_3469, ShiftRowsOutput[66]}), .c ({new_AGEMA_signal_3690, new_AGEMA_signal_3689, new_AGEMA_signal_3688, RoundOutput[66]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_67_U1 ( .s (MuxRound_n18), .b ({ciphertext_s3[67], ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}), .a ({new_AGEMA_signal_3480, new_AGEMA_signal_3479, new_AGEMA_signal_3478, ShiftRowsOutput[67]}), .c ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, new_AGEMA_signal_3691, RoundOutput[67]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_68_U1 ( .s (MuxRound_n17), .b ({ciphertext_s3[68], ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .a ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, new_AGEMA_signal_2353, ShiftRowsOutput[68]}), .c ({new_AGEMA_signal_3696, new_AGEMA_signal_3695, new_AGEMA_signal_3694, RoundOutput[68]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_69_U1 ( .s (MuxRound_n17), .b ({ciphertext_s3[69], ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}), .a ({new_AGEMA_signal_2364, new_AGEMA_signal_2363, new_AGEMA_signal_2362, ShiftRowsOutput[69]}), .c ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, new_AGEMA_signal_3697, RoundOutput[69]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_70_U1 ( .s (MuxRound_n17), .b ({ciphertext_s3[70], ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}), .a ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, new_AGEMA_signal_2371, ShiftRowsOutput[70]}), .c ({new_AGEMA_signal_3702, new_AGEMA_signal_3701, new_AGEMA_signal_3700, RoundOutput[70]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_71_U1 ( .s (MuxRound_n17), .b ({ciphertext_s3[71], ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .a ({new_AGEMA_signal_2382, new_AGEMA_signal_2381, new_AGEMA_signal_2380, ShiftRowsOutput[71]}), .c ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, new_AGEMA_signal_3703, RoundOutput[71]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_72_U1 ( .s (MuxRound_n17), .b ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .a ({new_AGEMA_signal_3390, new_AGEMA_signal_3389, new_AGEMA_signal_3388, ShiftRowsOutput[72]}), .c ({new_AGEMA_signal_3708, new_AGEMA_signal_3707, new_AGEMA_signal_3706, RoundOutput[72]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_73_U1 ( .s (MuxRound_n17), .b ({ciphertext_s3[105], ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .a ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, new_AGEMA_signal_3487, ShiftRowsOutput[73]}), .c ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, new_AGEMA_signal_3709, RoundOutput[73]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_74_U1 ( .s (MuxRound_n17), .b ({ciphertext_s3[106], ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .a ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, new_AGEMA_signal_2443, ShiftRowsOutput[74]}), .c ({new_AGEMA_signal_3714, new_AGEMA_signal_3713, new_AGEMA_signal_3712, RoundOutput[74]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_75_U1 ( .s (MuxRound_n17), .b ({ciphertext_s3[107], ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}), .a ({new_AGEMA_signal_2544, new_AGEMA_signal_2543, new_AGEMA_signal_2542, ShiftRowsOutput[75]}), .c ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, new_AGEMA_signal_3715, RoundOutput[75]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_76_U1 ( .s (MuxRound_n17), .b ({ciphertext_s3[108], ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .a ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, new_AGEMA_signal_2623, ShiftRowsOutput[76]}), .c ({new_AGEMA_signal_3720, new_AGEMA_signal_3719, new_AGEMA_signal_3718, RoundOutput[76]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_77_U1 ( .s (MuxRound_n17), .b ({ciphertext_s3[109], ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}), .a ({new_AGEMA_signal_2634, new_AGEMA_signal_2633, new_AGEMA_signal_2632, ShiftRowsOutput[77]}), .c ({new_AGEMA_signal_3723, new_AGEMA_signal_3722, new_AGEMA_signal_3721, RoundOutput[77]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_78_U1 ( .s (MuxRound_n17), .b ({ciphertext_s3[110], ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}), .a ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, new_AGEMA_signal_2641, ShiftRowsOutput[78]}), .c ({new_AGEMA_signal_3726, new_AGEMA_signal_3725, new_AGEMA_signal_3724, RoundOutput[78]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_79_U1 ( .s (MuxRound_n17), .b ({ciphertext_s3[111], ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .a ({new_AGEMA_signal_2652, new_AGEMA_signal_2651, new_AGEMA_signal_2650, ShiftRowsOutput[79]}), .c ({new_AGEMA_signal_3729, new_AGEMA_signal_3728, new_AGEMA_signal_3727, RoundOutput[79]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_80_U1 ( .s (MuxRound_n16), .b ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .a ({new_AGEMA_signal_2976, new_AGEMA_signal_2975, new_AGEMA_signal_2974, ShiftRowsOutput[80]}), .c ({new_AGEMA_signal_3732, new_AGEMA_signal_3731, new_AGEMA_signal_3730, RoundOutput[80]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_81_U1 ( .s (MuxRound_n16), .b ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .a ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, new_AGEMA_signal_2983, ShiftRowsOutput[81]}), .c ({new_AGEMA_signal_3735, new_AGEMA_signal_3734, new_AGEMA_signal_3733, RoundOutput[81]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_82_U1 ( .s (MuxRound_n16), .b ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .a ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, new_AGEMA_signal_3001, ShiftRowsOutput[82]}), .c ({new_AGEMA_signal_3738, new_AGEMA_signal_3737, new_AGEMA_signal_3736, RoundOutput[82]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_83_U1 ( .s (MuxRound_n16), .b ({ciphertext_s3[19], ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .a ({new_AGEMA_signal_3012, new_AGEMA_signal_3011, new_AGEMA_signal_3010, ShiftRowsOutput[83]}), .c ({new_AGEMA_signal_3741, new_AGEMA_signal_3740, new_AGEMA_signal_3739, RoundOutput[83]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_84_U1 ( .s (MuxRound_n16), .b ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .a ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, new_AGEMA_signal_3019, ShiftRowsOutput[84]}), .c ({new_AGEMA_signal_3744, new_AGEMA_signal_3743, new_AGEMA_signal_3742, RoundOutput[84]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_85_U1 ( .s (MuxRound_n16), .b ({ciphertext_s3[21], ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .a ({new_AGEMA_signal_3030, new_AGEMA_signal_3029, new_AGEMA_signal_3028, ShiftRowsOutput[85]}), .c ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, new_AGEMA_signal_3745, RoundOutput[85]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_86_U1 ( .s (MuxRound_n16), .b ({ciphertext_s3[22], ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .a ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, new_AGEMA_signal_3037, ShiftRowsOutput[86]}), .c ({new_AGEMA_signal_3750, new_AGEMA_signal_3749, new_AGEMA_signal_3748, RoundOutput[86]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_87_U1 ( .s (MuxRound_n16), .b ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .a ({new_AGEMA_signal_3048, new_AGEMA_signal_3047, new_AGEMA_signal_3046, ShiftRowsOutput[87]}), .c ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, new_AGEMA_signal_3751, RoundOutput[87]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_88_U1 ( .s (MuxRound_n16), .b ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .a ({new_AGEMA_signal_3372, new_AGEMA_signal_3371, new_AGEMA_signal_3370, ShiftRowsOutput[88]}), .c ({new_AGEMA_signal_3756, new_AGEMA_signal_3755, new_AGEMA_signal_3754, RoundOutput[88]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_89_U1 ( .s (MuxRound_n16), .b ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .a ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, new_AGEMA_signal_3379, ShiftRowsOutput[89]}), .c ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, new_AGEMA_signal_3757, RoundOutput[89]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_90_U1 ( .s (MuxRound_n16), .b ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .a ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, new_AGEMA_signal_3397, ShiftRowsOutput[90]}), .c ({new_AGEMA_signal_3762, new_AGEMA_signal_3761, new_AGEMA_signal_3760, RoundOutput[90]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_91_U1 ( .s (MuxRound_n16), .b ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .a ({new_AGEMA_signal_3408, new_AGEMA_signal_3407, new_AGEMA_signal_3406, ShiftRowsOutput[91]}), .c ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, new_AGEMA_signal_3763, RoundOutput[91]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_92_U1 ( .s (MuxRound_n15), .b ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .a ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, new_AGEMA_signal_3415, ShiftRowsOutput[92]}), .c ({new_AGEMA_signal_3768, new_AGEMA_signal_3767, new_AGEMA_signal_3766, RoundOutput[92]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_93_U1 ( .s (MuxRound_n15), .b ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .a ({new_AGEMA_signal_3426, new_AGEMA_signal_3425, new_AGEMA_signal_3424, ShiftRowsOutput[93]}), .c ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, new_AGEMA_signal_3769, RoundOutput[93]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_94_U1 ( .s (MuxRound_n15), .b ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .a ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, new_AGEMA_signal_3433, ShiftRowsOutput[94]}), .c ({new_AGEMA_signal_3774, new_AGEMA_signal_3773, new_AGEMA_signal_3772, RoundOutput[94]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_95_U1 ( .s (MuxRound_n15), .b ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .a ({new_AGEMA_signal_3444, new_AGEMA_signal_3443, new_AGEMA_signal_3442, ShiftRowsOutput[95]}), .c ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, new_AGEMA_signal_3775, RoundOutput[95]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_96_U1 ( .s (MuxRound_n15), .b ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .a ({new_AGEMA_signal_2346, new_AGEMA_signal_2345, new_AGEMA_signal_2344, ShiftRowsOutput[96]}), .c ({new_AGEMA_signal_3780, new_AGEMA_signal_3779, new_AGEMA_signal_3778, RoundOutput[96]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_97_U1 ( .s (MuxRound_n15), .b ({ciphertext_s3[97], ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .a ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, new_AGEMA_signal_2695, ShiftRowsOutput[97]}), .c ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, new_AGEMA_signal_3781, RoundOutput[97]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_98_U1 ( .s (MuxRound_n15), .b ({ciphertext_s3[98], ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .a ({new_AGEMA_signal_2796, new_AGEMA_signal_2795, new_AGEMA_signal_2794, ShiftRowsOutput[98]}), .c ({new_AGEMA_signal_3786, new_AGEMA_signal_3785, new_AGEMA_signal_3784, RoundOutput[98]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_99_U1 ( .s (MuxRound_n15), .b ({ciphertext_s3[99], ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}), .a ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, new_AGEMA_signal_2893, ShiftRowsOutput[99]}), .c ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, new_AGEMA_signal_3787, RoundOutput[99]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_100_U1 ( .s (MuxRound_n15), .b ({ciphertext_s3[100], ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .a ({new_AGEMA_signal_2994, new_AGEMA_signal_2993, new_AGEMA_signal_2992, ShiftRowsOutput[100]}), .c ({new_AGEMA_signal_3792, new_AGEMA_signal_3791, new_AGEMA_signal_3790, RoundOutput[100]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_101_U1 ( .s (MuxRound_n15), .b ({ciphertext_s3[101], ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}), .a ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, new_AGEMA_signal_3091, ShiftRowsOutput[101]}), .c ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, new_AGEMA_signal_3793, RoundOutput[101]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_102_U1 ( .s (MuxRound_n15), .b ({ciphertext_s3[102], ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}), .a ({new_AGEMA_signal_3192, new_AGEMA_signal_3191, new_AGEMA_signal_3190, ShiftRowsOutput[102]}), .c ({new_AGEMA_signal_3798, new_AGEMA_signal_3797, new_AGEMA_signal_3796, RoundOutput[102]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_103_U1 ( .s (MuxRound_n15), .b ({ciphertext_s3[103], ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .a ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, new_AGEMA_signal_3289, ShiftRowsOutput[103]}), .c ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, new_AGEMA_signal_3799, RoundOutput[103]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_104_U1 ( .s (MuxRound_n14), .b ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .a ({new_AGEMA_signal_2904, new_AGEMA_signal_2903, new_AGEMA_signal_2902, ShiftRowsOutput[104]}), .c ({new_AGEMA_signal_3804, new_AGEMA_signal_3803, new_AGEMA_signal_3802, RoundOutput[104]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_105_U1 ( .s (MuxRound_n14), .b ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .a ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, new_AGEMA_signal_2911, ShiftRowsOutput[105]}), .c ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, new_AGEMA_signal_3805, RoundOutput[105]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_106_U1 ( .s (MuxRound_n14), .b ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .a ({new_AGEMA_signal_2922, new_AGEMA_signal_2921, new_AGEMA_signal_2920, ShiftRowsOutput[106]}), .c ({new_AGEMA_signal_3810, new_AGEMA_signal_3809, new_AGEMA_signal_3808, RoundOutput[106]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_107_U1 ( .s (MuxRound_n14), .b ({ciphertext_s3[11], ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .a ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, new_AGEMA_signal_2929, ShiftRowsOutput[107]}), .c ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, new_AGEMA_signal_3811, RoundOutput[107]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_108_U1 ( .s (MuxRound_n14), .b ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .a ({new_AGEMA_signal_2940, new_AGEMA_signal_2939, new_AGEMA_signal_2938, ShiftRowsOutput[108]}), .c ({new_AGEMA_signal_3816, new_AGEMA_signal_3815, new_AGEMA_signal_3814, RoundOutput[108]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_109_U1 ( .s (MuxRound_n14), .b ({ciphertext_s3[13], ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .a ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, new_AGEMA_signal_2947, ShiftRowsOutput[109]}), .c ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, new_AGEMA_signal_3817, RoundOutput[109]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_110_U1 ( .s (MuxRound_n14), .b ({ciphertext_s3[14], ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .a ({new_AGEMA_signal_2958, new_AGEMA_signal_2957, new_AGEMA_signal_2956, ShiftRowsOutput[110]}), .c ({new_AGEMA_signal_3822, new_AGEMA_signal_3821, new_AGEMA_signal_3820, RoundOutput[110]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_111_U1 ( .s (MuxRound_n14), .b ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .a ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, new_AGEMA_signal_2965, ShiftRowsOutput[111]}), .c ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, new_AGEMA_signal_3823, RoundOutput[111]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_112_U1 ( .s (MuxRound_n14), .b ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .a ({new_AGEMA_signal_3300, new_AGEMA_signal_3299, new_AGEMA_signal_3298, ShiftRowsOutput[112]}), .c ({new_AGEMA_signal_3828, new_AGEMA_signal_3827, new_AGEMA_signal_3826, RoundOutput[112]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_113_U1 ( .s (MuxRound_n14), .b ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .a ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, new_AGEMA_signal_3307, ShiftRowsOutput[113]}), .c ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, new_AGEMA_signal_3829, RoundOutput[113]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_114_U1 ( .s (MuxRound_n14), .b ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .a ({new_AGEMA_signal_3318, new_AGEMA_signal_3317, new_AGEMA_signal_3316, ShiftRowsOutput[114]}), .c ({new_AGEMA_signal_3834, new_AGEMA_signal_3833, new_AGEMA_signal_3832, RoundOutput[114]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_115_U1 ( .s (MuxRound_n14), .b ({ciphertext_s3[51], ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .a ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, new_AGEMA_signal_3325, ShiftRowsOutput[115]}), .c ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, new_AGEMA_signal_3835, RoundOutput[115]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_116_U1 ( .s (MuxRound_n13), .b ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .a ({new_AGEMA_signal_3336, new_AGEMA_signal_3335, new_AGEMA_signal_3334, ShiftRowsOutput[116]}), .c ({new_AGEMA_signal_3840, new_AGEMA_signal_3839, new_AGEMA_signal_3838, RoundOutput[116]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_117_U1 ( .s (MuxRound_n13), .b ({ciphertext_s3[53], ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .a ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, new_AGEMA_signal_3343, ShiftRowsOutput[117]}), .c ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, new_AGEMA_signal_3841, RoundOutput[117]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_118_U1 ( .s (MuxRound_n13), .b ({ciphertext_s3[54], ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .a ({new_AGEMA_signal_3354, new_AGEMA_signal_3353, new_AGEMA_signal_3352, ShiftRowsOutput[118]}), .c ({new_AGEMA_signal_3846, new_AGEMA_signal_3845, new_AGEMA_signal_3844, RoundOutput[118]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_119_U1 ( .s (MuxRound_n13), .b ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .a ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, new_AGEMA_signal_3361, ShiftRowsOutput[119]}), .c ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, new_AGEMA_signal_3847, RoundOutput[119]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_120_U1 ( .s (MuxRound_n13), .b ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .a ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, new_AGEMA_signal_2551, ShiftRowsOutput[120]}), .c ({new_AGEMA_signal_3852, new_AGEMA_signal_3851, new_AGEMA_signal_3850, RoundOutput[120]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_121_U1 ( .s (MuxRound_n13), .b ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .a ({new_AGEMA_signal_2562, new_AGEMA_signal_2561, new_AGEMA_signal_2560, ShiftRowsOutput[121]}), .c ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, new_AGEMA_signal_3853, RoundOutput[121]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_122_U1 ( .s (MuxRound_n13), .b ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .a ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, new_AGEMA_signal_2569, ShiftRowsOutput[122]}), .c ({new_AGEMA_signal_3858, new_AGEMA_signal_3857, new_AGEMA_signal_3856, RoundOutput[122]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_123_U1 ( .s (MuxRound_n13), .b ({ciphertext_s3[91], ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .a ({new_AGEMA_signal_2580, new_AGEMA_signal_2579, new_AGEMA_signal_2578, ShiftRowsOutput[123]}), .c ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, new_AGEMA_signal_3859, RoundOutput[123]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_124_U1 ( .s (MuxRound_n13), .b ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .a ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, new_AGEMA_signal_2587, ShiftRowsOutput[124]}), .c ({new_AGEMA_signal_3864, new_AGEMA_signal_3863, new_AGEMA_signal_3862, RoundOutput[124]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_125_U1 ( .s (MuxRound_n13), .b ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .a ({new_AGEMA_signal_2598, new_AGEMA_signal_2597, new_AGEMA_signal_2596, ShiftRowsOutput[125]}), .c ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, new_AGEMA_signal_3865, RoundOutput[125]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_126_U1 ( .s (MuxRound_n13), .b ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .a ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, new_AGEMA_signal_2605, ShiftRowsOutput[126]}), .c ({new_AGEMA_signal_3870, new_AGEMA_signal_3869, new_AGEMA_signal_3868, RoundOutput[126]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_127_U1 ( .s (MuxRound_n13), .b ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .a ({new_AGEMA_signal_2616, new_AGEMA_signal_2615, new_AGEMA_signal_2614, ShiftRowsOutput[127]}), .c ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, new_AGEMA_signal_3871, RoundOutput[127]}) ) ;
    INV_X1 MuxKeyExpansion_U8 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n14) ) ;
    INV_X1 MuxKeyExpansion_U7 ( .A (AKSRnotDone), .ZN (MuxKeyExpansion_n21) ) ;
    INV_X1 MuxKeyExpansion_U6 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n16) ) ;
    INV_X1 MuxKeyExpansion_U5 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n17) ) ;
    INV_X1 MuxKeyExpansion_U4 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n18) ) ;
    INV_X1 MuxKeyExpansion_U3 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n19) ) ;
    INV_X1 MuxKeyExpansion_U2 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n20) ) ;
    INV_X1 MuxKeyExpansion_U1 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n15) ) ;
    NOR2_X1 RoundCounterIns_U11 ( .A1 (reset), .A2 (RoundCounterIns_n10), .ZN (RoundCounterIns_n45) ) ;
    XNOR2_X1 RoundCounterIns_U10 ( .A (RoundCounter[0]), .B (AKSRnotDone), .ZN (RoundCounterIns_n10) ) ;
    NOR2_X1 RoundCounterIns_U9 ( .A1 (reset), .A2 (RoundCounterIns_n9), .ZN (RoundCounterIns_n44) ) ;
    XOR2_X1 RoundCounterIns_U8 ( .A (RoundCounter[1]), .B (RoundCounterIns_n8), .Z (RoundCounterIns_n9) ) ;
    NOR2_X1 RoundCounterIns_U7 ( .A1 (reset), .A2 (RoundCounterIns_n7), .ZN (RoundCounterIns_n42) ) ;
    XOR2_X1 RoundCounterIns_U6 ( .A (RoundCounter[3]), .B (RoundCounterIns_n6), .Z (RoundCounterIns_n7) ) ;
    NAND2_X1 RoundCounterIns_U5 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounter[2]), .ZN (RoundCounterIns_n6) ) ;
    NOR2_X1 RoundCounterIns_U4 ( .A1 (reset), .A2 (RoundCounterIns_n4), .ZN (RoundCounterIns_n1) ) ;
    XNOR2_X1 RoundCounterIns_U3 ( .A (RoundCounter[2]), .B (RoundCounterIns_n5), .ZN (RoundCounterIns_n4) ) ;
    NOR2_X1 RoundCounterIns_U2 ( .A1 (RoundCounterIns_n2), .A2 (RoundCounterIns_n8), .ZN (RoundCounterIns_n5) ) ;
    NAND2_X1 RoundCounterIns_U1 ( .A1 (AKSRnotDone), .A2 (RoundCounter[0]), .ZN (RoundCounterIns_n8) ) ;
    INV_X1 RoundCounterIns_count_reg_1__U1 ( .A (RoundCounter[1]), .ZN (RoundCounterIns_n2) ) ;
    NOR2_X1 InRoundCounterIns_U13 ( .A1 (reset), .A2 (InRoundCounterIns_n12), .ZN (InRoundCounterIns_n41) ) ;
    XOR2_X1 InRoundCounterIns_U12 ( .A (InRoundCounter[0]), .B (InRoundCounterIns_n11), .Z (InRoundCounterIns_n12) ) ;
    NAND2_X1 InRoundCounterIns_U11 ( .A1 (InRoundCounterIns_n10), .A2 (1'b1), .ZN (InRoundCounterIns_n11) ) ;
    NAND2_X1 InRoundCounterIns_U10 ( .A1 (InRoundCounterIns_n9), .A2 (InRoundCounter[2]), .ZN (InRoundCounterIns_n10) ) ;
    NAND2_X1 InRoundCounterIns_U9 ( .A1 (InRoundCounter[0]), .A2 (InRoundCounter[1]), .ZN (InRoundCounterIns_n9) ) ;
    NOR2_X1 InRoundCounterIns_U8 ( .A1 (reset), .A2 (InRoundCounterIns_n8), .ZN (InRoundCounterIns_n40) ) ;
    MUX2_X1 InRoundCounterIns_U7 ( .S (InRoundCounter[1]), .A (InRoundCounterIns_n7), .B (InRoundCounterIns_n5), .Z (InRoundCounterIns_n8) ) ;
    NOR2_X1 InRoundCounterIns_U6 ( .A1 (reset), .A2 (InRoundCounterIns_n4), .ZN (InRoundCounterIns_n39) ) ;
    NOR2_X1 InRoundCounterIns_U5 ( .A1 (InRoundCounterIns_n3), .A2 (InRoundCounterIns_n2), .ZN (InRoundCounterIns_n4) ) ;
    NOR2_X1 InRoundCounterIns_U4 ( .A1 (InRoundCounterIns_n1), .A2 (InRoundCounterIns_n7), .ZN (InRoundCounterIns_n2) ) ;
    NAND2_X1 InRoundCounterIns_U3 ( .A1 (InRoundCounterIns_n5), .A2 (InRoundCounterIns_n6), .ZN (InRoundCounterIns_n7) ) ;
    AND2_X1 InRoundCounterIns_U2 ( .A1 (InRoundCounter[0]), .A2 (1'b1), .ZN (InRoundCounterIns_n5) ) ;
    NOR2_X1 InRoundCounterIns_U1 ( .A1 (1'b1), .A2 (InRoundCounterIns_n6), .ZN (InRoundCounterIns_n3) ) ;
    INV_X1 InRoundCounterIns_count_reg_1__U1 ( .A (InRoundCounter[1]), .ZN (InRoundCounterIns_n1) ) ;
    INV_X1 InRoundCounterIns_count_reg_2__U1 ( .A (InRoundCounter[2]), .ZN (InRoundCounterIns_n6) ) ;

    /* cells in depth 1 */
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_4578, new_AGEMA_signal_4577, new_AGEMA_signal_4576, SubBytesIns_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_4572, new_AGEMA_signal_4571, new_AGEMA_signal_4570, SubBytesIns_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_4689, new_AGEMA_signal_4688, new_AGEMA_signal_4687, SubBytesIns_Inst_Sbox_0_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_4683, new_AGEMA_signal_4682, new_AGEMA_signal_4681, SubBytesIns_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_4668, new_AGEMA_signal_4667, new_AGEMA_signal_4666, SubBytesIns_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_4830, new_AGEMA_signal_4829, new_AGEMA_signal_4828, SubBytesIns_Inst_Sbox_0_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_9889, new_AGEMA_signal_9888, new_AGEMA_signal_9887, new_AGEMA_signal_9886}), .b ({new_AGEMA_signal_4689, new_AGEMA_signal_4688, new_AGEMA_signal_4687, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, new_AGEMA_signal_4831, SubBytesIns_Inst_Sbox_0_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_4587, new_AGEMA_signal_4586, new_AGEMA_signal_4585, SubBytesIns_Inst_Sbox_0_T19}), .b ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, new_AGEMA_signal_3493, SubBytesInput[0]}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_4692, new_AGEMA_signal_4691, new_AGEMA_signal_4690, SubBytesIns_Inst_Sbox_0_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_4692, new_AGEMA_signal_4691, new_AGEMA_signal_4690, SubBytesIns_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_4689, new_AGEMA_signal_4688, new_AGEMA_signal_4687, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_4836, new_AGEMA_signal_4835, new_AGEMA_signal_4834, SubBytesIns_Inst_Sbox_0_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_4458, new_AGEMA_signal_4457, new_AGEMA_signal_4456, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_4584, new_AGEMA_signal_4583, new_AGEMA_signal_4582, SubBytesIns_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_4695, new_AGEMA_signal_4694, new_AGEMA_signal_4693, SubBytesIns_Inst_Sbox_0_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_4590, new_AGEMA_signal_4589, new_AGEMA_signal_4588, SubBytesIns_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, new_AGEMA_signal_4573, SubBytesIns_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_4698, new_AGEMA_signal_4697, new_AGEMA_signal_4696, SubBytesIns_Inst_Sbox_0_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_9893, new_AGEMA_signal_9892, new_AGEMA_signal_9891, new_AGEMA_signal_9890}), .b ({new_AGEMA_signal_4695, new_AGEMA_signal_4694, new_AGEMA_signal_4693, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_4839, new_AGEMA_signal_4838, new_AGEMA_signal_4837, SubBytesIns_Inst_Sbox_0_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_4680, new_AGEMA_signal_4679, new_AGEMA_signal_4678, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_4677, new_AGEMA_signal_4676, new_AGEMA_signal_4675, SubBytesIns_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_4842, new_AGEMA_signal_4841, new_AGEMA_signal_4840, SubBytesIns_Inst_Sbox_0_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_4842, new_AGEMA_signal_4841, new_AGEMA_signal_4840, SubBytesIns_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_4695, new_AGEMA_signal_4694, new_AGEMA_signal_4693, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_4932, new_AGEMA_signal_4931, new_AGEMA_signal_4930, SubBytesIns_Inst_Sbox_0_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_4452, new_AGEMA_signal_4451, new_AGEMA_signal_4450, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, new_AGEMA_signal_4579, SubBytesIns_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_4701, new_AGEMA_signal_4700, new_AGEMA_signal_4699, SubBytesIns_Inst_Sbox_0_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_4461, new_AGEMA_signal_4460, new_AGEMA_signal_4459, SubBytesIns_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, new_AGEMA_signal_4591, SubBytesIns_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90], Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_4704, new_AGEMA_signal_4703, new_AGEMA_signal_4702, SubBytesIns_Inst_Sbox_0_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_4704, new_AGEMA_signal_4703, new_AGEMA_signal_4702, SubBytesIns_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_4701, new_AGEMA_signal_4700, new_AGEMA_signal_4699, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_4845, new_AGEMA_signal_4844, new_AGEMA_signal_4843, SubBytesIns_Inst_Sbox_0_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_4455, new_AGEMA_signal_4454, new_AGEMA_signal_4453, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, new_AGEMA_signal_4669, SubBytesIns_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_4848, new_AGEMA_signal_4847, new_AGEMA_signal_4846, SubBytesIns_Inst_Sbox_0_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_4848, new_AGEMA_signal_4847, new_AGEMA_signal_4846, SubBytesIns_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_4701, new_AGEMA_signal_4700, new_AGEMA_signal_4699, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_4935, new_AGEMA_signal_4934, new_AGEMA_signal_4933, SubBytesIns_Inst_Sbox_0_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, new_AGEMA_signal_4831, SubBytesIns_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_4830, new_AGEMA_signal_4829, new_AGEMA_signal_4828, SubBytesIns_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_4938, new_AGEMA_signal_4937, new_AGEMA_signal_4936, SubBytesIns_Inst_Sbox_0_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_4836, new_AGEMA_signal_4835, new_AGEMA_signal_4834, SubBytesIns_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_9897, new_AGEMA_signal_9896, new_AGEMA_signal_9895, new_AGEMA_signal_9894}), .c ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, new_AGEMA_signal_4939, SubBytesIns_Inst_Sbox_0_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_4839, new_AGEMA_signal_4838, new_AGEMA_signal_4837, SubBytesIns_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_4698, new_AGEMA_signal_4697, new_AGEMA_signal_4696, SubBytesIns_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_4944, new_AGEMA_signal_4943, new_AGEMA_signal_4942, SubBytesIns_Inst_Sbox_0_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_4932, new_AGEMA_signal_4931, new_AGEMA_signal_4930, SubBytesIns_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_4935, new_AGEMA_signal_4934, new_AGEMA_signal_4933, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_4992, new_AGEMA_signal_4991, new_AGEMA_signal_4990, SubBytesIns_Inst_Sbox_0_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_4938, new_AGEMA_signal_4937, new_AGEMA_signal_4936, SubBytesIns_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_4845, new_AGEMA_signal_4844, new_AGEMA_signal_4843, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, new_AGEMA_signal_4993, SubBytesIns_Inst_Sbox_0_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, new_AGEMA_signal_4939, SubBytesIns_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_4935, new_AGEMA_signal_4934, new_AGEMA_signal_4933, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_4998, new_AGEMA_signal_4997, new_AGEMA_signal_4996, SubBytesIns_Inst_Sbox_0_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_4944, new_AGEMA_signal_4943, new_AGEMA_signal_4942, SubBytesIns_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_4845, new_AGEMA_signal_4844, new_AGEMA_signal_4843, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, new_AGEMA_signal_4999, SubBytesIns_Inst_Sbox_0_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_4992, new_AGEMA_signal_4991, new_AGEMA_signal_4990, SubBytesIns_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_9901, new_AGEMA_signal_9900, new_AGEMA_signal_9899, new_AGEMA_signal_9898}), .c ({new_AGEMA_signal_5040, new_AGEMA_signal_5039, new_AGEMA_signal_5038, SubBytesIns_Inst_Sbox_0_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, new_AGEMA_signal_4999, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_5040, new_AGEMA_signal_5039, new_AGEMA_signal_5038, SubBytesIns_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_5088, new_AGEMA_signal_5087, new_AGEMA_signal_5086, SubBytesIns_Inst_Sbox_0_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, new_AGEMA_signal_4993, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_4998, new_AGEMA_signal_4997, new_AGEMA_signal_4996, SubBytesIns_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_5046, new_AGEMA_signal_5045, new_AGEMA_signal_5044, SubBytesIns_Inst_Sbox_0_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_4602, new_AGEMA_signal_4601, new_AGEMA_signal_4600, SubBytesIns_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_4596, new_AGEMA_signal_4595, new_AGEMA_signal_4594, SubBytesIns_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_4728, new_AGEMA_signal_4727, new_AGEMA_signal_4726, SubBytesIns_Inst_Sbox_1_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_4722, new_AGEMA_signal_4721, new_AGEMA_signal_4720, SubBytesIns_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_4707, new_AGEMA_signal_4706, new_AGEMA_signal_4705, SubBytesIns_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_4857, new_AGEMA_signal_4856, new_AGEMA_signal_4855, SubBytesIns_Inst_Sbox_1_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_9905, new_AGEMA_signal_9904, new_AGEMA_signal_9903, new_AGEMA_signal_9902}), .b ({new_AGEMA_signal_4728, new_AGEMA_signal_4727, new_AGEMA_signal_4726, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, new_AGEMA_signal_4858, SubBytesIns_Inst_Sbox_1_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_4611, new_AGEMA_signal_4610, new_AGEMA_signal_4609, SubBytesIns_Inst_Sbox_1_T19}), .b ({new_AGEMA_signal_3492, new_AGEMA_signal_3491, new_AGEMA_signal_3490, SubBytesInput[8]}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, new_AGEMA_signal_4729, SubBytesIns_Inst_Sbox_1_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, new_AGEMA_signal_4729, SubBytesIns_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_4728, new_AGEMA_signal_4727, new_AGEMA_signal_4726, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_4863, new_AGEMA_signal_4862, new_AGEMA_signal_4861, SubBytesIns_Inst_Sbox_1_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_4488, new_AGEMA_signal_4487, new_AGEMA_signal_4486, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_4608, new_AGEMA_signal_4607, new_AGEMA_signal_4606, SubBytesIns_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150], Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_4734, new_AGEMA_signal_4733, new_AGEMA_signal_4732, SubBytesIns_Inst_Sbox_1_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_4614, new_AGEMA_signal_4613, new_AGEMA_signal_4612, SubBytesIns_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, new_AGEMA_signal_4597, SubBytesIns_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, new_AGEMA_signal_4735, SubBytesIns_Inst_Sbox_1_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_9909, new_AGEMA_signal_9908, new_AGEMA_signal_9907, new_AGEMA_signal_9906}), .b ({new_AGEMA_signal_4734, new_AGEMA_signal_4733, new_AGEMA_signal_4732, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_4866, new_AGEMA_signal_4865, new_AGEMA_signal_4864, SubBytesIns_Inst_Sbox_1_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, new_AGEMA_signal_4717, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_4716, new_AGEMA_signal_4715, new_AGEMA_signal_4714, SubBytesIns_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, SubBytesIns_Inst_Sbox_1_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, SubBytesIns_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_4734, new_AGEMA_signal_4733, new_AGEMA_signal_4732, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, new_AGEMA_signal_4945, SubBytesIns_Inst_Sbox_1_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_4482, new_AGEMA_signal_4481, new_AGEMA_signal_4480, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_4605, new_AGEMA_signal_4604, new_AGEMA_signal_4603, SubBytesIns_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_4740, new_AGEMA_signal_4739, new_AGEMA_signal_4738, SubBytesIns_Inst_Sbox_1_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_4491, new_AGEMA_signal_4490, new_AGEMA_signal_4489, SubBytesIns_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, new_AGEMA_signal_4615, SubBytesIns_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, new_AGEMA_signal_4741, SubBytesIns_Inst_Sbox_1_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, new_AGEMA_signal_4741, SubBytesIns_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_4740, new_AGEMA_signal_4739, new_AGEMA_signal_4738, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_4872, new_AGEMA_signal_4871, new_AGEMA_signal_4870, SubBytesIns_Inst_Sbox_1_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_4485, new_AGEMA_signal_4484, new_AGEMA_signal_4483, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_4710, new_AGEMA_signal_4709, new_AGEMA_signal_4708, SubBytesIns_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210], Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_4875, new_AGEMA_signal_4874, new_AGEMA_signal_4873, SubBytesIns_Inst_Sbox_1_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_4875, new_AGEMA_signal_4874, new_AGEMA_signal_4873, SubBytesIns_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_4740, new_AGEMA_signal_4739, new_AGEMA_signal_4738, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, SubBytesIns_Inst_Sbox_1_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, new_AGEMA_signal_4858, SubBytesIns_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_4857, new_AGEMA_signal_4856, new_AGEMA_signal_4855, SubBytesIns_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_4953, new_AGEMA_signal_4952, new_AGEMA_signal_4951, SubBytesIns_Inst_Sbox_1_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_4863, new_AGEMA_signal_4862, new_AGEMA_signal_4861, SubBytesIns_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_9913, new_AGEMA_signal_9912, new_AGEMA_signal_9911, new_AGEMA_signal_9910}), .c ({new_AGEMA_signal_4956, new_AGEMA_signal_4955, new_AGEMA_signal_4954, SubBytesIns_Inst_Sbox_1_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_4866, new_AGEMA_signal_4865, new_AGEMA_signal_4864, SubBytesIns_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, new_AGEMA_signal_4735, SubBytesIns_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, new_AGEMA_signal_4957, SubBytesIns_Inst_Sbox_1_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, new_AGEMA_signal_4945, SubBytesIns_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, SubBytesIns_Inst_Sbox_1_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_4953, new_AGEMA_signal_4952, new_AGEMA_signal_4951, SubBytesIns_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_4872, new_AGEMA_signal_4871, new_AGEMA_signal_4870, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_5007, new_AGEMA_signal_5006, new_AGEMA_signal_5005, SubBytesIns_Inst_Sbox_1_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_4956, new_AGEMA_signal_4955, new_AGEMA_signal_4954, SubBytesIns_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_5010, new_AGEMA_signal_5009, new_AGEMA_signal_5008, SubBytesIns_Inst_Sbox_1_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, new_AGEMA_signal_4957, SubBytesIns_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_4872, new_AGEMA_signal_4871, new_AGEMA_signal_4870, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, new_AGEMA_signal_5011, SubBytesIns_Inst_Sbox_1_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, SubBytesIns_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_9917, new_AGEMA_signal_9916, new_AGEMA_signal_9915, new_AGEMA_signal_9914}), .c ({new_AGEMA_signal_5052, new_AGEMA_signal_5051, new_AGEMA_signal_5050, SubBytesIns_Inst_Sbox_1_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, new_AGEMA_signal_5011, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_5052, new_AGEMA_signal_5051, new_AGEMA_signal_5050, SubBytesIns_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_5103, new_AGEMA_signal_5102, new_AGEMA_signal_5101, SubBytesIns_Inst_Sbox_1_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_5007, new_AGEMA_signal_5006, new_AGEMA_signal_5005, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_5010, new_AGEMA_signal_5009, new_AGEMA_signal_5008, SubBytesIns_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_5058, new_AGEMA_signal_5057, new_AGEMA_signal_5056, SubBytesIns_Inst_Sbox_1_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_4626, new_AGEMA_signal_4625, new_AGEMA_signal_4624, SubBytesIns_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_4620, new_AGEMA_signal_4619, new_AGEMA_signal_4618, SubBytesIns_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, new_AGEMA_signal_4765, SubBytesIns_Inst_Sbox_2_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, new_AGEMA_signal_4759, SubBytesIns_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_4746, new_AGEMA_signal_4745, new_AGEMA_signal_4744, SubBytesIns_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_4884, new_AGEMA_signal_4883, new_AGEMA_signal_4882, SubBytesIns_Inst_Sbox_2_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_9921, new_AGEMA_signal_9920, new_AGEMA_signal_9919, new_AGEMA_signal_9918}), .b ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, new_AGEMA_signal_4765, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, SubBytesIns_Inst_Sbox_2_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_4635, new_AGEMA_signal_4634, new_AGEMA_signal_4633, SubBytesIns_Inst_Sbox_2_T19}), .b ({new_AGEMA_signal_3540, new_AGEMA_signal_3539, new_AGEMA_signal_3538, SubBytesInput[16]}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_4770, new_AGEMA_signal_4769, new_AGEMA_signal_4768, SubBytesIns_Inst_Sbox_2_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_4770, new_AGEMA_signal_4769, new_AGEMA_signal_4768, SubBytesIns_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, new_AGEMA_signal_4765, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_4890, new_AGEMA_signal_4889, new_AGEMA_signal_4888, SubBytesIns_Inst_Sbox_2_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_4518, new_AGEMA_signal_4517, new_AGEMA_signal_4516, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_4632, new_AGEMA_signal_4631, new_AGEMA_signal_4630, SubBytesIns_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, new_AGEMA_signal_4771, SubBytesIns_Inst_Sbox_2_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_4638, new_AGEMA_signal_4637, new_AGEMA_signal_4636, SubBytesIns_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_4623, new_AGEMA_signal_4622, new_AGEMA_signal_4621, SubBytesIns_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270], Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_4776, new_AGEMA_signal_4775, new_AGEMA_signal_4774, SubBytesIns_Inst_Sbox_2_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_9925, new_AGEMA_signal_9924, new_AGEMA_signal_9923, new_AGEMA_signal_9922}), .b ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, new_AGEMA_signal_4771, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_4893, new_AGEMA_signal_4892, new_AGEMA_signal_4891, SubBytesIns_Inst_Sbox_2_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_4758, new_AGEMA_signal_4757, new_AGEMA_signal_4756, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, new_AGEMA_signal_4753, SubBytesIns_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_4896, new_AGEMA_signal_4895, new_AGEMA_signal_4894, SubBytesIns_Inst_Sbox_2_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_4896, new_AGEMA_signal_4895, new_AGEMA_signal_4894, SubBytesIns_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, new_AGEMA_signal_4771, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_4962, new_AGEMA_signal_4961, new_AGEMA_signal_4960, SubBytesIns_Inst_Sbox_2_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_4512, new_AGEMA_signal_4511, new_AGEMA_signal_4510, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_4629, new_AGEMA_signal_4628, new_AGEMA_signal_4627, SubBytesIns_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, new_AGEMA_signal_4777, SubBytesIns_Inst_Sbox_2_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_4521, new_AGEMA_signal_4520, new_AGEMA_signal_4519, SubBytesIns_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_4641, new_AGEMA_signal_4640, new_AGEMA_signal_4639, SubBytesIns_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_4782, new_AGEMA_signal_4781, new_AGEMA_signal_4780, SubBytesIns_Inst_Sbox_2_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_4782, new_AGEMA_signal_4781, new_AGEMA_signal_4780, SubBytesIns_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, new_AGEMA_signal_4777, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_4899, new_AGEMA_signal_4898, new_AGEMA_signal_4897, SubBytesIns_Inst_Sbox_2_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_4515, new_AGEMA_signal_4514, new_AGEMA_signal_4513, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, new_AGEMA_signal_4747, SubBytesIns_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_4902, new_AGEMA_signal_4901, new_AGEMA_signal_4900, SubBytesIns_Inst_Sbox_2_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_4902, new_AGEMA_signal_4901, new_AGEMA_signal_4900, SubBytesIns_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, new_AGEMA_signal_4777, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, new_AGEMA_signal_4963, SubBytesIns_Inst_Sbox_2_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, SubBytesIns_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_4884, new_AGEMA_signal_4883, new_AGEMA_signal_4882, SubBytesIns_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, SubBytesIns_Inst_Sbox_2_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_4890, new_AGEMA_signal_4889, new_AGEMA_signal_4888, SubBytesIns_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_9929, new_AGEMA_signal_9928, new_AGEMA_signal_9927, new_AGEMA_signal_9926}), .c ({new_AGEMA_signal_4971, new_AGEMA_signal_4970, new_AGEMA_signal_4969, SubBytesIns_Inst_Sbox_2_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_4893, new_AGEMA_signal_4892, new_AGEMA_signal_4891, SubBytesIns_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_4776, new_AGEMA_signal_4775, new_AGEMA_signal_4774, SubBytesIns_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_4974, new_AGEMA_signal_4973, new_AGEMA_signal_4972, SubBytesIns_Inst_Sbox_2_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_4962, new_AGEMA_signal_4961, new_AGEMA_signal_4960, SubBytesIns_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, new_AGEMA_signal_4963, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_5016, new_AGEMA_signal_5015, new_AGEMA_signal_5014, SubBytesIns_Inst_Sbox_2_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, SubBytesIns_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_4899, new_AGEMA_signal_4898, new_AGEMA_signal_4897, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, new_AGEMA_signal_5017, SubBytesIns_Inst_Sbox_2_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_4971, new_AGEMA_signal_4970, new_AGEMA_signal_4969, SubBytesIns_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, new_AGEMA_signal_4963, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, SubBytesIns_Inst_Sbox_2_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_4974, new_AGEMA_signal_4973, new_AGEMA_signal_4972, SubBytesIns_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_4899, new_AGEMA_signal_4898, new_AGEMA_signal_4897, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_5025, new_AGEMA_signal_5024, new_AGEMA_signal_5023, SubBytesIns_Inst_Sbox_2_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_5016, new_AGEMA_signal_5015, new_AGEMA_signal_5014, SubBytesIns_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_9933, new_AGEMA_signal_9932, new_AGEMA_signal_9931, new_AGEMA_signal_9930}), .c ({new_AGEMA_signal_5064, new_AGEMA_signal_5063, new_AGEMA_signal_5062, SubBytesIns_Inst_Sbox_2_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_5025, new_AGEMA_signal_5024, new_AGEMA_signal_5023, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_5064, new_AGEMA_signal_5063, new_AGEMA_signal_5062, SubBytesIns_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_5118, new_AGEMA_signal_5117, new_AGEMA_signal_5116, SubBytesIns_Inst_Sbox_2_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, new_AGEMA_signal_5017, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, SubBytesIns_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_5070, new_AGEMA_signal_5069, new_AGEMA_signal_5068, SubBytesIns_Inst_Sbox_2_M27}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_4650, new_AGEMA_signal_4649, new_AGEMA_signal_4648, SubBytesIns_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_4644, new_AGEMA_signal_4643, new_AGEMA_signal_4642, SubBytesIns_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330], Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_4806, new_AGEMA_signal_4805, new_AGEMA_signal_4804, SubBytesIns_Inst_Sbox_3_M1}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_4800, new_AGEMA_signal_4799, new_AGEMA_signal_4798, SubBytesIns_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_4785, new_AGEMA_signal_4784, new_AGEMA_signal_4783, SubBytesIns_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, new_AGEMA_signal_4909, SubBytesIns_Inst_Sbox_3_M2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_9937, new_AGEMA_signal_9936, new_AGEMA_signal_9935, new_AGEMA_signal_9934}), .b ({new_AGEMA_signal_4806, new_AGEMA_signal_4805, new_AGEMA_signal_4804, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, new_AGEMA_signal_4912, SubBytesIns_Inst_Sbox_3_M3}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_4659, new_AGEMA_signal_4658, new_AGEMA_signal_4657, SubBytesIns_Inst_Sbox_3_T19}), .b ({new_AGEMA_signal_3564, new_AGEMA_signal_3563, new_AGEMA_signal_3562, SubBytesInput[24]}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_4809, new_AGEMA_signal_4808, new_AGEMA_signal_4807, SubBytesIns_Inst_Sbox_3_M4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_4809, new_AGEMA_signal_4808, new_AGEMA_signal_4807, SubBytesIns_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_4806, new_AGEMA_signal_4805, new_AGEMA_signal_4804, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_4917, new_AGEMA_signal_4916, new_AGEMA_signal_4915, SubBytesIns_Inst_Sbox_3_M5}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_4548, new_AGEMA_signal_4547, new_AGEMA_signal_4546, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_4656, new_AGEMA_signal_4655, new_AGEMA_signal_4654, SubBytesIns_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_4812, new_AGEMA_signal_4811, new_AGEMA_signal_4810, SubBytesIns_Inst_Sbox_3_M6}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_4662, new_AGEMA_signal_4661, new_AGEMA_signal_4660, SubBytesIns_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, new_AGEMA_signal_4645, SubBytesIns_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, new_AGEMA_signal_4813, SubBytesIns_Inst_Sbox_3_M7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_9941, new_AGEMA_signal_9940, new_AGEMA_signal_9939, new_AGEMA_signal_9938}), .b ({new_AGEMA_signal_4812, new_AGEMA_signal_4811, new_AGEMA_signal_4810, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_4920, new_AGEMA_signal_4919, new_AGEMA_signal_4918, SubBytesIns_Inst_Sbox_3_M8}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, new_AGEMA_signal_4795, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_4794, new_AGEMA_signal_4793, new_AGEMA_signal_4792, SubBytesIns_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390], Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, new_AGEMA_signal_4921, SubBytesIns_Inst_Sbox_3_M9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, new_AGEMA_signal_4921, SubBytesIns_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_4812, new_AGEMA_signal_4811, new_AGEMA_signal_4810, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_4977, new_AGEMA_signal_4976, new_AGEMA_signal_4975, SubBytesIns_Inst_Sbox_3_M10}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_4542, new_AGEMA_signal_4541, new_AGEMA_signal_4540, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, SubBytesIns_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_4818, new_AGEMA_signal_4817, new_AGEMA_signal_4816, SubBytesIns_Inst_Sbox_3_M11}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_4551, new_AGEMA_signal_4550, new_AGEMA_signal_4549, SubBytesIns_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_4665, new_AGEMA_signal_4664, new_AGEMA_signal_4663, SubBytesIns_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_4821, new_AGEMA_signal_4820, new_AGEMA_signal_4819, SubBytesIns_Inst_Sbox_3_M12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_4821, new_AGEMA_signal_4820, new_AGEMA_signal_4819, SubBytesIns_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_4818, new_AGEMA_signal_4817, new_AGEMA_signal_4816, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_4926, new_AGEMA_signal_4925, new_AGEMA_signal_4924, SubBytesIns_Inst_Sbox_3_M13}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_4545, new_AGEMA_signal_4544, new_AGEMA_signal_4543, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_4788, new_AGEMA_signal_4787, new_AGEMA_signal_4786, SubBytesIns_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, new_AGEMA_signal_4927, SubBytesIns_Inst_Sbox_3_M14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, new_AGEMA_signal_4927, SubBytesIns_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_4818, new_AGEMA_signal_4817, new_AGEMA_signal_4816, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_4980, new_AGEMA_signal_4979, new_AGEMA_signal_4978, SubBytesIns_Inst_Sbox_3_M15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, new_AGEMA_signal_4912, SubBytesIns_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, new_AGEMA_signal_4909, SubBytesIns_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_4983, new_AGEMA_signal_4982, new_AGEMA_signal_4981, SubBytesIns_Inst_Sbox_3_M16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_4917, new_AGEMA_signal_4916, new_AGEMA_signal_4915, SubBytesIns_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_9945, new_AGEMA_signal_9944, new_AGEMA_signal_9943, new_AGEMA_signal_9942}), .c ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, new_AGEMA_signal_4984, SubBytesIns_Inst_Sbox_3_M17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_4920, new_AGEMA_signal_4919, new_AGEMA_signal_4918, SubBytesIns_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, new_AGEMA_signal_4813, SubBytesIns_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_4989, new_AGEMA_signal_4988, new_AGEMA_signal_4987, SubBytesIns_Inst_Sbox_3_M18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_4977, new_AGEMA_signal_4976, new_AGEMA_signal_4975, SubBytesIns_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_4980, new_AGEMA_signal_4979, new_AGEMA_signal_4978, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_5028, new_AGEMA_signal_5027, new_AGEMA_signal_5026, SubBytesIns_Inst_Sbox_3_M19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_4983, new_AGEMA_signal_4982, new_AGEMA_signal_4981, SubBytesIns_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_4926, new_AGEMA_signal_4925, new_AGEMA_signal_4924, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, new_AGEMA_signal_5029, SubBytesIns_Inst_Sbox_3_M20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, new_AGEMA_signal_4984, SubBytesIns_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_4980, new_AGEMA_signal_4979, new_AGEMA_signal_4978, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_5034, new_AGEMA_signal_5033, new_AGEMA_signal_5032, SubBytesIns_Inst_Sbox_3_M21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_4989, new_AGEMA_signal_4988, new_AGEMA_signal_4987, SubBytesIns_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_4926, new_AGEMA_signal_4925, new_AGEMA_signal_4924, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, new_AGEMA_signal_5035, SubBytesIns_Inst_Sbox_3_M22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_5028, new_AGEMA_signal_5027, new_AGEMA_signal_5026, SubBytesIns_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_9949, new_AGEMA_signal_9948, new_AGEMA_signal_9947, new_AGEMA_signal_9946}), .c ({new_AGEMA_signal_5076, new_AGEMA_signal_5075, new_AGEMA_signal_5074, SubBytesIns_Inst_Sbox_3_M23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, new_AGEMA_signal_5035, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_5076, new_AGEMA_signal_5075, new_AGEMA_signal_5074, SubBytesIns_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_5133, new_AGEMA_signal_5132, new_AGEMA_signal_5131, SubBytesIns_Inst_Sbox_3_M24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, new_AGEMA_signal_5029, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_5034, new_AGEMA_signal_5033, new_AGEMA_signal_5032, SubBytesIns_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_5082, new_AGEMA_signal_5081, new_AGEMA_signal_5080, SubBytesIns_Inst_Sbox_3_M27}) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2061 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T14), .Q (new_AGEMA_signal_9886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2062 ( .C (clk), .D (new_AGEMA_signal_4672), .Q (new_AGEMA_signal_9887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2063 ( .C (clk), .D (new_AGEMA_signal_4673), .Q (new_AGEMA_signal_9888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2064 ( .C (clk), .D (new_AGEMA_signal_4674), .Q (new_AGEMA_signal_9889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2065 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T26), .Q (new_AGEMA_signal_9890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2066 ( .C (clk), .D (new_AGEMA_signal_4684), .Q (new_AGEMA_signal_9891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2067 ( .C (clk), .D (new_AGEMA_signal_4685), .Q (new_AGEMA_signal_9892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2068 ( .C (clk), .D (new_AGEMA_signal_4686), .Q (new_AGEMA_signal_9893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2069 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T24), .Q (new_AGEMA_signal_9894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2070 ( .C (clk), .D (new_AGEMA_signal_4822), .Q (new_AGEMA_signal_9895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2071 ( .C (clk), .D (new_AGEMA_signal_4823), .Q (new_AGEMA_signal_9896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2072 ( .C (clk), .D (new_AGEMA_signal_4824), .Q (new_AGEMA_signal_9897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2073 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T25), .Q (new_AGEMA_signal_9898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2074 ( .C (clk), .D (new_AGEMA_signal_4825), .Q (new_AGEMA_signal_9899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2075 ( .C (clk), .D (new_AGEMA_signal_4826), .Q (new_AGEMA_signal_9900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2076 ( .C (clk), .D (new_AGEMA_signal_4827), .Q (new_AGEMA_signal_9901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2077 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T14), .Q (new_AGEMA_signal_9902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2078 ( .C (clk), .D (new_AGEMA_signal_4711), .Q (new_AGEMA_signal_9903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2079 ( .C (clk), .D (new_AGEMA_signal_4712), .Q (new_AGEMA_signal_9904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2080 ( .C (clk), .D (new_AGEMA_signal_4713), .Q (new_AGEMA_signal_9905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2081 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T26), .Q (new_AGEMA_signal_9906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2082 ( .C (clk), .D (new_AGEMA_signal_4723), .Q (new_AGEMA_signal_9907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2083 ( .C (clk), .D (new_AGEMA_signal_4724), .Q (new_AGEMA_signal_9908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2084 ( .C (clk), .D (new_AGEMA_signal_4725), .Q (new_AGEMA_signal_9909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2085 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T24), .Q (new_AGEMA_signal_9910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2086 ( .C (clk), .D (new_AGEMA_signal_4849), .Q (new_AGEMA_signal_9911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2087 ( .C (clk), .D (new_AGEMA_signal_4850), .Q (new_AGEMA_signal_9912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2088 ( .C (clk), .D (new_AGEMA_signal_4851), .Q (new_AGEMA_signal_9913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2089 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T25), .Q (new_AGEMA_signal_9914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2090 ( .C (clk), .D (new_AGEMA_signal_4852), .Q (new_AGEMA_signal_9915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2091 ( .C (clk), .D (new_AGEMA_signal_4853), .Q (new_AGEMA_signal_9916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2092 ( .C (clk), .D (new_AGEMA_signal_4854), .Q (new_AGEMA_signal_9917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2093 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T14), .Q (new_AGEMA_signal_9918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2094 ( .C (clk), .D (new_AGEMA_signal_4750), .Q (new_AGEMA_signal_9919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2095 ( .C (clk), .D (new_AGEMA_signal_4751), .Q (new_AGEMA_signal_9920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2096 ( .C (clk), .D (new_AGEMA_signal_4752), .Q (new_AGEMA_signal_9921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2097 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T26), .Q (new_AGEMA_signal_9922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2098 ( .C (clk), .D (new_AGEMA_signal_4762), .Q (new_AGEMA_signal_9923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2099 ( .C (clk), .D (new_AGEMA_signal_4763), .Q (new_AGEMA_signal_9924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2100 ( .C (clk), .D (new_AGEMA_signal_4764), .Q (new_AGEMA_signal_9925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2101 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T24), .Q (new_AGEMA_signal_9926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2102 ( .C (clk), .D (new_AGEMA_signal_4876), .Q (new_AGEMA_signal_9927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2103 ( .C (clk), .D (new_AGEMA_signal_4877), .Q (new_AGEMA_signal_9928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2104 ( .C (clk), .D (new_AGEMA_signal_4878), .Q (new_AGEMA_signal_9929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2105 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T25), .Q (new_AGEMA_signal_9930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2106 ( .C (clk), .D (new_AGEMA_signal_4879), .Q (new_AGEMA_signal_9931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2107 ( .C (clk), .D (new_AGEMA_signal_4880), .Q (new_AGEMA_signal_9932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2108 ( .C (clk), .D (new_AGEMA_signal_4881), .Q (new_AGEMA_signal_9933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2109 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T14), .Q (new_AGEMA_signal_9934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2110 ( .C (clk), .D (new_AGEMA_signal_4789), .Q (new_AGEMA_signal_9935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2111 ( .C (clk), .D (new_AGEMA_signal_4790), .Q (new_AGEMA_signal_9936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2112 ( .C (clk), .D (new_AGEMA_signal_4791), .Q (new_AGEMA_signal_9937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2113 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T26), .Q (new_AGEMA_signal_9938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2114 ( .C (clk), .D (new_AGEMA_signal_4801), .Q (new_AGEMA_signal_9939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2115 ( .C (clk), .D (new_AGEMA_signal_4802), .Q (new_AGEMA_signal_9940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2116 ( .C (clk), .D (new_AGEMA_signal_4803), .Q (new_AGEMA_signal_9941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2117 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T24), .Q (new_AGEMA_signal_9942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2118 ( .C (clk), .D (new_AGEMA_signal_4903), .Q (new_AGEMA_signal_9943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2119 ( .C (clk), .D (new_AGEMA_signal_4904), .Q (new_AGEMA_signal_9944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2120 ( .C (clk), .D (new_AGEMA_signal_4905), .Q (new_AGEMA_signal_9945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2121 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T25), .Q (new_AGEMA_signal_9946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2122 ( .C (clk), .D (new_AGEMA_signal_4906), .Q (new_AGEMA_signal_9947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2123 ( .C (clk), .D (new_AGEMA_signal_4907), .Q (new_AGEMA_signal_9948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2124 ( .C (clk), .D (new_AGEMA_signal_4908), .Q (new_AGEMA_signal_9949) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C (clk), .D (reset), .Q (new_AGEMA_signal_10078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2257 ( .C (clk), .D (plaintext_s0[0]), .Q (new_AGEMA_signal_10082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2261 ( .C (clk), .D (plaintext_s1[0]), .Q (new_AGEMA_signal_10086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2265 ( .C (clk), .D (plaintext_s2[0]), .Q (new_AGEMA_signal_10090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2269 ( .C (clk), .D (plaintext_s3[0]), .Q (new_AGEMA_signal_10094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2273 ( .C (clk), .D (plaintext_s0[1]), .Q (new_AGEMA_signal_10098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2277 ( .C (clk), .D (plaintext_s1[1]), .Q (new_AGEMA_signal_10102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2281 ( .C (clk), .D (plaintext_s2[1]), .Q (new_AGEMA_signal_10106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2285 ( .C (clk), .D (plaintext_s3[1]), .Q (new_AGEMA_signal_10110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2289 ( .C (clk), .D (plaintext_s0[2]), .Q (new_AGEMA_signal_10114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2293 ( .C (clk), .D (plaintext_s1[2]), .Q (new_AGEMA_signal_10118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2297 ( .C (clk), .D (plaintext_s2[2]), .Q (new_AGEMA_signal_10122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2301 ( .C (clk), .D (plaintext_s3[2]), .Q (new_AGEMA_signal_10126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2305 ( .C (clk), .D (plaintext_s0[3]), .Q (new_AGEMA_signal_10130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2309 ( .C (clk), .D (plaintext_s1[3]), .Q (new_AGEMA_signal_10134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2313 ( .C (clk), .D (plaintext_s2[3]), .Q (new_AGEMA_signal_10138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2317 ( .C (clk), .D (plaintext_s3[3]), .Q (new_AGEMA_signal_10142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2321 ( .C (clk), .D (plaintext_s0[4]), .Q (new_AGEMA_signal_10146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2325 ( .C (clk), .D (plaintext_s1[4]), .Q (new_AGEMA_signal_10150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2329 ( .C (clk), .D (plaintext_s2[4]), .Q (new_AGEMA_signal_10154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2333 ( .C (clk), .D (plaintext_s3[4]), .Q (new_AGEMA_signal_10158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2337 ( .C (clk), .D (plaintext_s0[5]), .Q (new_AGEMA_signal_10162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2341 ( .C (clk), .D (plaintext_s1[5]), .Q (new_AGEMA_signal_10166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2345 ( .C (clk), .D (plaintext_s2[5]), .Q (new_AGEMA_signal_10170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2349 ( .C (clk), .D (plaintext_s3[5]), .Q (new_AGEMA_signal_10174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2353 ( .C (clk), .D (plaintext_s0[6]), .Q (new_AGEMA_signal_10178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2357 ( .C (clk), .D (plaintext_s1[6]), .Q (new_AGEMA_signal_10182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2361 ( .C (clk), .D (plaintext_s2[6]), .Q (new_AGEMA_signal_10186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2365 ( .C (clk), .D (plaintext_s3[6]), .Q (new_AGEMA_signal_10190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2369 ( .C (clk), .D (plaintext_s0[7]), .Q (new_AGEMA_signal_10194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2373 ( .C (clk), .D (plaintext_s1[7]), .Q (new_AGEMA_signal_10198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2377 ( .C (clk), .D (plaintext_s2[7]), .Q (new_AGEMA_signal_10202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2381 ( .C (clk), .D (plaintext_s3[7]), .Q (new_AGEMA_signal_10206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2385 ( .C (clk), .D (plaintext_s0[8]), .Q (new_AGEMA_signal_10210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2389 ( .C (clk), .D (plaintext_s1[8]), .Q (new_AGEMA_signal_10214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2393 ( .C (clk), .D (plaintext_s2[8]), .Q (new_AGEMA_signal_10218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2397 ( .C (clk), .D (plaintext_s3[8]), .Q (new_AGEMA_signal_10222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2401 ( .C (clk), .D (plaintext_s0[9]), .Q (new_AGEMA_signal_10226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2405 ( .C (clk), .D (plaintext_s1[9]), .Q (new_AGEMA_signal_10230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2409 ( .C (clk), .D (plaintext_s2[9]), .Q (new_AGEMA_signal_10234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2413 ( .C (clk), .D (plaintext_s3[9]), .Q (new_AGEMA_signal_10238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2417 ( .C (clk), .D (plaintext_s0[10]), .Q (new_AGEMA_signal_10242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2421 ( .C (clk), .D (plaintext_s1[10]), .Q (new_AGEMA_signal_10246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2425 ( .C (clk), .D (plaintext_s2[10]), .Q (new_AGEMA_signal_10250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2429 ( .C (clk), .D (plaintext_s3[10]), .Q (new_AGEMA_signal_10254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2433 ( .C (clk), .D (plaintext_s0[11]), .Q (new_AGEMA_signal_10258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2437 ( .C (clk), .D (plaintext_s1[11]), .Q (new_AGEMA_signal_10262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2441 ( .C (clk), .D (plaintext_s2[11]), .Q (new_AGEMA_signal_10266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2445 ( .C (clk), .D (plaintext_s3[11]), .Q (new_AGEMA_signal_10270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2449 ( .C (clk), .D (plaintext_s0[12]), .Q (new_AGEMA_signal_10274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2453 ( .C (clk), .D (plaintext_s1[12]), .Q (new_AGEMA_signal_10278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2457 ( .C (clk), .D (plaintext_s2[12]), .Q (new_AGEMA_signal_10282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2461 ( .C (clk), .D (plaintext_s3[12]), .Q (new_AGEMA_signal_10286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2465 ( .C (clk), .D (plaintext_s0[13]), .Q (new_AGEMA_signal_10290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2469 ( .C (clk), .D (plaintext_s1[13]), .Q (new_AGEMA_signal_10294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2473 ( .C (clk), .D (plaintext_s2[13]), .Q (new_AGEMA_signal_10298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2477 ( .C (clk), .D (plaintext_s3[13]), .Q (new_AGEMA_signal_10302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2481 ( .C (clk), .D (plaintext_s0[14]), .Q (new_AGEMA_signal_10306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2485 ( .C (clk), .D (plaintext_s1[14]), .Q (new_AGEMA_signal_10310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2489 ( .C (clk), .D (plaintext_s2[14]), .Q (new_AGEMA_signal_10314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2493 ( .C (clk), .D (plaintext_s3[14]), .Q (new_AGEMA_signal_10318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2497 ( .C (clk), .D (plaintext_s0[15]), .Q (new_AGEMA_signal_10322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2501 ( .C (clk), .D (plaintext_s1[15]), .Q (new_AGEMA_signal_10326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2505 ( .C (clk), .D (plaintext_s2[15]), .Q (new_AGEMA_signal_10330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2509 ( .C (clk), .D (plaintext_s3[15]), .Q (new_AGEMA_signal_10334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2513 ( .C (clk), .D (plaintext_s0[16]), .Q (new_AGEMA_signal_10338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2517 ( .C (clk), .D (plaintext_s1[16]), .Q (new_AGEMA_signal_10342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2521 ( .C (clk), .D (plaintext_s2[16]), .Q (new_AGEMA_signal_10346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2525 ( .C (clk), .D (plaintext_s3[16]), .Q (new_AGEMA_signal_10350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2529 ( .C (clk), .D (plaintext_s0[17]), .Q (new_AGEMA_signal_10354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2533 ( .C (clk), .D (plaintext_s1[17]), .Q (new_AGEMA_signal_10358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2537 ( .C (clk), .D (plaintext_s2[17]), .Q (new_AGEMA_signal_10362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2541 ( .C (clk), .D (plaintext_s3[17]), .Q (new_AGEMA_signal_10366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2545 ( .C (clk), .D (plaintext_s0[18]), .Q (new_AGEMA_signal_10370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2549 ( .C (clk), .D (plaintext_s1[18]), .Q (new_AGEMA_signal_10374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2553 ( .C (clk), .D (plaintext_s2[18]), .Q (new_AGEMA_signal_10378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2557 ( .C (clk), .D (plaintext_s3[18]), .Q (new_AGEMA_signal_10382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2561 ( .C (clk), .D (plaintext_s0[19]), .Q (new_AGEMA_signal_10386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2565 ( .C (clk), .D (plaintext_s1[19]), .Q (new_AGEMA_signal_10390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2569 ( .C (clk), .D (plaintext_s2[19]), .Q (new_AGEMA_signal_10394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2573 ( .C (clk), .D (plaintext_s3[19]), .Q (new_AGEMA_signal_10398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2577 ( .C (clk), .D (plaintext_s0[20]), .Q (new_AGEMA_signal_10402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2581 ( .C (clk), .D (plaintext_s1[20]), .Q (new_AGEMA_signal_10406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2585 ( .C (clk), .D (plaintext_s2[20]), .Q (new_AGEMA_signal_10410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2589 ( .C (clk), .D (plaintext_s3[20]), .Q (new_AGEMA_signal_10414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2593 ( .C (clk), .D (plaintext_s0[21]), .Q (new_AGEMA_signal_10418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2597 ( .C (clk), .D (plaintext_s1[21]), .Q (new_AGEMA_signal_10422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2601 ( .C (clk), .D (plaintext_s2[21]), .Q (new_AGEMA_signal_10426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2605 ( .C (clk), .D (plaintext_s3[21]), .Q (new_AGEMA_signal_10430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2609 ( .C (clk), .D (plaintext_s0[22]), .Q (new_AGEMA_signal_10434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2613 ( .C (clk), .D (plaintext_s1[22]), .Q (new_AGEMA_signal_10438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2617 ( .C (clk), .D (plaintext_s2[22]), .Q (new_AGEMA_signal_10442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2621 ( .C (clk), .D (plaintext_s3[22]), .Q (new_AGEMA_signal_10446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2625 ( .C (clk), .D (plaintext_s0[23]), .Q (new_AGEMA_signal_10450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2629 ( .C (clk), .D (plaintext_s1[23]), .Q (new_AGEMA_signal_10454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2633 ( .C (clk), .D (plaintext_s2[23]), .Q (new_AGEMA_signal_10458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2637 ( .C (clk), .D (plaintext_s3[23]), .Q (new_AGEMA_signal_10462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2641 ( .C (clk), .D (plaintext_s0[24]), .Q (new_AGEMA_signal_10466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2645 ( .C (clk), .D (plaintext_s1[24]), .Q (new_AGEMA_signal_10470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2649 ( .C (clk), .D (plaintext_s2[24]), .Q (new_AGEMA_signal_10474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2653 ( .C (clk), .D (plaintext_s3[24]), .Q (new_AGEMA_signal_10478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2657 ( .C (clk), .D (plaintext_s0[25]), .Q (new_AGEMA_signal_10482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2661 ( .C (clk), .D (plaintext_s1[25]), .Q (new_AGEMA_signal_10486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2665 ( .C (clk), .D (plaintext_s2[25]), .Q (new_AGEMA_signal_10490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2669 ( .C (clk), .D (plaintext_s3[25]), .Q (new_AGEMA_signal_10494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2673 ( .C (clk), .D (plaintext_s0[26]), .Q (new_AGEMA_signal_10498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2677 ( .C (clk), .D (plaintext_s1[26]), .Q (new_AGEMA_signal_10502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2681 ( .C (clk), .D (plaintext_s2[26]), .Q (new_AGEMA_signal_10506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2685 ( .C (clk), .D (plaintext_s3[26]), .Q (new_AGEMA_signal_10510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2689 ( .C (clk), .D (plaintext_s0[27]), .Q (new_AGEMA_signal_10514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2693 ( .C (clk), .D (plaintext_s1[27]), .Q (new_AGEMA_signal_10518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2697 ( .C (clk), .D (plaintext_s2[27]), .Q (new_AGEMA_signal_10522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2701 ( .C (clk), .D (plaintext_s3[27]), .Q (new_AGEMA_signal_10526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2705 ( .C (clk), .D (plaintext_s0[28]), .Q (new_AGEMA_signal_10530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2709 ( .C (clk), .D (plaintext_s1[28]), .Q (new_AGEMA_signal_10534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2713 ( .C (clk), .D (plaintext_s2[28]), .Q (new_AGEMA_signal_10538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2717 ( .C (clk), .D (plaintext_s3[28]), .Q (new_AGEMA_signal_10542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2721 ( .C (clk), .D (plaintext_s0[29]), .Q (new_AGEMA_signal_10546) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2725 ( .C (clk), .D (plaintext_s1[29]), .Q (new_AGEMA_signal_10550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2729 ( .C (clk), .D (plaintext_s2[29]), .Q (new_AGEMA_signal_10554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2733 ( .C (clk), .D (plaintext_s3[29]), .Q (new_AGEMA_signal_10558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2737 ( .C (clk), .D (plaintext_s0[30]), .Q (new_AGEMA_signal_10562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2741 ( .C (clk), .D (plaintext_s1[30]), .Q (new_AGEMA_signal_10566) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2745 ( .C (clk), .D (plaintext_s2[30]), .Q (new_AGEMA_signal_10570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2749 ( .C (clk), .D (plaintext_s3[30]), .Q (new_AGEMA_signal_10574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2753 ( .C (clk), .D (plaintext_s0[31]), .Q (new_AGEMA_signal_10578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2757 ( .C (clk), .D (plaintext_s1[31]), .Q (new_AGEMA_signal_10582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2761 ( .C (clk), .D (plaintext_s2[31]), .Q (new_AGEMA_signal_10586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2765 ( .C (clk), .D (plaintext_s3[31]), .Q (new_AGEMA_signal_10590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2769 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T6), .Q (new_AGEMA_signal_10594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2772 ( .C (clk), .D (new_AGEMA_signal_4570), .Q (new_AGEMA_signal_10597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2775 ( .C (clk), .D (new_AGEMA_signal_4571), .Q (new_AGEMA_signal_10600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2778 ( .C (clk), .D (new_AGEMA_signal_4572), .Q (new_AGEMA_signal_10603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2781 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T8), .Q (new_AGEMA_signal_10606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2784 ( .C (clk), .D (new_AGEMA_signal_4666), .Q (new_AGEMA_signal_10609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2787 ( .C (clk), .D (new_AGEMA_signal_4667), .Q (new_AGEMA_signal_10612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2790 ( .C (clk), .D (new_AGEMA_signal_4668), .Q (new_AGEMA_signal_10615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2793 ( .C (clk), .D (SubBytesInput[0]), .Q (new_AGEMA_signal_10618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2796 ( .C (clk), .D (new_AGEMA_signal_3493), .Q (new_AGEMA_signal_10621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2799 ( .C (clk), .D (new_AGEMA_signal_3494), .Q (new_AGEMA_signal_10624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2802 ( .C (clk), .D (new_AGEMA_signal_3495), .Q (new_AGEMA_signal_10627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2805 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T16), .Q (new_AGEMA_signal_10630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2808 ( .C (clk), .D (new_AGEMA_signal_4582), .Q (new_AGEMA_signal_10633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2811 ( .C (clk), .D (new_AGEMA_signal_4583), .Q (new_AGEMA_signal_10636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2814 ( .C (clk), .D (new_AGEMA_signal_4584), .Q (new_AGEMA_signal_10639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2817 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T9), .Q (new_AGEMA_signal_10642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2820 ( .C (clk), .D (new_AGEMA_signal_4573), .Q (new_AGEMA_signal_10645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2823 ( .C (clk), .D (new_AGEMA_signal_4574), .Q (new_AGEMA_signal_10648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2826 ( .C (clk), .D (new_AGEMA_signal_4575), .Q (new_AGEMA_signal_10651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2829 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T17), .Q (new_AGEMA_signal_10654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2832 ( .C (clk), .D (new_AGEMA_signal_4675), .Q (new_AGEMA_signal_10657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2835 ( .C (clk), .D (new_AGEMA_signal_4676), .Q (new_AGEMA_signal_10660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2838 ( .C (clk), .D (new_AGEMA_signal_4677), .Q (new_AGEMA_signal_10663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2841 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T15), .Q (new_AGEMA_signal_10666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2844 ( .C (clk), .D (new_AGEMA_signal_4579), .Q (new_AGEMA_signal_10669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2847 ( .C (clk), .D (new_AGEMA_signal_4580), .Q (new_AGEMA_signal_10672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2850 ( .C (clk), .D (new_AGEMA_signal_4581), .Q (new_AGEMA_signal_10675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2853 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T27), .Q (new_AGEMA_signal_10678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2856 ( .C (clk), .D (new_AGEMA_signal_4591), .Q (new_AGEMA_signal_10681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2859 ( .C (clk), .D (new_AGEMA_signal_4592), .Q (new_AGEMA_signal_10684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2862 ( .C (clk), .D (new_AGEMA_signal_4593), .Q (new_AGEMA_signal_10687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2865 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T10), .Q (new_AGEMA_signal_10690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2868 ( .C (clk), .D (new_AGEMA_signal_4669), .Q (new_AGEMA_signal_10693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2871 ( .C (clk), .D (new_AGEMA_signal_4670), .Q (new_AGEMA_signal_10696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2874 ( .C (clk), .D (new_AGEMA_signal_4671), .Q (new_AGEMA_signal_10699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2877 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T13), .Q (new_AGEMA_signal_10702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2880 ( .C (clk), .D (new_AGEMA_signal_4576), .Q (new_AGEMA_signal_10705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2883 ( .C (clk), .D (new_AGEMA_signal_4577), .Q (new_AGEMA_signal_10708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2886 ( .C (clk), .D (new_AGEMA_signal_4578), .Q (new_AGEMA_signal_10711) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2889 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T23), .Q (new_AGEMA_signal_10714) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2892 ( .C (clk), .D (new_AGEMA_signal_4681), .Q (new_AGEMA_signal_10717) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2895 ( .C (clk), .D (new_AGEMA_signal_4682), .Q (new_AGEMA_signal_10720) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2898 ( .C (clk), .D (new_AGEMA_signal_4683), .Q (new_AGEMA_signal_10723) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2901 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T19), .Q (new_AGEMA_signal_10726) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2904 ( .C (clk), .D (new_AGEMA_signal_4585), .Q (new_AGEMA_signal_10729) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2907 ( .C (clk), .D (new_AGEMA_signal_4586), .Q (new_AGEMA_signal_10732) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2910 ( .C (clk), .D (new_AGEMA_signal_4587), .Q (new_AGEMA_signal_10735) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2913 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T3), .Q (new_AGEMA_signal_10738) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2916 ( .C (clk), .D (new_AGEMA_signal_4456), .Q (new_AGEMA_signal_10741) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2919 ( .C (clk), .D (new_AGEMA_signal_4457), .Q (new_AGEMA_signal_10744) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2922 ( .C (clk), .D (new_AGEMA_signal_4458), .Q (new_AGEMA_signal_10747) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2925 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T22), .Q (new_AGEMA_signal_10750) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2928 ( .C (clk), .D (new_AGEMA_signal_4588), .Q (new_AGEMA_signal_10753) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2931 ( .C (clk), .D (new_AGEMA_signal_4589), .Q (new_AGEMA_signal_10756) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2934 ( .C (clk), .D (new_AGEMA_signal_4590), .Q (new_AGEMA_signal_10759) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2937 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T20), .Q (new_AGEMA_signal_10762) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2940 ( .C (clk), .D (new_AGEMA_signal_4678), .Q (new_AGEMA_signal_10765) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2943 ( .C (clk), .D (new_AGEMA_signal_4679), .Q (new_AGEMA_signal_10768) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2946 ( .C (clk), .D (new_AGEMA_signal_4680), .Q (new_AGEMA_signal_10771) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2949 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T1), .Q (new_AGEMA_signal_10774) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2952 ( .C (clk), .D (new_AGEMA_signal_4450), .Q (new_AGEMA_signal_10777) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2955 ( .C (clk), .D (new_AGEMA_signal_4451), .Q (new_AGEMA_signal_10780) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2958 ( .C (clk), .D (new_AGEMA_signal_4452), .Q (new_AGEMA_signal_10783) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2961 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T4), .Q (new_AGEMA_signal_10786) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2964 ( .C (clk), .D (new_AGEMA_signal_4459), .Q (new_AGEMA_signal_10789) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2967 ( .C (clk), .D (new_AGEMA_signal_4460), .Q (new_AGEMA_signal_10792) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2970 ( .C (clk), .D (new_AGEMA_signal_4461), .Q (new_AGEMA_signal_10795) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2973 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T2), .Q (new_AGEMA_signal_10798) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2976 ( .C (clk), .D (new_AGEMA_signal_4453), .Q (new_AGEMA_signal_10801) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2979 ( .C (clk), .D (new_AGEMA_signal_4454), .Q (new_AGEMA_signal_10804) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2982 ( .C (clk), .D (new_AGEMA_signal_4455), .Q (new_AGEMA_signal_10807) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2985 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T6), .Q (new_AGEMA_signal_10810) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2988 ( .C (clk), .D (new_AGEMA_signal_4594), .Q (new_AGEMA_signal_10813) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2991 ( .C (clk), .D (new_AGEMA_signal_4595), .Q (new_AGEMA_signal_10816) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2994 ( .C (clk), .D (new_AGEMA_signal_4596), .Q (new_AGEMA_signal_10819) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2997 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T8), .Q (new_AGEMA_signal_10822) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3000 ( .C (clk), .D (new_AGEMA_signal_4705), .Q (new_AGEMA_signal_10825) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3003 ( .C (clk), .D (new_AGEMA_signal_4706), .Q (new_AGEMA_signal_10828) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3006 ( .C (clk), .D (new_AGEMA_signal_4707), .Q (new_AGEMA_signal_10831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3009 ( .C (clk), .D (SubBytesInput[8]), .Q (new_AGEMA_signal_10834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3012 ( .C (clk), .D (new_AGEMA_signal_3490), .Q (new_AGEMA_signal_10837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3015 ( .C (clk), .D (new_AGEMA_signal_3491), .Q (new_AGEMA_signal_10840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3018 ( .C (clk), .D (new_AGEMA_signal_3492), .Q (new_AGEMA_signal_10843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3021 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T16), .Q (new_AGEMA_signal_10846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3024 ( .C (clk), .D (new_AGEMA_signal_4606), .Q (new_AGEMA_signal_10849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3027 ( .C (clk), .D (new_AGEMA_signal_4607), .Q (new_AGEMA_signal_10852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3030 ( .C (clk), .D (new_AGEMA_signal_4608), .Q (new_AGEMA_signal_10855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3033 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T9), .Q (new_AGEMA_signal_10858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3036 ( .C (clk), .D (new_AGEMA_signal_4597), .Q (new_AGEMA_signal_10861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3039 ( .C (clk), .D (new_AGEMA_signal_4598), .Q (new_AGEMA_signal_10864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3042 ( .C (clk), .D (new_AGEMA_signal_4599), .Q (new_AGEMA_signal_10867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3045 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T17), .Q (new_AGEMA_signal_10870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3048 ( .C (clk), .D (new_AGEMA_signal_4714), .Q (new_AGEMA_signal_10873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3051 ( .C (clk), .D (new_AGEMA_signal_4715), .Q (new_AGEMA_signal_10876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3054 ( .C (clk), .D (new_AGEMA_signal_4716), .Q (new_AGEMA_signal_10879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3057 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T15), .Q (new_AGEMA_signal_10882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3060 ( .C (clk), .D (new_AGEMA_signal_4603), .Q (new_AGEMA_signal_10885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3063 ( .C (clk), .D (new_AGEMA_signal_4604), .Q (new_AGEMA_signal_10888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3066 ( .C (clk), .D (new_AGEMA_signal_4605), .Q (new_AGEMA_signal_10891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3069 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T27), .Q (new_AGEMA_signal_10894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3072 ( .C (clk), .D (new_AGEMA_signal_4615), .Q (new_AGEMA_signal_10897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3075 ( .C (clk), .D (new_AGEMA_signal_4616), .Q (new_AGEMA_signal_10900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3078 ( .C (clk), .D (new_AGEMA_signal_4617), .Q (new_AGEMA_signal_10903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3081 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T10), .Q (new_AGEMA_signal_10906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3084 ( .C (clk), .D (new_AGEMA_signal_4708), .Q (new_AGEMA_signal_10909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3087 ( .C (clk), .D (new_AGEMA_signal_4709), .Q (new_AGEMA_signal_10912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3090 ( .C (clk), .D (new_AGEMA_signal_4710), .Q (new_AGEMA_signal_10915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3093 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T13), .Q (new_AGEMA_signal_10918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3096 ( .C (clk), .D (new_AGEMA_signal_4600), .Q (new_AGEMA_signal_10921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3099 ( .C (clk), .D (new_AGEMA_signal_4601), .Q (new_AGEMA_signal_10924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3102 ( .C (clk), .D (new_AGEMA_signal_4602), .Q (new_AGEMA_signal_10927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3105 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T23), .Q (new_AGEMA_signal_10930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3108 ( .C (clk), .D (new_AGEMA_signal_4720), .Q (new_AGEMA_signal_10933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3111 ( .C (clk), .D (new_AGEMA_signal_4721), .Q (new_AGEMA_signal_10936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3114 ( .C (clk), .D (new_AGEMA_signal_4722), .Q (new_AGEMA_signal_10939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3117 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T19), .Q (new_AGEMA_signal_10942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3120 ( .C (clk), .D (new_AGEMA_signal_4609), .Q (new_AGEMA_signal_10945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3123 ( .C (clk), .D (new_AGEMA_signal_4610), .Q (new_AGEMA_signal_10948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3126 ( .C (clk), .D (new_AGEMA_signal_4611), .Q (new_AGEMA_signal_10951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3129 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T3), .Q (new_AGEMA_signal_10954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3132 ( .C (clk), .D (new_AGEMA_signal_4486), .Q (new_AGEMA_signal_10957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3135 ( .C (clk), .D (new_AGEMA_signal_4487), .Q (new_AGEMA_signal_10960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3138 ( .C (clk), .D (new_AGEMA_signal_4488), .Q (new_AGEMA_signal_10963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3141 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T22), .Q (new_AGEMA_signal_10966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3144 ( .C (clk), .D (new_AGEMA_signal_4612), .Q (new_AGEMA_signal_10969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3147 ( .C (clk), .D (new_AGEMA_signal_4613), .Q (new_AGEMA_signal_10972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3150 ( .C (clk), .D (new_AGEMA_signal_4614), .Q (new_AGEMA_signal_10975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3153 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T20), .Q (new_AGEMA_signal_10978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3156 ( .C (clk), .D (new_AGEMA_signal_4717), .Q (new_AGEMA_signal_10981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3159 ( .C (clk), .D (new_AGEMA_signal_4718), .Q (new_AGEMA_signal_10984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3162 ( .C (clk), .D (new_AGEMA_signal_4719), .Q (new_AGEMA_signal_10987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3165 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T1), .Q (new_AGEMA_signal_10990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3168 ( .C (clk), .D (new_AGEMA_signal_4480), .Q (new_AGEMA_signal_10993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3171 ( .C (clk), .D (new_AGEMA_signal_4481), .Q (new_AGEMA_signal_10996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3174 ( .C (clk), .D (new_AGEMA_signal_4482), .Q (new_AGEMA_signal_10999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3177 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T4), .Q (new_AGEMA_signal_11002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3180 ( .C (clk), .D (new_AGEMA_signal_4489), .Q (new_AGEMA_signal_11005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3183 ( .C (clk), .D (new_AGEMA_signal_4490), .Q (new_AGEMA_signal_11008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3186 ( .C (clk), .D (new_AGEMA_signal_4491), .Q (new_AGEMA_signal_11011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3189 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T2), .Q (new_AGEMA_signal_11014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3192 ( .C (clk), .D (new_AGEMA_signal_4483), .Q (new_AGEMA_signal_11017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3195 ( .C (clk), .D (new_AGEMA_signal_4484), .Q (new_AGEMA_signal_11020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3198 ( .C (clk), .D (new_AGEMA_signal_4485), .Q (new_AGEMA_signal_11023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3201 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T6), .Q (new_AGEMA_signal_11026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3204 ( .C (clk), .D (new_AGEMA_signal_4618), .Q (new_AGEMA_signal_11029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3207 ( .C (clk), .D (new_AGEMA_signal_4619), .Q (new_AGEMA_signal_11032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3210 ( .C (clk), .D (new_AGEMA_signal_4620), .Q (new_AGEMA_signal_11035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3213 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T8), .Q (new_AGEMA_signal_11038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3216 ( .C (clk), .D (new_AGEMA_signal_4744), .Q (new_AGEMA_signal_11041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3219 ( .C (clk), .D (new_AGEMA_signal_4745), .Q (new_AGEMA_signal_11044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3222 ( .C (clk), .D (new_AGEMA_signal_4746), .Q (new_AGEMA_signal_11047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3225 ( .C (clk), .D (SubBytesInput[16]), .Q (new_AGEMA_signal_11050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3228 ( .C (clk), .D (new_AGEMA_signal_3538), .Q (new_AGEMA_signal_11053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3231 ( .C (clk), .D (new_AGEMA_signal_3539), .Q (new_AGEMA_signal_11056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3234 ( .C (clk), .D (new_AGEMA_signal_3540), .Q (new_AGEMA_signal_11059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3237 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T16), .Q (new_AGEMA_signal_11062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3240 ( .C (clk), .D (new_AGEMA_signal_4630), .Q (new_AGEMA_signal_11065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3243 ( .C (clk), .D (new_AGEMA_signal_4631), .Q (new_AGEMA_signal_11068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3246 ( .C (clk), .D (new_AGEMA_signal_4632), .Q (new_AGEMA_signal_11071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3249 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T9), .Q (new_AGEMA_signal_11074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3252 ( .C (clk), .D (new_AGEMA_signal_4621), .Q (new_AGEMA_signal_11077) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3255 ( .C (clk), .D (new_AGEMA_signal_4622), .Q (new_AGEMA_signal_11080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3258 ( .C (clk), .D (new_AGEMA_signal_4623), .Q (new_AGEMA_signal_11083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3261 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T17), .Q (new_AGEMA_signal_11086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3264 ( .C (clk), .D (new_AGEMA_signal_4753), .Q (new_AGEMA_signal_11089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3267 ( .C (clk), .D (new_AGEMA_signal_4754), .Q (new_AGEMA_signal_11092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3270 ( .C (clk), .D (new_AGEMA_signal_4755), .Q (new_AGEMA_signal_11095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3273 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T15), .Q (new_AGEMA_signal_11098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3276 ( .C (clk), .D (new_AGEMA_signal_4627), .Q (new_AGEMA_signal_11101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3279 ( .C (clk), .D (new_AGEMA_signal_4628), .Q (new_AGEMA_signal_11104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3282 ( .C (clk), .D (new_AGEMA_signal_4629), .Q (new_AGEMA_signal_11107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3285 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T27), .Q (new_AGEMA_signal_11110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3288 ( .C (clk), .D (new_AGEMA_signal_4639), .Q (new_AGEMA_signal_11113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3291 ( .C (clk), .D (new_AGEMA_signal_4640), .Q (new_AGEMA_signal_11116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3294 ( .C (clk), .D (new_AGEMA_signal_4641), .Q (new_AGEMA_signal_11119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3297 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T10), .Q (new_AGEMA_signal_11122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3300 ( .C (clk), .D (new_AGEMA_signal_4747), .Q (new_AGEMA_signal_11125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3303 ( .C (clk), .D (new_AGEMA_signal_4748), .Q (new_AGEMA_signal_11128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3306 ( .C (clk), .D (new_AGEMA_signal_4749), .Q (new_AGEMA_signal_11131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3309 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T13), .Q (new_AGEMA_signal_11134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3312 ( .C (clk), .D (new_AGEMA_signal_4624), .Q (new_AGEMA_signal_11137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3315 ( .C (clk), .D (new_AGEMA_signal_4625), .Q (new_AGEMA_signal_11140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3318 ( .C (clk), .D (new_AGEMA_signal_4626), .Q (new_AGEMA_signal_11143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3321 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T23), .Q (new_AGEMA_signal_11146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3324 ( .C (clk), .D (new_AGEMA_signal_4759), .Q (new_AGEMA_signal_11149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3327 ( .C (clk), .D (new_AGEMA_signal_4760), .Q (new_AGEMA_signal_11152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3330 ( .C (clk), .D (new_AGEMA_signal_4761), .Q (new_AGEMA_signal_11155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3333 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T19), .Q (new_AGEMA_signal_11158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3336 ( .C (clk), .D (new_AGEMA_signal_4633), .Q (new_AGEMA_signal_11161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3339 ( .C (clk), .D (new_AGEMA_signal_4634), .Q (new_AGEMA_signal_11164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3342 ( .C (clk), .D (new_AGEMA_signal_4635), .Q (new_AGEMA_signal_11167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3345 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T3), .Q (new_AGEMA_signal_11170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3348 ( .C (clk), .D (new_AGEMA_signal_4516), .Q (new_AGEMA_signal_11173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3351 ( .C (clk), .D (new_AGEMA_signal_4517), .Q (new_AGEMA_signal_11176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3354 ( .C (clk), .D (new_AGEMA_signal_4518), .Q (new_AGEMA_signal_11179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3357 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T22), .Q (new_AGEMA_signal_11182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3360 ( .C (clk), .D (new_AGEMA_signal_4636), .Q (new_AGEMA_signal_11185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3363 ( .C (clk), .D (new_AGEMA_signal_4637), .Q (new_AGEMA_signal_11188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3366 ( .C (clk), .D (new_AGEMA_signal_4638), .Q (new_AGEMA_signal_11191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3369 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T20), .Q (new_AGEMA_signal_11194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3372 ( .C (clk), .D (new_AGEMA_signal_4756), .Q (new_AGEMA_signal_11197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3375 ( .C (clk), .D (new_AGEMA_signal_4757), .Q (new_AGEMA_signal_11200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3378 ( .C (clk), .D (new_AGEMA_signal_4758), .Q (new_AGEMA_signal_11203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3381 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T1), .Q (new_AGEMA_signal_11206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3384 ( .C (clk), .D (new_AGEMA_signal_4510), .Q (new_AGEMA_signal_11209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3387 ( .C (clk), .D (new_AGEMA_signal_4511), .Q (new_AGEMA_signal_11212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3390 ( .C (clk), .D (new_AGEMA_signal_4512), .Q (new_AGEMA_signal_11215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3393 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T4), .Q (new_AGEMA_signal_11218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3396 ( .C (clk), .D (new_AGEMA_signal_4519), .Q (new_AGEMA_signal_11221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3399 ( .C (clk), .D (new_AGEMA_signal_4520), .Q (new_AGEMA_signal_11224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3402 ( .C (clk), .D (new_AGEMA_signal_4521), .Q (new_AGEMA_signal_11227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3405 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T2), .Q (new_AGEMA_signal_11230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3408 ( .C (clk), .D (new_AGEMA_signal_4513), .Q (new_AGEMA_signal_11233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3411 ( .C (clk), .D (new_AGEMA_signal_4514), .Q (new_AGEMA_signal_11236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3414 ( .C (clk), .D (new_AGEMA_signal_4515), .Q (new_AGEMA_signal_11239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3417 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T6), .Q (new_AGEMA_signal_11242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3420 ( .C (clk), .D (new_AGEMA_signal_4642), .Q (new_AGEMA_signal_11245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3423 ( .C (clk), .D (new_AGEMA_signal_4643), .Q (new_AGEMA_signal_11248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3426 ( .C (clk), .D (new_AGEMA_signal_4644), .Q (new_AGEMA_signal_11251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3429 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T8), .Q (new_AGEMA_signal_11254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3432 ( .C (clk), .D (new_AGEMA_signal_4783), .Q (new_AGEMA_signal_11257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3435 ( .C (clk), .D (new_AGEMA_signal_4784), .Q (new_AGEMA_signal_11260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3438 ( .C (clk), .D (new_AGEMA_signal_4785), .Q (new_AGEMA_signal_11263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3441 ( .C (clk), .D (SubBytesInput[24]), .Q (new_AGEMA_signal_11266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3444 ( .C (clk), .D (new_AGEMA_signal_3562), .Q (new_AGEMA_signal_11269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3447 ( .C (clk), .D (new_AGEMA_signal_3563), .Q (new_AGEMA_signal_11272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3450 ( .C (clk), .D (new_AGEMA_signal_3564), .Q (new_AGEMA_signal_11275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3453 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T16), .Q (new_AGEMA_signal_11278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3456 ( .C (clk), .D (new_AGEMA_signal_4654), .Q (new_AGEMA_signal_11281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3459 ( .C (clk), .D (new_AGEMA_signal_4655), .Q (new_AGEMA_signal_11284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3462 ( .C (clk), .D (new_AGEMA_signal_4656), .Q (new_AGEMA_signal_11287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3465 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T9), .Q (new_AGEMA_signal_11290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3468 ( .C (clk), .D (new_AGEMA_signal_4645), .Q (new_AGEMA_signal_11293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3471 ( .C (clk), .D (new_AGEMA_signal_4646), .Q (new_AGEMA_signal_11296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3474 ( .C (clk), .D (new_AGEMA_signal_4647), .Q (new_AGEMA_signal_11299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3477 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T17), .Q (new_AGEMA_signal_11302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3480 ( .C (clk), .D (new_AGEMA_signal_4792), .Q (new_AGEMA_signal_11305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3483 ( .C (clk), .D (new_AGEMA_signal_4793), .Q (new_AGEMA_signal_11308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3486 ( .C (clk), .D (new_AGEMA_signal_4794), .Q (new_AGEMA_signal_11311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3489 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T15), .Q (new_AGEMA_signal_11314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3492 ( .C (clk), .D (new_AGEMA_signal_4651), .Q (new_AGEMA_signal_11317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3495 ( .C (clk), .D (new_AGEMA_signal_4652), .Q (new_AGEMA_signal_11320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3498 ( .C (clk), .D (new_AGEMA_signal_4653), .Q (new_AGEMA_signal_11323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3501 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T27), .Q (new_AGEMA_signal_11326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3504 ( .C (clk), .D (new_AGEMA_signal_4663), .Q (new_AGEMA_signal_11329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3507 ( .C (clk), .D (new_AGEMA_signal_4664), .Q (new_AGEMA_signal_11332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3510 ( .C (clk), .D (new_AGEMA_signal_4665), .Q (new_AGEMA_signal_11335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3513 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T10), .Q (new_AGEMA_signal_11338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3516 ( .C (clk), .D (new_AGEMA_signal_4786), .Q (new_AGEMA_signal_11341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3519 ( .C (clk), .D (new_AGEMA_signal_4787), .Q (new_AGEMA_signal_11344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3522 ( .C (clk), .D (new_AGEMA_signal_4788), .Q (new_AGEMA_signal_11347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3525 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T13), .Q (new_AGEMA_signal_11350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3528 ( .C (clk), .D (new_AGEMA_signal_4648), .Q (new_AGEMA_signal_11353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3531 ( .C (clk), .D (new_AGEMA_signal_4649), .Q (new_AGEMA_signal_11356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3534 ( .C (clk), .D (new_AGEMA_signal_4650), .Q (new_AGEMA_signal_11359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3537 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T23), .Q (new_AGEMA_signal_11362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3540 ( .C (clk), .D (new_AGEMA_signal_4798), .Q (new_AGEMA_signal_11365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3543 ( .C (clk), .D (new_AGEMA_signal_4799), .Q (new_AGEMA_signal_11368) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3546 ( .C (clk), .D (new_AGEMA_signal_4800), .Q (new_AGEMA_signal_11371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3549 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T19), .Q (new_AGEMA_signal_11374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3552 ( .C (clk), .D (new_AGEMA_signal_4657), .Q (new_AGEMA_signal_11377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3555 ( .C (clk), .D (new_AGEMA_signal_4658), .Q (new_AGEMA_signal_11380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3558 ( .C (clk), .D (new_AGEMA_signal_4659), .Q (new_AGEMA_signal_11383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3561 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T3), .Q (new_AGEMA_signal_11386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3564 ( .C (clk), .D (new_AGEMA_signal_4546), .Q (new_AGEMA_signal_11389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3567 ( .C (clk), .D (new_AGEMA_signal_4547), .Q (new_AGEMA_signal_11392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3570 ( .C (clk), .D (new_AGEMA_signal_4548), .Q (new_AGEMA_signal_11395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3573 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T22), .Q (new_AGEMA_signal_11398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3576 ( .C (clk), .D (new_AGEMA_signal_4660), .Q (new_AGEMA_signal_11401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3579 ( .C (clk), .D (new_AGEMA_signal_4661), .Q (new_AGEMA_signal_11404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3582 ( .C (clk), .D (new_AGEMA_signal_4662), .Q (new_AGEMA_signal_11407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3585 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T20), .Q (new_AGEMA_signal_11410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3588 ( .C (clk), .D (new_AGEMA_signal_4795), .Q (new_AGEMA_signal_11413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3591 ( .C (clk), .D (new_AGEMA_signal_4796), .Q (new_AGEMA_signal_11416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3594 ( .C (clk), .D (new_AGEMA_signal_4797), .Q (new_AGEMA_signal_11419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3597 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T1), .Q (new_AGEMA_signal_11422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3600 ( .C (clk), .D (new_AGEMA_signal_4540), .Q (new_AGEMA_signal_11425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3603 ( .C (clk), .D (new_AGEMA_signal_4541), .Q (new_AGEMA_signal_11428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3606 ( .C (clk), .D (new_AGEMA_signal_4542), .Q (new_AGEMA_signal_11431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3609 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T4), .Q (new_AGEMA_signal_11434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3612 ( .C (clk), .D (new_AGEMA_signal_4549), .Q (new_AGEMA_signal_11437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3615 ( .C (clk), .D (new_AGEMA_signal_4550), .Q (new_AGEMA_signal_11440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3618 ( .C (clk), .D (new_AGEMA_signal_4551), .Q (new_AGEMA_signal_11443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3621 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T2), .Q (new_AGEMA_signal_11446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3624 ( .C (clk), .D (new_AGEMA_signal_4543), .Q (new_AGEMA_signal_11449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3627 ( .C (clk), .D (new_AGEMA_signal_4544), .Q (new_AGEMA_signal_11452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3630 ( .C (clk), .D (new_AGEMA_signal_4545), .Q (new_AGEMA_signal_11455) ) ;
    buf_clk new_AGEMA_reg_buffer_3633 ( .C (clk), .D (MuxMCOut_n5), .Q (new_AGEMA_signal_11458) ) ;
    buf_clk new_AGEMA_reg_buffer_3637 ( .C (clk), .D (LastRoundorDone), .Q (new_AGEMA_signal_11462) ) ;
    buf_clk new_AGEMA_reg_buffer_3641 ( .C (clk), .D (MuxMCOut_n4), .Q (new_AGEMA_signal_11466) ) ;
    buf_clk new_AGEMA_reg_buffer_3645 ( .C (clk), .D (AKSRnotDone), .Q (new_AGEMA_signal_11470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3649 ( .C (clk), .D (ShiftRowsOutput[0]), .Q (new_AGEMA_signal_11474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3653 ( .C (clk), .D (new_AGEMA_signal_2821), .Q (new_AGEMA_signal_11478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3657 ( .C (clk), .D (new_AGEMA_signal_2822), .Q (new_AGEMA_signal_11482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3661 ( .C (clk), .D (new_AGEMA_signal_2823), .Q (new_AGEMA_signal_11486) ) ;
    buf_clk new_AGEMA_reg_buffer_3665 ( .C (clk), .D (MuxRound_n13), .Q (new_AGEMA_signal_11490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3669 ( .C (clk), .D (ShiftRowsOutput[1]), .Q (new_AGEMA_signal_11494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3673 ( .C (clk), .D (new_AGEMA_signal_2830), .Q (new_AGEMA_signal_11498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3677 ( .C (clk), .D (new_AGEMA_signal_2831), .Q (new_AGEMA_signal_11502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3681 ( .C (clk), .D (new_AGEMA_signal_2832), .Q (new_AGEMA_signal_11506) ) ;
    buf_clk new_AGEMA_reg_buffer_3685 ( .C (clk), .D (MuxRound_n14), .Q (new_AGEMA_signal_11510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3689 ( .C (clk), .D (ShiftRowsOutput[2]), .Q (new_AGEMA_signal_11514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3693 ( .C (clk), .D (new_AGEMA_signal_2839), .Q (new_AGEMA_signal_11518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3697 ( .C (clk), .D (new_AGEMA_signal_2840), .Q (new_AGEMA_signal_11522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3701 ( .C (clk), .D (new_AGEMA_signal_2841), .Q (new_AGEMA_signal_11526) ) ;
    buf_clk new_AGEMA_reg_buffer_3705 ( .C (clk), .D (MuxRound_n15), .Q (new_AGEMA_signal_11530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3709 ( .C (clk), .D (ShiftRowsOutput[3]), .Q (new_AGEMA_signal_11534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3713 ( .C (clk), .D (new_AGEMA_signal_2848), .Q (new_AGEMA_signal_11538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3717 ( .C (clk), .D (new_AGEMA_signal_2849), .Q (new_AGEMA_signal_11542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3721 ( .C (clk), .D (new_AGEMA_signal_2850), .Q (new_AGEMA_signal_11546) ) ;
    buf_clk new_AGEMA_reg_buffer_3725 ( .C (clk), .D (MuxRound_n16), .Q (new_AGEMA_signal_11550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3729 ( .C (clk), .D (ShiftRowsOutput[4]), .Q (new_AGEMA_signal_11554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3733 ( .C (clk), .D (new_AGEMA_signal_2857), .Q (new_AGEMA_signal_11558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3737 ( .C (clk), .D (new_AGEMA_signal_2858), .Q (new_AGEMA_signal_11562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3741 ( .C (clk), .D (new_AGEMA_signal_2859), .Q (new_AGEMA_signal_11566) ) ;
    buf_clk new_AGEMA_reg_buffer_3745 ( .C (clk), .D (MuxRound_n17), .Q (new_AGEMA_signal_11570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3749 ( .C (clk), .D (ShiftRowsOutput[5]), .Q (new_AGEMA_signal_11574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3753 ( .C (clk), .D (new_AGEMA_signal_2866), .Q (new_AGEMA_signal_11578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3757 ( .C (clk), .D (new_AGEMA_signal_2867), .Q (new_AGEMA_signal_11582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3761 ( .C (clk), .D (new_AGEMA_signal_2868), .Q (new_AGEMA_signal_11586) ) ;
    buf_clk new_AGEMA_reg_buffer_3765 ( .C (clk), .D (MuxRound_n18), .Q (new_AGEMA_signal_11590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3769 ( .C (clk), .D (ShiftRowsOutput[6]), .Q (new_AGEMA_signal_11594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3773 ( .C (clk), .D (new_AGEMA_signal_2875), .Q (new_AGEMA_signal_11598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3777 ( .C (clk), .D (new_AGEMA_signal_2876), .Q (new_AGEMA_signal_11602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3781 ( .C (clk), .D (new_AGEMA_signal_2877), .Q (new_AGEMA_signal_11606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3785 ( .C (clk), .D (ShiftRowsOutput[7]), .Q (new_AGEMA_signal_11610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3789 ( .C (clk), .D (new_AGEMA_signal_2884), .Q (new_AGEMA_signal_11614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3793 ( .C (clk), .D (new_AGEMA_signal_2885), .Q (new_AGEMA_signal_11618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3797 ( .C (clk), .D (new_AGEMA_signal_2886), .Q (new_AGEMA_signal_11622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3801 ( .C (clk), .D (ShiftRowsOutput[8]), .Q (new_AGEMA_signal_11626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3805 ( .C (clk), .D (new_AGEMA_signal_3217), .Q (new_AGEMA_signal_11630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3809 ( .C (clk), .D (new_AGEMA_signal_3218), .Q (new_AGEMA_signal_11634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3813 ( .C (clk), .D (new_AGEMA_signal_3219), .Q (new_AGEMA_signal_11638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3817 ( .C (clk), .D (ShiftRowsOutput[9]), .Q (new_AGEMA_signal_11642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3821 ( .C (clk), .D (new_AGEMA_signal_3226), .Q (new_AGEMA_signal_11646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3825 ( .C (clk), .D (new_AGEMA_signal_3227), .Q (new_AGEMA_signal_11650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3829 ( .C (clk), .D (new_AGEMA_signal_3228), .Q (new_AGEMA_signal_11654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3833 ( .C (clk), .D (ShiftRowsOutput[10]), .Q (new_AGEMA_signal_11658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3837 ( .C (clk), .D (new_AGEMA_signal_3235), .Q (new_AGEMA_signal_11662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3841 ( .C (clk), .D (new_AGEMA_signal_3236), .Q (new_AGEMA_signal_11666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3845 ( .C (clk), .D (new_AGEMA_signal_3237), .Q (new_AGEMA_signal_11670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3849 ( .C (clk), .D (ShiftRowsOutput[11]), .Q (new_AGEMA_signal_11674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3853 ( .C (clk), .D (new_AGEMA_signal_3244), .Q (new_AGEMA_signal_11678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3857 ( .C (clk), .D (new_AGEMA_signal_3245), .Q (new_AGEMA_signal_11682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3861 ( .C (clk), .D (new_AGEMA_signal_3246), .Q (new_AGEMA_signal_11686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3865 ( .C (clk), .D (ShiftRowsOutput[12]), .Q (new_AGEMA_signal_11690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3869 ( .C (clk), .D (new_AGEMA_signal_3253), .Q (new_AGEMA_signal_11694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3873 ( .C (clk), .D (new_AGEMA_signal_3254), .Q (new_AGEMA_signal_11698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3877 ( .C (clk), .D (new_AGEMA_signal_3255), .Q (new_AGEMA_signal_11702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3881 ( .C (clk), .D (ShiftRowsOutput[13]), .Q (new_AGEMA_signal_11706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3885 ( .C (clk), .D (new_AGEMA_signal_3262), .Q (new_AGEMA_signal_11710) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3889 ( .C (clk), .D (new_AGEMA_signal_3263), .Q (new_AGEMA_signal_11714) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3893 ( .C (clk), .D (new_AGEMA_signal_3264), .Q (new_AGEMA_signal_11718) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3897 ( .C (clk), .D (ShiftRowsOutput[14]), .Q (new_AGEMA_signal_11722) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3901 ( .C (clk), .D (new_AGEMA_signal_3271), .Q (new_AGEMA_signal_11726) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3905 ( .C (clk), .D (new_AGEMA_signal_3272), .Q (new_AGEMA_signal_11730) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3909 ( .C (clk), .D (new_AGEMA_signal_3273), .Q (new_AGEMA_signal_11734) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3913 ( .C (clk), .D (ShiftRowsOutput[15]), .Q (new_AGEMA_signal_11738) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3917 ( .C (clk), .D (new_AGEMA_signal_3280), .Q (new_AGEMA_signal_11742) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3921 ( .C (clk), .D (new_AGEMA_signal_3281), .Q (new_AGEMA_signal_11746) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3925 ( .C (clk), .D (new_AGEMA_signal_3282), .Q (new_AGEMA_signal_11750) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3929 ( .C (clk), .D (ShiftRowsOutput[16]), .Q (new_AGEMA_signal_11754) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3933 ( .C (clk), .D (new_AGEMA_signal_2470), .Q (new_AGEMA_signal_11758) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3937 ( .C (clk), .D (new_AGEMA_signal_2471), .Q (new_AGEMA_signal_11762) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3941 ( .C (clk), .D (new_AGEMA_signal_2472), .Q (new_AGEMA_signal_11766) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3945 ( .C (clk), .D (ShiftRowsOutput[17]), .Q (new_AGEMA_signal_11770) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3949 ( .C (clk), .D (new_AGEMA_signal_2479), .Q (new_AGEMA_signal_11774) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3953 ( .C (clk), .D (new_AGEMA_signal_2480), .Q (new_AGEMA_signal_11778) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3957 ( .C (clk), .D (new_AGEMA_signal_2481), .Q (new_AGEMA_signal_11782) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3961 ( .C (clk), .D (ShiftRowsOutput[18]), .Q (new_AGEMA_signal_11786) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3965 ( .C (clk), .D (new_AGEMA_signal_2488), .Q (new_AGEMA_signal_11790) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3969 ( .C (clk), .D (new_AGEMA_signal_2489), .Q (new_AGEMA_signal_11794) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3973 ( .C (clk), .D (new_AGEMA_signal_2490), .Q (new_AGEMA_signal_11798) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3977 ( .C (clk), .D (ShiftRowsOutput[19]), .Q (new_AGEMA_signal_11802) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3981 ( .C (clk), .D (new_AGEMA_signal_2497), .Q (new_AGEMA_signal_11806) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3985 ( .C (clk), .D (new_AGEMA_signal_2498), .Q (new_AGEMA_signal_11810) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3989 ( .C (clk), .D (new_AGEMA_signal_2499), .Q (new_AGEMA_signal_11814) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3993 ( .C (clk), .D (ShiftRowsOutput[20]), .Q (new_AGEMA_signal_11818) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3997 ( .C (clk), .D (new_AGEMA_signal_2506), .Q (new_AGEMA_signal_11822) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4001 ( .C (clk), .D (new_AGEMA_signal_2507), .Q (new_AGEMA_signal_11826) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4005 ( .C (clk), .D (new_AGEMA_signal_2508), .Q (new_AGEMA_signal_11830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4009 ( .C (clk), .D (ShiftRowsOutput[21]), .Q (new_AGEMA_signal_11834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4013 ( .C (clk), .D (new_AGEMA_signal_2515), .Q (new_AGEMA_signal_11838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4017 ( .C (clk), .D (new_AGEMA_signal_2516), .Q (new_AGEMA_signal_11842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4021 ( .C (clk), .D (new_AGEMA_signal_2517), .Q (new_AGEMA_signal_11846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4025 ( .C (clk), .D (ShiftRowsOutput[22]), .Q (new_AGEMA_signal_11850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4029 ( .C (clk), .D (new_AGEMA_signal_2524), .Q (new_AGEMA_signal_11854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4033 ( .C (clk), .D (new_AGEMA_signal_2525), .Q (new_AGEMA_signal_11858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4037 ( .C (clk), .D (new_AGEMA_signal_2526), .Q (new_AGEMA_signal_11862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4041 ( .C (clk), .D (ShiftRowsOutput[23]), .Q (new_AGEMA_signal_11866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4045 ( .C (clk), .D (new_AGEMA_signal_2533), .Q (new_AGEMA_signal_11870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4049 ( .C (clk), .D (new_AGEMA_signal_2534), .Q (new_AGEMA_signal_11874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4053 ( .C (clk), .D (new_AGEMA_signal_2535), .Q (new_AGEMA_signal_11878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4057 ( .C (clk), .D (ShiftRowsOutput[24]), .Q (new_AGEMA_signal_11882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4061 ( .C (clk), .D (new_AGEMA_signal_2740), .Q (new_AGEMA_signal_11886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4065 ( .C (clk), .D (new_AGEMA_signal_2741), .Q (new_AGEMA_signal_11890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4069 ( .C (clk), .D (new_AGEMA_signal_2742), .Q (new_AGEMA_signal_11894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4073 ( .C (clk), .D (ShiftRowsOutput[25]), .Q (new_AGEMA_signal_11898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4077 ( .C (clk), .D (new_AGEMA_signal_2749), .Q (new_AGEMA_signal_11902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4081 ( .C (clk), .D (new_AGEMA_signal_2750), .Q (new_AGEMA_signal_11906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4085 ( .C (clk), .D (new_AGEMA_signal_2751), .Q (new_AGEMA_signal_11910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4089 ( .C (clk), .D (ShiftRowsOutput[26]), .Q (new_AGEMA_signal_11914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4093 ( .C (clk), .D (new_AGEMA_signal_2758), .Q (new_AGEMA_signal_11918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4097 ( .C (clk), .D (new_AGEMA_signal_2759), .Q (new_AGEMA_signal_11922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4101 ( .C (clk), .D (new_AGEMA_signal_2760), .Q (new_AGEMA_signal_11926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4105 ( .C (clk), .D (ShiftRowsOutput[27]), .Q (new_AGEMA_signal_11930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4109 ( .C (clk), .D (new_AGEMA_signal_2767), .Q (new_AGEMA_signal_11934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4113 ( .C (clk), .D (new_AGEMA_signal_2768), .Q (new_AGEMA_signal_11938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4117 ( .C (clk), .D (new_AGEMA_signal_2769), .Q (new_AGEMA_signal_11942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4121 ( .C (clk), .D (ShiftRowsOutput[28]), .Q (new_AGEMA_signal_11946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4125 ( .C (clk), .D (new_AGEMA_signal_2776), .Q (new_AGEMA_signal_11950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4129 ( .C (clk), .D (new_AGEMA_signal_2777), .Q (new_AGEMA_signal_11954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4133 ( .C (clk), .D (new_AGEMA_signal_2778), .Q (new_AGEMA_signal_11958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4137 ( .C (clk), .D (ShiftRowsOutput[29]), .Q (new_AGEMA_signal_11962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4141 ( .C (clk), .D (new_AGEMA_signal_2785), .Q (new_AGEMA_signal_11966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4145 ( .C (clk), .D (new_AGEMA_signal_2786), .Q (new_AGEMA_signal_11970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4149 ( .C (clk), .D (new_AGEMA_signal_2787), .Q (new_AGEMA_signal_11974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4153 ( .C (clk), .D (ShiftRowsOutput[30]), .Q (new_AGEMA_signal_11978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4157 ( .C (clk), .D (new_AGEMA_signal_2803), .Q (new_AGEMA_signal_11982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4161 ( .C (clk), .D (new_AGEMA_signal_2804), .Q (new_AGEMA_signal_11986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4165 ( .C (clk), .D (new_AGEMA_signal_2805), .Q (new_AGEMA_signal_11990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4169 ( .C (clk), .D (ShiftRowsOutput[31]), .Q (new_AGEMA_signal_11994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4173 ( .C (clk), .D (new_AGEMA_signal_2812), .Q (new_AGEMA_signal_11998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4177 ( .C (clk), .D (new_AGEMA_signal_2813), .Q (new_AGEMA_signal_12002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4181 ( .C (clk), .D (new_AGEMA_signal_2814), .Q (new_AGEMA_signal_12006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4185 ( .C (clk), .D (key_s0[0]), .Q (new_AGEMA_signal_12010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4189 ( .C (clk), .D (key_s1[0]), .Q (new_AGEMA_signal_12014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4193 ( .C (clk), .D (key_s2[0]), .Q (new_AGEMA_signal_12018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4197 ( .C (clk), .D (key_s3[0]), .Q (new_AGEMA_signal_12022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4201 ( .C (clk), .D (key_s0[1]), .Q (new_AGEMA_signal_12026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4205 ( .C (clk), .D (key_s1[1]), .Q (new_AGEMA_signal_12030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4209 ( .C (clk), .D (key_s2[1]), .Q (new_AGEMA_signal_12034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4213 ( .C (clk), .D (key_s3[1]), .Q (new_AGEMA_signal_12038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4217 ( .C (clk), .D (key_s0[2]), .Q (new_AGEMA_signal_12042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4221 ( .C (clk), .D (key_s1[2]), .Q (new_AGEMA_signal_12046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4225 ( .C (clk), .D (key_s2[2]), .Q (new_AGEMA_signal_12050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4229 ( .C (clk), .D (key_s3[2]), .Q (new_AGEMA_signal_12054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4233 ( .C (clk), .D (key_s0[3]), .Q (new_AGEMA_signal_12058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4237 ( .C (clk), .D (key_s1[3]), .Q (new_AGEMA_signal_12062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4241 ( .C (clk), .D (key_s2[3]), .Q (new_AGEMA_signal_12066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4245 ( .C (clk), .D (key_s3[3]), .Q (new_AGEMA_signal_12070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4249 ( .C (clk), .D (key_s0[4]), .Q (new_AGEMA_signal_12074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4253 ( .C (clk), .D (key_s1[4]), .Q (new_AGEMA_signal_12078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4257 ( .C (clk), .D (key_s2[4]), .Q (new_AGEMA_signal_12082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4261 ( .C (clk), .D (key_s3[4]), .Q (new_AGEMA_signal_12086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4265 ( .C (clk), .D (key_s0[5]), .Q (new_AGEMA_signal_12090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4269 ( .C (clk), .D (key_s1[5]), .Q (new_AGEMA_signal_12094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4273 ( .C (clk), .D (key_s2[5]), .Q (new_AGEMA_signal_12098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4277 ( .C (clk), .D (key_s3[5]), .Q (new_AGEMA_signal_12102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4281 ( .C (clk), .D (key_s0[6]), .Q (new_AGEMA_signal_12106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4285 ( .C (clk), .D (key_s1[6]), .Q (new_AGEMA_signal_12110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4289 ( .C (clk), .D (key_s2[6]), .Q (new_AGEMA_signal_12114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4293 ( .C (clk), .D (key_s3[6]), .Q (new_AGEMA_signal_12118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4297 ( .C (clk), .D (key_s0[7]), .Q (new_AGEMA_signal_12122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4301 ( .C (clk), .D (key_s1[7]), .Q (new_AGEMA_signal_12126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4305 ( .C (clk), .D (key_s2[7]), .Q (new_AGEMA_signal_12130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4309 ( .C (clk), .D (key_s3[7]), .Q (new_AGEMA_signal_12134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4313 ( .C (clk), .D (key_s0[8]), .Q (new_AGEMA_signal_12138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4317 ( .C (clk), .D (key_s1[8]), .Q (new_AGEMA_signal_12142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4321 ( .C (clk), .D (key_s2[8]), .Q (new_AGEMA_signal_12146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4325 ( .C (clk), .D (key_s3[8]), .Q (new_AGEMA_signal_12150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4329 ( .C (clk), .D (key_s0[9]), .Q (new_AGEMA_signal_12154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4333 ( .C (clk), .D (key_s1[9]), .Q (new_AGEMA_signal_12158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4337 ( .C (clk), .D (key_s2[9]), .Q (new_AGEMA_signal_12162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4341 ( .C (clk), .D (key_s3[9]), .Q (new_AGEMA_signal_12166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4345 ( .C (clk), .D (key_s0[10]), .Q (new_AGEMA_signal_12170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4349 ( .C (clk), .D (key_s1[10]), .Q (new_AGEMA_signal_12174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4353 ( .C (clk), .D (key_s2[10]), .Q (new_AGEMA_signal_12178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4357 ( .C (clk), .D (key_s3[10]), .Q (new_AGEMA_signal_12182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4361 ( .C (clk), .D (key_s0[11]), .Q (new_AGEMA_signal_12186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4365 ( .C (clk), .D (key_s1[11]), .Q (new_AGEMA_signal_12190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4369 ( .C (clk), .D (key_s2[11]), .Q (new_AGEMA_signal_12194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4373 ( .C (clk), .D (key_s3[11]), .Q (new_AGEMA_signal_12198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4377 ( .C (clk), .D (key_s0[12]), .Q (new_AGEMA_signal_12202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4381 ( .C (clk), .D (key_s1[12]), .Q (new_AGEMA_signal_12206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4385 ( .C (clk), .D (key_s2[12]), .Q (new_AGEMA_signal_12210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4389 ( .C (clk), .D (key_s3[12]), .Q (new_AGEMA_signal_12214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4393 ( .C (clk), .D (key_s0[13]), .Q (new_AGEMA_signal_12218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4397 ( .C (clk), .D (key_s1[13]), .Q (new_AGEMA_signal_12222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4401 ( .C (clk), .D (key_s2[13]), .Q (new_AGEMA_signal_12226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4405 ( .C (clk), .D (key_s3[13]), .Q (new_AGEMA_signal_12230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4409 ( .C (clk), .D (key_s0[14]), .Q (new_AGEMA_signal_12234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4413 ( .C (clk), .D (key_s1[14]), .Q (new_AGEMA_signal_12238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4417 ( .C (clk), .D (key_s2[14]), .Q (new_AGEMA_signal_12242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4421 ( .C (clk), .D (key_s3[14]), .Q (new_AGEMA_signal_12246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4425 ( .C (clk), .D (key_s0[15]), .Q (new_AGEMA_signal_12250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4429 ( .C (clk), .D (key_s1[15]), .Q (new_AGEMA_signal_12254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4433 ( .C (clk), .D (key_s2[15]), .Q (new_AGEMA_signal_12258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4437 ( .C (clk), .D (key_s3[15]), .Q (new_AGEMA_signal_12262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4441 ( .C (clk), .D (key_s0[16]), .Q (new_AGEMA_signal_12266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4445 ( .C (clk), .D (key_s1[16]), .Q (new_AGEMA_signal_12270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4449 ( .C (clk), .D (key_s2[16]), .Q (new_AGEMA_signal_12274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4453 ( .C (clk), .D (key_s3[16]), .Q (new_AGEMA_signal_12278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4457 ( .C (clk), .D (key_s0[17]), .Q (new_AGEMA_signal_12282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4461 ( .C (clk), .D (key_s1[17]), .Q (new_AGEMA_signal_12286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4465 ( .C (clk), .D (key_s2[17]), .Q (new_AGEMA_signal_12290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4469 ( .C (clk), .D (key_s3[17]), .Q (new_AGEMA_signal_12294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4473 ( .C (clk), .D (key_s0[18]), .Q (new_AGEMA_signal_12298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4477 ( .C (clk), .D (key_s1[18]), .Q (new_AGEMA_signal_12302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4481 ( .C (clk), .D (key_s2[18]), .Q (new_AGEMA_signal_12306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4485 ( .C (clk), .D (key_s3[18]), .Q (new_AGEMA_signal_12310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4489 ( .C (clk), .D (key_s0[19]), .Q (new_AGEMA_signal_12314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4493 ( .C (clk), .D (key_s1[19]), .Q (new_AGEMA_signal_12318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4497 ( .C (clk), .D (key_s2[19]), .Q (new_AGEMA_signal_12322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4501 ( .C (clk), .D (key_s3[19]), .Q (new_AGEMA_signal_12326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4505 ( .C (clk), .D (key_s0[20]), .Q (new_AGEMA_signal_12330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4509 ( .C (clk), .D (key_s1[20]), .Q (new_AGEMA_signal_12334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4513 ( .C (clk), .D (key_s2[20]), .Q (new_AGEMA_signal_12338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4517 ( .C (clk), .D (key_s3[20]), .Q (new_AGEMA_signal_12342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4521 ( .C (clk), .D (key_s0[21]), .Q (new_AGEMA_signal_12346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4525 ( .C (clk), .D (key_s1[21]), .Q (new_AGEMA_signal_12350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4529 ( .C (clk), .D (key_s2[21]), .Q (new_AGEMA_signal_12354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4533 ( .C (clk), .D (key_s3[21]), .Q (new_AGEMA_signal_12358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4537 ( .C (clk), .D (key_s0[22]), .Q (new_AGEMA_signal_12362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4541 ( .C (clk), .D (key_s1[22]), .Q (new_AGEMA_signal_12366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4545 ( .C (clk), .D (key_s2[22]), .Q (new_AGEMA_signal_12370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4549 ( .C (clk), .D (key_s3[22]), .Q (new_AGEMA_signal_12374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4553 ( .C (clk), .D (key_s0[23]), .Q (new_AGEMA_signal_12378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4557 ( .C (clk), .D (key_s1[23]), .Q (new_AGEMA_signal_12382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4561 ( .C (clk), .D (key_s2[23]), .Q (new_AGEMA_signal_12386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4565 ( .C (clk), .D (key_s3[23]), .Q (new_AGEMA_signal_12390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4569 ( .C (clk), .D (key_s0[24]), .Q (new_AGEMA_signal_12394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4573 ( .C (clk), .D (key_s1[24]), .Q (new_AGEMA_signal_12398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4577 ( .C (clk), .D (key_s2[24]), .Q (new_AGEMA_signal_12402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4581 ( .C (clk), .D (key_s3[24]), .Q (new_AGEMA_signal_12406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4585 ( .C (clk), .D (key_s0[25]), .Q (new_AGEMA_signal_12410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4589 ( .C (clk), .D (key_s1[25]), .Q (new_AGEMA_signal_12414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4593 ( .C (clk), .D (key_s2[25]), .Q (new_AGEMA_signal_12418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4597 ( .C (clk), .D (key_s3[25]), .Q (new_AGEMA_signal_12422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4601 ( .C (clk), .D (key_s0[26]), .Q (new_AGEMA_signal_12426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4605 ( .C (clk), .D (key_s1[26]), .Q (new_AGEMA_signal_12430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4609 ( .C (clk), .D (key_s2[26]), .Q (new_AGEMA_signal_12434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4613 ( .C (clk), .D (key_s3[26]), .Q (new_AGEMA_signal_12438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4617 ( .C (clk), .D (key_s0[27]), .Q (new_AGEMA_signal_12442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4621 ( .C (clk), .D (key_s1[27]), .Q (new_AGEMA_signal_12446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4625 ( .C (clk), .D (key_s2[27]), .Q (new_AGEMA_signal_12450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4629 ( .C (clk), .D (key_s3[27]), .Q (new_AGEMA_signal_12454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4633 ( .C (clk), .D (key_s0[28]), .Q (new_AGEMA_signal_12458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4637 ( .C (clk), .D (key_s1[28]), .Q (new_AGEMA_signal_12462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4641 ( .C (clk), .D (key_s2[28]), .Q (new_AGEMA_signal_12466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4645 ( .C (clk), .D (key_s3[28]), .Q (new_AGEMA_signal_12470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4649 ( .C (clk), .D (key_s0[29]), .Q (new_AGEMA_signal_12474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4653 ( .C (clk), .D (key_s1[29]), .Q (new_AGEMA_signal_12478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4657 ( .C (clk), .D (key_s2[29]), .Q (new_AGEMA_signal_12482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4661 ( .C (clk), .D (key_s3[29]), .Q (new_AGEMA_signal_12486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4665 ( .C (clk), .D (key_s0[30]), .Q (new_AGEMA_signal_12490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4669 ( .C (clk), .D (key_s1[30]), .Q (new_AGEMA_signal_12494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4673 ( .C (clk), .D (key_s2[30]), .Q (new_AGEMA_signal_12498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4677 ( .C (clk), .D (key_s3[30]), .Q (new_AGEMA_signal_12502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4681 ( .C (clk), .D (key_s0[31]), .Q (new_AGEMA_signal_12506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4685 ( .C (clk), .D (key_s1[31]), .Q (new_AGEMA_signal_12510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4689 ( .C (clk), .D (key_s2[31]), .Q (new_AGEMA_signal_12514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4693 ( .C (clk), .D (key_s3[31]), .Q (new_AGEMA_signal_12518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4697 ( .C (clk), .D (key_s0[32]), .Q (new_AGEMA_signal_12522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4701 ( .C (clk), .D (key_s1[32]), .Q (new_AGEMA_signal_12526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4705 ( .C (clk), .D (key_s2[32]), .Q (new_AGEMA_signal_12530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4709 ( .C (clk), .D (key_s3[32]), .Q (new_AGEMA_signal_12534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4713 ( .C (clk), .D (key_s0[33]), .Q (new_AGEMA_signal_12538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4717 ( .C (clk), .D (key_s1[33]), .Q (new_AGEMA_signal_12542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4721 ( .C (clk), .D (key_s2[33]), .Q (new_AGEMA_signal_12546) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4725 ( .C (clk), .D (key_s3[33]), .Q (new_AGEMA_signal_12550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4729 ( .C (clk), .D (key_s0[34]), .Q (new_AGEMA_signal_12554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4733 ( .C (clk), .D (key_s1[34]), .Q (new_AGEMA_signal_12558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4737 ( .C (clk), .D (key_s2[34]), .Q (new_AGEMA_signal_12562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4741 ( .C (clk), .D (key_s3[34]), .Q (new_AGEMA_signal_12566) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4745 ( .C (clk), .D (key_s0[35]), .Q (new_AGEMA_signal_12570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4749 ( .C (clk), .D (key_s1[35]), .Q (new_AGEMA_signal_12574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4753 ( .C (clk), .D (key_s2[35]), .Q (new_AGEMA_signal_12578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4757 ( .C (clk), .D (key_s3[35]), .Q (new_AGEMA_signal_12582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4761 ( .C (clk), .D (key_s0[36]), .Q (new_AGEMA_signal_12586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4765 ( .C (clk), .D (key_s1[36]), .Q (new_AGEMA_signal_12590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4769 ( .C (clk), .D (key_s2[36]), .Q (new_AGEMA_signal_12594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4773 ( .C (clk), .D (key_s3[36]), .Q (new_AGEMA_signal_12598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4777 ( .C (clk), .D (key_s0[37]), .Q (new_AGEMA_signal_12602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4781 ( .C (clk), .D (key_s1[37]), .Q (new_AGEMA_signal_12606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4785 ( .C (clk), .D (key_s2[37]), .Q (new_AGEMA_signal_12610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4789 ( .C (clk), .D (key_s3[37]), .Q (new_AGEMA_signal_12614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4793 ( .C (clk), .D (key_s0[38]), .Q (new_AGEMA_signal_12618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4797 ( .C (clk), .D (key_s1[38]), .Q (new_AGEMA_signal_12622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4801 ( .C (clk), .D (key_s2[38]), .Q (new_AGEMA_signal_12626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4805 ( .C (clk), .D (key_s3[38]), .Q (new_AGEMA_signal_12630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4809 ( .C (clk), .D (key_s0[39]), .Q (new_AGEMA_signal_12634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4813 ( .C (clk), .D (key_s1[39]), .Q (new_AGEMA_signal_12638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4817 ( .C (clk), .D (key_s2[39]), .Q (new_AGEMA_signal_12642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4821 ( .C (clk), .D (key_s3[39]), .Q (new_AGEMA_signal_12646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4825 ( .C (clk), .D (key_s0[40]), .Q (new_AGEMA_signal_12650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4829 ( .C (clk), .D (key_s1[40]), .Q (new_AGEMA_signal_12654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4833 ( .C (clk), .D (key_s2[40]), .Q (new_AGEMA_signal_12658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4837 ( .C (clk), .D (key_s3[40]), .Q (new_AGEMA_signal_12662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4841 ( .C (clk), .D (key_s0[41]), .Q (new_AGEMA_signal_12666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4845 ( .C (clk), .D (key_s1[41]), .Q (new_AGEMA_signal_12670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4849 ( .C (clk), .D (key_s2[41]), .Q (new_AGEMA_signal_12674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4853 ( .C (clk), .D (key_s3[41]), .Q (new_AGEMA_signal_12678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4857 ( .C (clk), .D (key_s0[42]), .Q (new_AGEMA_signal_12682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4861 ( .C (clk), .D (key_s1[42]), .Q (new_AGEMA_signal_12686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4865 ( .C (clk), .D (key_s2[42]), .Q (new_AGEMA_signal_12690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4869 ( .C (clk), .D (key_s3[42]), .Q (new_AGEMA_signal_12694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4873 ( .C (clk), .D (key_s0[43]), .Q (new_AGEMA_signal_12698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4877 ( .C (clk), .D (key_s1[43]), .Q (new_AGEMA_signal_12702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4881 ( .C (clk), .D (key_s2[43]), .Q (new_AGEMA_signal_12706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4885 ( .C (clk), .D (key_s3[43]), .Q (new_AGEMA_signal_12710) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4889 ( .C (clk), .D (key_s0[44]), .Q (new_AGEMA_signal_12714) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4893 ( .C (clk), .D (key_s1[44]), .Q (new_AGEMA_signal_12718) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4897 ( .C (clk), .D (key_s2[44]), .Q (new_AGEMA_signal_12722) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4901 ( .C (clk), .D (key_s3[44]), .Q (new_AGEMA_signal_12726) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4905 ( .C (clk), .D (key_s0[45]), .Q (new_AGEMA_signal_12730) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4909 ( .C (clk), .D (key_s1[45]), .Q (new_AGEMA_signal_12734) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4913 ( .C (clk), .D (key_s2[45]), .Q (new_AGEMA_signal_12738) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4917 ( .C (clk), .D (key_s3[45]), .Q (new_AGEMA_signal_12742) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4921 ( .C (clk), .D (key_s0[46]), .Q (new_AGEMA_signal_12746) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4925 ( .C (clk), .D (key_s1[46]), .Q (new_AGEMA_signal_12750) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4929 ( .C (clk), .D (key_s2[46]), .Q (new_AGEMA_signal_12754) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4933 ( .C (clk), .D (key_s3[46]), .Q (new_AGEMA_signal_12758) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4937 ( .C (clk), .D (key_s0[47]), .Q (new_AGEMA_signal_12762) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4941 ( .C (clk), .D (key_s1[47]), .Q (new_AGEMA_signal_12766) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4945 ( .C (clk), .D (key_s2[47]), .Q (new_AGEMA_signal_12770) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4949 ( .C (clk), .D (key_s3[47]), .Q (new_AGEMA_signal_12774) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4953 ( .C (clk), .D (key_s0[48]), .Q (new_AGEMA_signal_12778) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4957 ( .C (clk), .D (key_s1[48]), .Q (new_AGEMA_signal_12782) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4961 ( .C (clk), .D (key_s2[48]), .Q (new_AGEMA_signal_12786) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4965 ( .C (clk), .D (key_s3[48]), .Q (new_AGEMA_signal_12790) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4969 ( .C (clk), .D (key_s0[49]), .Q (new_AGEMA_signal_12794) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4973 ( .C (clk), .D (key_s1[49]), .Q (new_AGEMA_signal_12798) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4977 ( .C (clk), .D (key_s2[49]), .Q (new_AGEMA_signal_12802) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4981 ( .C (clk), .D (key_s3[49]), .Q (new_AGEMA_signal_12806) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4985 ( .C (clk), .D (key_s0[50]), .Q (new_AGEMA_signal_12810) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4989 ( .C (clk), .D (key_s1[50]), .Q (new_AGEMA_signal_12814) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4993 ( .C (clk), .D (key_s2[50]), .Q (new_AGEMA_signal_12818) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4997 ( .C (clk), .D (key_s3[50]), .Q (new_AGEMA_signal_12822) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5001 ( .C (clk), .D (key_s0[51]), .Q (new_AGEMA_signal_12826) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5005 ( .C (clk), .D (key_s1[51]), .Q (new_AGEMA_signal_12830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5009 ( .C (clk), .D (key_s2[51]), .Q (new_AGEMA_signal_12834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5013 ( .C (clk), .D (key_s3[51]), .Q (new_AGEMA_signal_12838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5017 ( .C (clk), .D (key_s0[52]), .Q (new_AGEMA_signal_12842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5021 ( .C (clk), .D (key_s1[52]), .Q (new_AGEMA_signal_12846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5025 ( .C (clk), .D (key_s2[52]), .Q (new_AGEMA_signal_12850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5029 ( .C (clk), .D (key_s3[52]), .Q (new_AGEMA_signal_12854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5033 ( .C (clk), .D (key_s0[53]), .Q (new_AGEMA_signal_12858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5037 ( .C (clk), .D (key_s1[53]), .Q (new_AGEMA_signal_12862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5041 ( .C (clk), .D (key_s2[53]), .Q (new_AGEMA_signal_12866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5045 ( .C (clk), .D (key_s3[53]), .Q (new_AGEMA_signal_12870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5049 ( .C (clk), .D (key_s0[54]), .Q (new_AGEMA_signal_12874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5053 ( .C (clk), .D (key_s1[54]), .Q (new_AGEMA_signal_12878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5057 ( .C (clk), .D (key_s2[54]), .Q (new_AGEMA_signal_12882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5061 ( .C (clk), .D (key_s3[54]), .Q (new_AGEMA_signal_12886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5065 ( .C (clk), .D (key_s0[55]), .Q (new_AGEMA_signal_12890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5069 ( .C (clk), .D (key_s1[55]), .Q (new_AGEMA_signal_12894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5073 ( .C (clk), .D (key_s2[55]), .Q (new_AGEMA_signal_12898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5077 ( .C (clk), .D (key_s3[55]), .Q (new_AGEMA_signal_12902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5081 ( .C (clk), .D (key_s0[56]), .Q (new_AGEMA_signal_12906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5085 ( .C (clk), .D (key_s1[56]), .Q (new_AGEMA_signal_12910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5089 ( .C (clk), .D (key_s2[56]), .Q (new_AGEMA_signal_12914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5093 ( .C (clk), .D (key_s3[56]), .Q (new_AGEMA_signal_12918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5097 ( .C (clk), .D (key_s0[57]), .Q (new_AGEMA_signal_12922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5101 ( .C (clk), .D (key_s1[57]), .Q (new_AGEMA_signal_12926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5105 ( .C (clk), .D (key_s2[57]), .Q (new_AGEMA_signal_12930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5109 ( .C (clk), .D (key_s3[57]), .Q (new_AGEMA_signal_12934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5113 ( .C (clk), .D (key_s0[58]), .Q (new_AGEMA_signal_12938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5117 ( .C (clk), .D (key_s1[58]), .Q (new_AGEMA_signal_12942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5121 ( .C (clk), .D (key_s2[58]), .Q (new_AGEMA_signal_12946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5125 ( .C (clk), .D (key_s3[58]), .Q (new_AGEMA_signal_12950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5129 ( .C (clk), .D (key_s0[59]), .Q (new_AGEMA_signal_12954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5133 ( .C (clk), .D (key_s1[59]), .Q (new_AGEMA_signal_12958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5137 ( .C (clk), .D (key_s2[59]), .Q (new_AGEMA_signal_12962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5141 ( .C (clk), .D (key_s3[59]), .Q (new_AGEMA_signal_12966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5145 ( .C (clk), .D (key_s0[60]), .Q (new_AGEMA_signal_12970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5149 ( .C (clk), .D (key_s1[60]), .Q (new_AGEMA_signal_12974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5153 ( .C (clk), .D (key_s2[60]), .Q (new_AGEMA_signal_12978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5157 ( .C (clk), .D (key_s3[60]), .Q (new_AGEMA_signal_12982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5161 ( .C (clk), .D (key_s0[61]), .Q (new_AGEMA_signal_12986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5165 ( .C (clk), .D (key_s1[61]), .Q (new_AGEMA_signal_12990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5169 ( .C (clk), .D (key_s2[61]), .Q (new_AGEMA_signal_12994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5173 ( .C (clk), .D (key_s3[61]), .Q (new_AGEMA_signal_12998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5177 ( .C (clk), .D (key_s0[62]), .Q (new_AGEMA_signal_13002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5181 ( .C (clk), .D (key_s1[62]), .Q (new_AGEMA_signal_13006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5185 ( .C (clk), .D (key_s2[62]), .Q (new_AGEMA_signal_13010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5189 ( .C (clk), .D (key_s3[62]), .Q (new_AGEMA_signal_13014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5193 ( .C (clk), .D (key_s0[63]), .Q (new_AGEMA_signal_13018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5197 ( .C (clk), .D (key_s1[63]), .Q (new_AGEMA_signal_13022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5201 ( .C (clk), .D (key_s2[63]), .Q (new_AGEMA_signal_13026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5205 ( .C (clk), .D (key_s3[63]), .Q (new_AGEMA_signal_13030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5209 ( .C (clk), .D (key_s0[64]), .Q (new_AGEMA_signal_13034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5213 ( .C (clk), .D (key_s1[64]), .Q (new_AGEMA_signal_13038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5217 ( .C (clk), .D (key_s2[64]), .Q (new_AGEMA_signal_13042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5221 ( .C (clk), .D (key_s3[64]), .Q (new_AGEMA_signal_13046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5225 ( .C (clk), .D (key_s0[65]), .Q (new_AGEMA_signal_13050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5229 ( .C (clk), .D (key_s1[65]), .Q (new_AGEMA_signal_13054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5233 ( .C (clk), .D (key_s2[65]), .Q (new_AGEMA_signal_13058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5237 ( .C (clk), .D (key_s3[65]), .Q (new_AGEMA_signal_13062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5241 ( .C (clk), .D (key_s0[66]), .Q (new_AGEMA_signal_13066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5245 ( .C (clk), .D (key_s1[66]), .Q (new_AGEMA_signal_13070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5249 ( .C (clk), .D (key_s2[66]), .Q (new_AGEMA_signal_13074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5253 ( .C (clk), .D (key_s3[66]), .Q (new_AGEMA_signal_13078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5257 ( .C (clk), .D (key_s0[67]), .Q (new_AGEMA_signal_13082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5261 ( .C (clk), .D (key_s1[67]), .Q (new_AGEMA_signal_13086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5265 ( .C (clk), .D (key_s2[67]), .Q (new_AGEMA_signal_13090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5269 ( .C (clk), .D (key_s3[67]), .Q (new_AGEMA_signal_13094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5273 ( .C (clk), .D (key_s0[68]), .Q (new_AGEMA_signal_13098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5277 ( .C (clk), .D (key_s1[68]), .Q (new_AGEMA_signal_13102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5281 ( .C (clk), .D (key_s2[68]), .Q (new_AGEMA_signal_13106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5285 ( .C (clk), .D (key_s3[68]), .Q (new_AGEMA_signal_13110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5289 ( .C (clk), .D (key_s0[69]), .Q (new_AGEMA_signal_13114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5293 ( .C (clk), .D (key_s1[69]), .Q (new_AGEMA_signal_13118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5297 ( .C (clk), .D (key_s2[69]), .Q (new_AGEMA_signal_13122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5301 ( .C (clk), .D (key_s3[69]), .Q (new_AGEMA_signal_13126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5305 ( .C (clk), .D (key_s0[70]), .Q (new_AGEMA_signal_13130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5309 ( .C (clk), .D (key_s1[70]), .Q (new_AGEMA_signal_13134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5313 ( .C (clk), .D (key_s2[70]), .Q (new_AGEMA_signal_13138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5317 ( .C (clk), .D (key_s3[70]), .Q (new_AGEMA_signal_13142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5321 ( .C (clk), .D (key_s0[71]), .Q (new_AGEMA_signal_13146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5325 ( .C (clk), .D (key_s1[71]), .Q (new_AGEMA_signal_13150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5329 ( .C (clk), .D (key_s2[71]), .Q (new_AGEMA_signal_13154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5333 ( .C (clk), .D (key_s3[71]), .Q (new_AGEMA_signal_13158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5337 ( .C (clk), .D (key_s0[72]), .Q (new_AGEMA_signal_13162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5341 ( .C (clk), .D (key_s1[72]), .Q (new_AGEMA_signal_13166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5345 ( .C (clk), .D (key_s2[72]), .Q (new_AGEMA_signal_13170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5349 ( .C (clk), .D (key_s3[72]), .Q (new_AGEMA_signal_13174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5353 ( .C (clk), .D (key_s0[73]), .Q (new_AGEMA_signal_13178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5357 ( .C (clk), .D (key_s1[73]), .Q (new_AGEMA_signal_13182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5361 ( .C (clk), .D (key_s2[73]), .Q (new_AGEMA_signal_13186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5365 ( .C (clk), .D (key_s3[73]), .Q (new_AGEMA_signal_13190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5369 ( .C (clk), .D (key_s0[74]), .Q (new_AGEMA_signal_13194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5373 ( .C (clk), .D (key_s1[74]), .Q (new_AGEMA_signal_13198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5377 ( .C (clk), .D (key_s2[74]), .Q (new_AGEMA_signal_13202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5381 ( .C (clk), .D (key_s3[74]), .Q (new_AGEMA_signal_13206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5385 ( .C (clk), .D (key_s0[75]), .Q (new_AGEMA_signal_13210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5389 ( .C (clk), .D (key_s1[75]), .Q (new_AGEMA_signal_13214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5393 ( .C (clk), .D (key_s2[75]), .Q (new_AGEMA_signal_13218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5397 ( .C (clk), .D (key_s3[75]), .Q (new_AGEMA_signal_13222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5401 ( .C (clk), .D (key_s0[76]), .Q (new_AGEMA_signal_13226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5405 ( .C (clk), .D (key_s1[76]), .Q (new_AGEMA_signal_13230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5409 ( .C (clk), .D (key_s2[76]), .Q (new_AGEMA_signal_13234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5413 ( .C (clk), .D (key_s3[76]), .Q (new_AGEMA_signal_13238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5417 ( .C (clk), .D (key_s0[77]), .Q (new_AGEMA_signal_13242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5421 ( .C (clk), .D (key_s1[77]), .Q (new_AGEMA_signal_13246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5425 ( .C (clk), .D (key_s2[77]), .Q (new_AGEMA_signal_13250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5429 ( .C (clk), .D (key_s3[77]), .Q (new_AGEMA_signal_13254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5433 ( .C (clk), .D (key_s0[78]), .Q (new_AGEMA_signal_13258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5437 ( .C (clk), .D (key_s1[78]), .Q (new_AGEMA_signal_13262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5441 ( .C (clk), .D (key_s2[78]), .Q (new_AGEMA_signal_13266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5445 ( .C (clk), .D (key_s3[78]), .Q (new_AGEMA_signal_13270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5449 ( .C (clk), .D (key_s0[79]), .Q (new_AGEMA_signal_13274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5453 ( .C (clk), .D (key_s1[79]), .Q (new_AGEMA_signal_13278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5457 ( .C (clk), .D (key_s2[79]), .Q (new_AGEMA_signal_13282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5461 ( .C (clk), .D (key_s3[79]), .Q (new_AGEMA_signal_13286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5465 ( .C (clk), .D (key_s0[80]), .Q (new_AGEMA_signal_13290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5469 ( .C (clk), .D (key_s1[80]), .Q (new_AGEMA_signal_13294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5473 ( .C (clk), .D (key_s2[80]), .Q (new_AGEMA_signal_13298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5477 ( .C (clk), .D (key_s3[80]), .Q (new_AGEMA_signal_13302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5481 ( .C (clk), .D (key_s0[81]), .Q (new_AGEMA_signal_13306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5485 ( .C (clk), .D (key_s1[81]), .Q (new_AGEMA_signal_13310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5489 ( .C (clk), .D (key_s2[81]), .Q (new_AGEMA_signal_13314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5493 ( .C (clk), .D (key_s3[81]), .Q (new_AGEMA_signal_13318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5497 ( .C (clk), .D (key_s0[82]), .Q (new_AGEMA_signal_13322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5501 ( .C (clk), .D (key_s1[82]), .Q (new_AGEMA_signal_13326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5505 ( .C (clk), .D (key_s2[82]), .Q (new_AGEMA_signal_13330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5509 ( .C (clk), .D (key_s3[82]), .Q (new_AGEMA_signal_13334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5513 ( .C (clk), .D (key_s0[83]), .Q (new_AGEMA_signal_13338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5517 ( .C (clk), .D (key_s1[83]), .Q (new_AGEMA_signal_13342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5521 ( .C (clk), .D (key_s2[83]), .Q (new_AGEMA_signal_13346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5525 ( .C (clk), .D (key_s3[83]), .Q (new_AGEMA_signal_13350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5529 ( .C (clk), .D (key_s0[84]), .Q (new_AGEMA_signal_13354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5533 ( .C (clk), .D (key_s1[84]), .Q (new_AGEMA_signal_13358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5537 ( .C (clk), .D (key_s2[84]), .Q (new_AGEMA_signal_13362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5541 ( .C (clk), .D (key_s3[84]), .Q (new_AGEMA_signal_13366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5545 ( .C (clk), .D (key_s0[85]), .Q (new_AGEMA_signal_13370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5549 ( .C (clk), .D (key_s1[85]), .Q (new_AGEMA_signal_13374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5553 ( .C (clk), .D (key_s2[85]), .Q (new_AGEMA_signal_13378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5557 ( .C (clk), .D (key_s3[85]), .Q (new_AGEMA_signal_13382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5561 ( .C (clk), .D (key_s0[86]), .Q (new_AGEMA_signal_13386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5565 ( .C (clk), .D (key_s1[86]), .Q (new_AGEMA_signal_13390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5569 ( .C (clk), .D (key_s2[86]), .Q (new_AGEMA_signal_13394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5573 ( .C (clk), .D (key_s3[86]), .Q (new_AGEMA_signal_13398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5577 ( .C (clk), .D (key_s0[87]), .Q (new_AGEMA_signal_13402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5581 ( .C (clk), .D (key_s1[87]), .Q (new_AGEMA_signal_13406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5585 ( .C (clk), .D (key_s2[87]), .Q (new_AGEMA_signal_13410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5589 ( .C (clk), .D (key_s3[87]), .Q (new_AGEMA_signal_13414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5593 ( .C (clk), .D (key_s0[88]), .Q (new_AGEMA_signal_13418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5597 ( .C (clk), .D (key_s1[88]), .Q (new_AGEMA_signal_13422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5601 ( .C (clk), .D (key_s2[88]), .Q (new_AGEMA_signal_13426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5605 ( .C (clk), .D (key_s3[88]), .Q (new_AGEMA_signal_13430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5609 ( .C (clk), .D (key_s0[89]), .Q (new_AGEMA_signal_13434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5613 ( .C (clk), .D (key_s1[89]), .Q (new_AGEMA_signal_13438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5617 ( .C (clk), .D (key_s2[89]), .Q (new_AGEMA_signal_13442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5621 ( .C (clk), .D (key_s3[89]), .Q (new_AGEMA_signal_13446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5625 ( .C (clk), .D (key_s0[90]), .Q (new_AGEMA_signal_13450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5629 ( .C (clk), .D (key_s1[90]), .Q (new_AGEMA_signal_13454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5633 ( .C (clk), .D (key_s2[90]), .Q (new_AGEMA_signal_13458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5637 ( .C (clk), .D (key_s3[90]), .Q (new_AGEMA_signal_13462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5641 ( .C (clk), .D (key_s0[91]), .Q (new_AGEMA_signal_13466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5645 ( .C (clk), .D (key_s1[91]), .Q (new_AGEMA_signal_13470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5649 ( .C (clk), .D (key_s2[91]), .Q (new_AGEMA_signal_13474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5653 ( .C (clk), .D (key_s3[91]), .Q (new_AGEMA_signal_13478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5657 ( .C (clk), .D (key_s0[92]), .Q (new_AGEMA_signal_13482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5661 ( .C (clk), .D (key_s1[92]), .Q (new_AGEMA_signal_13486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5665 ( .C (clk), .D (key_s2[92]), .Q (new_AGEMA_signal_13490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5669 ( .C (clk), .D (key_s3[92]), .Q (new_AGEMA_signal_13494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5673 ( .C (clk), .D (key_s0[93]), .Q (new_AGEMA_signal_13498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5677 ( .C (clk), .D (key_s1[93]), .Q (new_AGEMA_signal_13502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5681 ( .C (clk), .D (key_s2[93]), .Q (new_AGEMA_signal_13506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5685 ( .C (clk), .D (key_s3[93]), .Q (new_AGEMA_signal_13510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5689 ( .C (clk), .D (key_s0[94]), .Q (new_AGEMA_signal_13514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5693 ( .C (clk), .D (key_s1[94]), .Q (new_AGEMA_signal_13518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5697 ( .C (clk), .D (key_s2[94]), .Q (new_AGEMA_signal_13522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5701 ( .C (clk), .D (key_s3[94]), .Q (new_AGEMA_signal_13526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5705 ( .C (clk), .D (key_s0[95]), .Q (new_AGEMA_signal_13530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5709 ( .C (clk), .D (key_s1[95]), .Q (new_AGEMA_signal_13534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5713 ( .C (clk), .D (key_s2[95]), .Q (new_AGEMA_signal_13538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5717 ( .C (clk), .D (key_s3[95]), .Q (new_AGEMA_signal_13542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5721 ( .C (clk), .D (key_s0[96]), .Q (new_AGEMA_signal_13546) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5725 ( .C (clk), .D (key_s1[96]), .Q (new_AGEMA_signal_13550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5729 ( .C (clk), .D (key_s2[96]), .Q (new_AGEMA_signal_13554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5733 ( .C (clk), .D (key_s3[96]), .Q (new_AGEMA_signal_13558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5737 ( .C (clk), .D (key_s0[97]), .Q (new_AGEMA_signal_13562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5741 ( .C (clk), .D (key_s1[97]), .Q (new_AGEMA_signal_13566) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5745 ( .C (clk), .D (key_s2[97]), .Q (new_AGEMA_signal_13570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5749 ( .C (clk), .D (key_s3[97]), .Q (new_AGEMA_signal_13574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5753 ( .C (clk), .D (key_s0[98]), .Q (new_AGEMA_signal_13578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5757 ( .C (clk), .D (key_s1[98]), .Q (new_AGEMA_signal_13582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5761 ( .C (clk), .D (key_s2[98]), .Q (new_AGEMA_signal_13586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5765 ( .C (clk), .D (key_s3[98]), .Q (new_AGEMA_signal_13590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5769 ( .C (clk), .D (key_s0[99]), .Q (new_AGEMA_signal_13594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5773 ( .C (clk), .D (key_s1[99]), .Q (new_AGEMA_signal_13598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5777 ( .C (clk), .D (key_s2[99]), .Q (new_AGEMA_signal_13602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5781 ( .C (clk), .D (key_s3[99]), .Q (new_AGEMA_signal_13606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5785 ( .C (clk), .D (key_s0[100]), .Q (new_AGEMA_signal_13610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5789 ( .C (clk), .D (key_s1[100]), .Q (new_AGEMA_signal_13614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5793 ( .C (clk), .D (key_s2[100]), .Q (new_AGEMA_signal_13618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5797 ( .C (clk), .D (key_s3[100]), .Q (new_AGEMA_signal_13622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5801 ( .C (clk), .D (key_s0[101]), .Q (new_AGEMA_signal_13626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5805 ( .C (clk), .D (key_s1[101]), .Q (new_AGEMA_signal_13630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5809 ( .C (clk), .D (key_s2[101]), .Q (new_AGEMA_signal_13634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5813 ( .C (clk), .D (key_s3[101]), .Q (new_AGEMA_signal_13638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5817 ( .C (clk), .D (key_s0[102]), .Q (new_AGEMA_signal_13642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5821 ( .C (clk), .D (key_s1[102]), .Q (new_AGEMA_signal_13646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5825 ( .C (clk), .D (key_s2[102]), .Q (new_AGEMA_signal_13650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5829 ( .C (clk), .D (key_s3[102]), .Q (new_AGEMA_signal_13654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5833 ( .C (clk), .D (key_s0[103]), .Q (new_AGEMA_signal_13658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5837 ( .C (clk), .D (key_s1[103]), .Q (new_AGEMA_signal_13662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5841 ( .C (clk), .D (key_s2[103]), .Q (new_AGEMA_signal_13666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5845 ( .C (clk), .D (key_s3[103]), .Q (new_AGEMA_signal_13670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5849 ( .C (clk), .D (key_s0[104]), .Q (new_AGEMA_signal_13674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5853 ( .C (clk), .D (key_s1[104]), .Q (new_AGEMA_signal_13678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5857 ( .C (clk), .D (key_s2[104]), .Q (new_AGEMA_signal_13682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5861 ( .C (clk), .D (key_s3[104]), .Q (new_AGEMA_signal_13686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5865 ( .C (clk), .D (key_s0[105]), .Q (new_AGEMA_signal_13690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5869 ( .C (clk), .D (key_s1[105]), .Q (new_AGEMA_signal_13694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5873 ( .C (clk), .D (key_s2[105]), .Q (new_AGEMA_signal_13698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5877 ( .C (clk), .D (key_s3[105]), .Q (new_AGEMA_signal_13702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5881 ( .C (clk), .D (key_s0[106]), .Q (new_AGEMA_signal_13706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5885 ( .C (clk), .D (key_s1[106]), .Q (new_AGEMA_signal_13710) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5889 ( .C (clk), .D (key_s2[106]), .Q (new_AGEMA_signal_13714) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5893 ( .C (clk), .D (key_s3[106]), .Q (new_AGEMA_signal_13718) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5897 ( .C (clk), .D (key_s0[107]), .Q (new_AGEMA_signal_13722) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5901 ( .C (clk), .D (key_s1[107]), .Q (new_AGEMA_signal_13726) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5905 ( .C (clk), .D (key_s2[107]), .Q (new_AGEMA_signal_13730) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5909 ( .C (clk), .D (key_s3[107]), .Q (new_AGEMA_signal_13734) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5913 ( .C (clk), .D (key_s0[108]), .Q (new_AGEMA_signal_13738) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5917 ( .C (clk), .D (key_s1[108]), .Q (new_AGEMA_signal_13742) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5921 ( .C (clk), .D (key_s2[108]), .Q (new_AGEMA_signal_13746) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5925 ( .C (clk), .D (key_s3[108]), .Q (new_AGEMA_signal_13750) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5929 ( .C (clk), .D (key_s0[109]), .Q (new_AGEMA_signal_13754) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5933 ( .C (clk), .D (key_s1[109]), .Q (new_AGEMA_signal_13758) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5937 ( .C (clk), .D (key_s2[109]), .Q (new_AGEMA_signal_13762) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5941 ( .C (clk), .D (key_s3[109]), .Q (new_AGEMA_signal_13766) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5945 ( .C (clk), .D (key_s0[110]), .Q (new_AGEMA_signal_13770) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5949 ( .C (clk), .D (key_s1[110]), .Q (new_AGEMA_signal_13774) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5953 ( .C (clk), .D (key_s2[110]), .Q (new_AGEMA_signal_13778) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5957 ( .C (clk), .D (key_s3[110]), .Q (new_AGEMA_signal_13782) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5961 ( .C (clk), .D (key_s0[111]), .Q (new_AGEMA_signal_13786) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5965 ( .C (clk), .D (key_s1[111]), .Q (new_AGEMA_signal_13790) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5969 ( .C (clk), .D (key_s2[111]), .Q (new_AGEMA_signal_13794) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5973 ( .C (clk), .D (key_s3[111]), .Q (new_AGEMA_signal_13798) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5977 ( .C (clk), .D (key_s0[112]), .Q (new_AGEMA_signal_13802) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5981 ( .C (clk), .D (key_s1[112]), .Q (new_AGEMA_signal_13806) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5985 ( .C (clk), .D (key_s2[112]), .Q (new_AGEMA_signal_13810) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5989 ( .C (clk), .D (key_s3[112]), .Q (new_AGEMA_signal_13814) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5993 ( .C (clk), .D (key_s0[113]), .Q (new_AGEMA_signal_13818) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5997 ( .C (clk), .D (key_s1[113]), .Q (new_AGEMA_signal_13822) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6001 ( .C (clk), .D (key_s2[113]), .Q (new_AGEMA_signal_13826) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6005 ( .C (clk), .D (key_s3[113]), .Q (new_AGEMA_signal_13830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6009 ( .C (clk), .D (key_s0[114]), .Q (new_AGEMA_signal_13834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6013 ( .C (clk), .D (key_s1[114]), .Q (new_AGEMA_signal_13838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6017 ( .C (clk), .D (key_s2[114]), .Q (new_AGEMA_signal_13842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6021 ( .C (clk), .D (key_s3[114]), .Q (new_AGEMA_signal_13846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6025 ( .C (clk), .D (key_s0[115]), .Q (new_AGEMA_signal_13850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6029 ( .C (clk), .D (key_s1[115]), .Q (new_AGEMA_signal_13854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6033 ( .C (clk), .D (key_s2[115]), .Q (new_AGEMA_signal_13858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6037 ( .C (clk), .D (key_s3[115]), .Q (new_AGEMA_signal_13862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6041 ( .C (clk), .D (key_s0[116]), .Q (new_AGEMA_signal_13866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6045 ( .C (clk), .D (key_s1[116]), .Q (new_AGEMA_signal_13870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6049 ( .C (clk), .D (key_s2[116]), .Q (new_AGEMA_signal_13874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6053 ( .C (clk), .D (key_s3[116]), .Q (new_AGEMA_signal_13878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6057 ( .C (clk), .D (key_s0[117]), .Q (new_AGEMA_signal_13882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6061 ( .C (clk), .D (key_s1[117]), .Q (new_AGEMA_signal_13886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6065 ( .C (clk), .D (key_s2[117]), .Q (new_AGEMA_signal_13890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6069 ( .C (clk), .D (key_s3[117]), .Q (new_AGEMA_signal_13894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6073 ( .C (clk), .D (key_s0[118]), .Q (new_AGEMA_signal_13898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6077 ( .C (clk), .D (key_s1[118]), .Q (new_AGEMA_signal_13902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6081 ( .C (clk), .D (key_s2[118]), .Q (new_AGEMA_signal_13906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6085 ( .C (clk), .D (key_s3[118]), .Q (new_AGEMA_signal_13910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6089 ( .C (clk), .D (key_s0[119]), .Q (new_AGEMA_signal_13914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6093 ( .C (clk), .D (key_s1[119]), .Q (new_AGEMA_signal_13918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6097 ( .C (clk), .D (key_s2[119]), .Q (new_AGEMA_signal_13922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6101 ( .C (clk), .D (key_s3[119]), .Q (new_AGEMA_signal_13926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6105 ( .C (clk), .D (key_s0[120]), .Q (new_AGEMA_signal_13930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6109 ( .C (clk), .D (key_s1[120]), .Q (new_AGEMA_signal_13934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6113 ( .C (clk), .D (key_s2[120]), .Q (new_AGEMA_signal_13938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6117 ( .C (clk), .D (key_s3[120]), .Q (new_AGEMA_signal_13942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6121 ( .C (clk), .D (key_s0[121]), .Q (new_AGEMA_signal_13946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6125 ( .C (clk), .D (key_s1[121]), .Q (new_AGEMA_signal_13950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6129 ( .C (clk), .D (key_s2[121]), .Q (new_AGEMA_signal_13954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6133 ( .C (clk), .D (key_s3[121]), .Q (new_AGEMA_signal_13958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6137 ( .C (clk), .D (key_s0[122]), .Q (new_AGEMA_signal_13962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6141 ( .C (clk), .D (key_s1[122]), .Q (new_AGEMA_signal_13966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6145 ( .C (clk), .D (key_s2[122]), .Q (new_AGEMA_signal_13970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6149 ( .C (clk), .D (key_s3[122]), .Q (new_AGEMA_signal_13974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6153 ( .C (clk), .D (key_s0[123]), .Q (new_AGEMA_signal_13978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6157 ( .C (clk), .D (key_s1[123]), .Q (new_AGEMA_signal_13982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6161 ( .C (clk), .D (key_s2[123]), .Q (new_AGEMA_signal_13986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6165 ( .C (clk), .D (key_s3[123]), .Q (new_AGEMA_signal_13990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6169 ( .C (clk), .D (key_s0[124]), .Q (new_AGEMA_signal_13994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6173 ( .C (clk), .D (key_s1[124]), .Q (new_AGEMA_signal_13998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6177 ( .C (clk), .D (key_s2[124]), .Q (new_AGEMA_signal_14002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6181 ( .C (clk), .D (key_s3[124]), .Q (new_AGEMA_signal_14006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6185 ( .C (clk), .D (key_s0[125]), .Q (new_AGEMA_signal_14010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6189 ( .C (clk), .D (key_s1[125]), .Q (new_AGEMA_signal_14014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6193 ( .C (clk), .D (key_s2[125]), .Q (new_AGEMA_signal_14018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6197 ( .C (clk), .D (key_s3[125]), .Q (new_AGEMA_signal_14022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6201 ( .C (clk), .D (key_s0[126]), .Q (new_AGEMA_signal_14026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6205 ( .C (clk), .D (key_s1[126]), .Q (new_AGEMA_signal_14030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6209 ( .C (clk), .D (key_s2[126]), .Q (new_AGEMA_signal_14034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6213 ( .C (clk), .D (key_s3[126]), .Q (new_AGEMA_signal_14038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6217 ( .C (clk), .D (key_s0[127]), .Q (new_AGEMA_signal_14042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6221 ( .C (clk), .D (key_s1[127]), .Q (new_AGEMA_signal_14046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6225 ( .C (clk), .D (key_s2[127]), .Q (new_AGEMA_signal_14050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6229 ( .C (clk), .D (key_s3[127]), .Q (new_AGEMA_signal_14054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6233 ( .C (clk), .D (KSSubBytesInput[9]), .Q (new_AGEMA_signal_14058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6237 ( .C (clk), .D (new_AGEMA_signal_3484), .Q (new_AGEMA_signal_14062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6241 ( .C (clk), .D (new_AGEMA_signal_3485), .Q (new_AGEMA_signal_14066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6245 ( .C (clk), .D (new_AGEMA_signal_3486), .Q (new_AGEMA_signal_14070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6249 ( .C (clk), .D (KSSubBytesInput[8]), .Q (new_AGEMA_signal_14074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6253 ( .C (clk), .D (new_AGEMA_signal_3385), .Q (new_AGEMA_signal_14078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6257 ( .C (clk), .D (new_AGEMA_signal_3386), .Q (new_AGEMA_signal_14082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6261 ( .C (clk), .D (new_AGEMA_signal_3387), .Q (new_AGEMA_signal_14086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6265 ( .C (clk), .D (KSSubBytesInput[23]), .Q (new_AGEMA_signal_14090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6269 ( .C (clk), .D (new_AGEMA_signal_3286), .Q (new_AGEMA_signal_14094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6273 ( .C (clk), .D (new_AGEMA_signal_3287), .Q (new_AGEMA_signal_14098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6277 ( .C (clk), .D (new_AGEMA_signal_3288), .Q (new_AGEMA_signal_14102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6281 ( .C (clk), .D (KSSubBytesInput[22]), .Q (new_AGEMA_signal_14106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6285 ( .C (clk), .D (new_AGEMA_signal_3187), .Q (new_AGEMA_signal_14110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6289 ( .C (clk), .D (new_AGEMA_signal_3188), .Q (new_AGEMA_signal_14114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6293 ( .C (clk), .D (new_AGEMA_signal_3189), .Q (new_AGEMA_signal_14118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6297 ( .C (clk), .D (KSSubBytesInput[21]), .Q (new_AGEMA_signal_14122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6301 ( .C (clk), .D (new_AGEMA_signal_3088), .Q (new_AGEMA_signal_14126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6305 ( .C (clk), .D (new_AGEMA_signal_3089), .Q (new_AGEMA_signal_14130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6309 ( .C (clk), .D (new_AGEMA_signal_3090), .Q (new_AGEMA_signal_14134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6313 ( .C (clk), .D (KSSubBytesInput[20]), .Q (new_AGEMA_signal_14138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6317 ( .C (clk), .D (new_AGEMA_signal_2989), .Q (new_AGEMA_signal_14142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6321 ( .C (clk), .D (new_AGEMA_signal_2990), .Q (new_AGEMA_signal_14146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6325 ( .C (clk), .D (new_AGEMA_signal_2991), .Q (new_AGEMA_signal_14150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6329 ( .C (clk), .D (RoundKey[41]), .Q (new_AGEMA_signal_14154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6333 ( .C (clk), .D (new_AGEMA_signal_2908), .Q (new_AGEMA_signal_14158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6337 ( .C (clk), .D (new_AGEMA_signal_2909), .Q (new_AGEMA_signal_14162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6341 ( .C (clk), .D (new_AGEMA_signal_2910), .Q (new_AGEMA_signal_14166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6345 ( .C (clk), .D (RoundKey[73]), .Q (new_AGEMA_signal_14170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6349 ( .C (clk), .D (new_AGEMA_signal_3223), .Q (new_AGEMA_signal_14174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6353 ( .C (clk), .D (new_AGEMA_signal_3224), .Q (new_AGEMA_signal_14178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6357 ( .C (clk), .D (new_AGEMA_signal_3225), .Q (new_AGEMA_signal_14182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6361 ( .C (clk), .D (RoundKey[40]), .Q (new_AGEMA_signal_14186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6365 ( .C (clk), .D (new_AGEMA_signal_2899), .Q (new_AGEMA_signal_14190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6369 ( .C (clk), .D (new_AGEMA_signal_2900), .Q (new_AGEMA_signal_14194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6373 ( .C (clk), .D (new_AGEMA_signal_2901), .Q (new_AGEMA_signal_14198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6377 ( .C (clk), .D (RoundKey[72]), .Q (new_AGEMA_signal_14202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6381 ( .C (clk), .D (new_AGEMA_signal_3214), .Q (new_AGEMA_signal_14206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6385 ( .C (clk), .D (new_AGEMA_signal_3215), .Q (new_AGEMA_signal_14210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6389 ( .C (clk), .D (new_AGEMA_signal_3216), .Q (new_AGEMA_signal_14214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6393 ( .C (clk), .D (KSSubBytesInput[19]), .Q (new_AGEMA_signal_14218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6397 ( .C (clk), .D (new_AGEMA_signal_2890), .Q (new_AGEMA_signal_14222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6401 ( .C (clk), .D (new_AGEMA_signal_2891), .Q (new_AGEMA_signal_14226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6405 ( .C (clk), .D (new_AGEMA_signal_2892), .Q (new_AGEMA_signal_14230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6409 ( .C (clk), .D (RoundKey[39]), .Q (new_AGEMA_signal_14234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6413 ( .C (clk), .D (new_AGEMA_signal_2881), .Q (new_AGEMA_signal_14238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6417 ( .C (clk), .D (new_AGEMA_signal_2882), .Q (new_AGEMA_signal_14242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6421 ( .C (clk), .D (new_AGEMA_signal_2883), .Q (new_AGEMA_signal_14246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6425 ( .C (clk), .D (RoundKey[71]), .Q (new_AGEMA_signal_14250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6429 ( .C (clk), .D (new_AGEMA_signal_3205), .Q (new_AGEMA_signal_14254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6433 ( .C (clk), .D (new_AGEMA_signal_3206), .Q (new_AGEMA_signal_14258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6437 ( .C (clk), .D (new_AGEMA_signal_3207), .Q (new_AGEMA_signal_14262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6441 ( .C (clk), .D (RoundKey[38]), .Q (new_AGEMA_signal_14266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6445 ( .C (clk), .D (new_AGEMA_signal_2872), .Q (new_AGEMA_signal_14270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6449 ( .C (clk), .D (new_AGEMA_signal_2873), .Q (new_AGEMA_signal_14274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6453 ( .C (clk), .D (new_AGEMA_signal_2874), .Q (new_AGEMA_signal_14278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6457 ( .C (clk), .D (RoundKey[70]), .Q (new_AGEMA_signal_14282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6461 ( .C (clk), .D (new_AGEMA_signal_3196), .Q (new_AGEMA_signal_14286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6465 ( .C (clk), .D (new_AGEMA_signal_3197), .Q (new_AGEMA_signal_14290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6469 ( .C (clk), .D (new_AGEMA_signal_3198), .Q (new_AGEMA_signal_14294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6473 ( .C (clk), .D (RoundKey[37]), .Q (new_AGEMA_signal_14298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6477 ( .C (clk), .D (new_AGEMA_signal_2863), .Q (new_AGEMA_signal_14302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6481 ( .C (clk), .D (new_AGEMA_signal_2864), .Q (new_AGEMA_signal_14306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6485 ( .C (clk), .D (new_AGEMA_signal_2865), .Q (new_AGEMA_signal_14310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6489 ( .C (clk), .D (RoundKey[69]), .Q (new_AGEMA_signal_14314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6493 ( .C (clk), .D (new_AGEMA_signal_3178), .Q (new_AGEMA_signal_14318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6497 ( .C (clk), .D (new_AGEMA_signal_3179), .Q (new_AGEMA_signal_14322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6501 ( .C (clk), .D (new_AGEMA_signal_3180), .Q (new_AGEMA_signal_14326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6505 ( .C (clk), .D (RoundKey[36]), .Q (new_AGEMA_signal_14330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6509 ( .C (clk), .D (new_AGEMA_signal_2854), .Q (new_AGEMA_signal_14334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6513 ( .C (clk), .D (new_AGEMA_signal_2855), .Q (new_AGEMA_signal_14338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6517 ( .C (clk), .D (new_AGEMA_signal_2856), .Q (new_AGEMA_signal_14342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6521 ( .C (clk), .D (RoundKey[68]), .Q (new_AGEMA_signal_14346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6525 ( .C (clk), .D (new_AGEMA_signal_3169), .Q (new_AGEMA_signal_14350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6529 ( .C (clk), .D (new_AGEMA_signal_3170), .Q (new_AGEMA_signal_14354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6533 ( .C (clk), .D (new_AGEMA_signal_3171), .Q (new_AGEMA_signal_14358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6537 ( .C (clk), .D (RoundKey[35]), .Q (new_AGEMA_signal_14362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6541 ( .C (clk), .D (new_AGEMA_signal_2845), .Q (new_AGEMA_signal_14366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6545 ( .C (clk), .D (new_AGEMA_signal_2846), .Q (new_AGEMA_signal_14370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6549 ( .C (clk), .D (new_AGEMA_signal_2847), .Q (new_AGEMA_signal_14374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6553 ( .C (clk), .D (RoundKey[67]), .Q (new_AGEMA_signal_14378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6557 ( .C (clk), .D (new_AGEMA_signal_3160), .Q (new_AGEMA_signal_14382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6561 ( .C (clk), .D (new_AGEMA_signal_3161), .Q (new_AGEMA_signal_14386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6565 ( .C (clk), .D (new_AGEMA_signal_3162), .Q (new_AGEMA_signal_14390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6569 ( .C (clk), .D (RoundKey[99]), .Q (new_AGEMA_signal_14394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6573 ( .C (clk), .D (new_AGEMA_signal_3475), .Q (new_AGEMA_signal_14398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6577 ( .C (clk), .D (new_AGEMA_signal_3476), .Q (new_AGEMA_signal_14402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6581 ( .C (clk), .D (new_AGEMA_signal_3477), .Q (new_AGEMA_signal_14406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6585 ( .C (clk), .D (KSSubBytesInput[31]), .Q (new_AGEMA_signal_14410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6589 ( .C (clk), .D (new_AGEMA_signal_2809), .Q (new_AGEMA_signal_14414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6593 ( .C (clk), .D (new_AGEMA_signal_2810), .Q (new_AGEMA_signal_14418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6597 ( .C (clk), .D (new_AGEMA_signal_2811), .Q (new_AGEMA_signal_14422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6601 ( .C (clk), .D (RoundKey[63]), .Q (new_AGEMA_signal_14426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6605 ( .C (clk), .D (new_AGEMA_signal_3124), .Q (new_AGEMA_signal_14430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6609 ( .C (clk), .D (new_AGEMA_signal_3125), .Q (new_AGEMA_signal_14434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6613 ( .C (clk), .D (new_AGEMA_signal_3126), .Q (new_AGEMA_signal_14438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6617 ( .C (clk), .D (RoundKey[95]), .Q (new_AGEMA_signal_14442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6621 ( .C (clk), .D (new_AGEMA_signal_3439), .Q (new_AGEMA_signal_14446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6625 ( .C (clk), .D (new_AGEMA_signal_3440), .Q (new_AGEMA_signal_14450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6629 ( .C (clk), .D (new_AGEMA_signal_3441), .Q (new_AGEMA_signal_14454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6633 ( .C (clk), .D (KSSubBytesInput[30]), .Q (new_AGEMA_signal_14458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6637 ( .C (clk), .D (new_AGEMA_signal_2800), .Q (new_AGEMA_signal_14462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6641 ( .C (clk), .D (new_AGEMA_signal_2801), .Q (new_AGEMA_signal_14466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6645 ( .C (clk), .D (new_AGEMA_signal_2802), .Q (new_AGEMA_signal_14470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6649 ( .C (clk), .D (RoundKey[62]), .Q (new_AGEMA_signal_14474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6653 ( .C (clk), .D (new_AGEMA_signal_3115), .Q (new_AGEMA_signal_14478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6657 ( .C (clk), .D (new_AGEMA_signal_3116), .Q (new_AGEMA_signal_14482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6661 ( .C (clk), .D (new_AGEMA_signal_3117), .Q (new_AGEMA_signal_14486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6665 ( .C (clk), .D (RoundKey[94]), .Q (new_AGEMA_signal_14490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6669 ( .C (clk), .D (new_AGEMA_signal_3430), .Q (new_AGEMA_signal_14494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6673 ( .C (clk), .D (new_AGEMA_signal_3431), .Q (new_AGEMA_signal_14498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6677 ( .C (clk), .D (new_AGEMA_signal_3432), .Q (new_AGEMA_signal_14502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6681 ( .C (clk), .D (KSSubBytesInput[18]), .Q (new_AGEMA_signal_14506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6685 ( .C (clk), .D (new_AGEMA_signal_2791), .Q (new_AGEMA_signal_14510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6689 ( .C (clk), .D (new_AGEMA_signal_2792), .Q (new_AGEMA_signal_14514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6693 ( .C (clk), .D (new_AGEMA_signal_2793), .Q (new_AGEMA_signal_14518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6697 ( .C (clk), .D (RoundKey[34]), .Q (new_AGEMA_signal_14522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6701 ( .C (clk), .D (new_AGEMA_signal_2836), .Q (new_AGEMA_signal_14526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6705 ( .C (clk), .D (new_AGEMA_signal_2837), .Q (new_AGEMA_signal_14530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6709 ( .C (clk), .D (new_AGEMA_signal_2838), .Q (new_AGEMA_signal_14534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6713 ( .C (clk), .D (RoundKey[66]), .Q (new_AGEMA_signal_14538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6717 ( .C (clk), .D (new_AGEMA_signal_3151), .Q (new_AGEMA_signal_14542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6721 ( .C (clk), .D (new_AGEMA_signal_3152), .Q (new_AGEMA_signal_14546) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6725 ( .C (clk), .D (new_AGEMA_signal_3153), .Q (new_AGEMA_signal_14550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6729 ( .C (clk), .D (RoundKey[98]), .Q (new_AGEMA_signal_14554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6733 ( .C (clk), .D (new_AGEMA_signal_3466), .Q (new_AGEMA_signal_14558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6737 ( .C (clk), .D (new_AGEMA_signal_3467), .Q (new_AGEMA_signal_14562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6741 ( .C (clk), .D (new_AGEMA_signal_3468), .Q (new_AGEMA_signal_14566) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6745 ( .C (clk), .D (KSSubBytesInput[29]), .Q (new_AGEMA_signal_14570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6749 ( .C (clk), .D (new_AGEMA_signal_2782), .Q (new_AGEMA_signal_14574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6753 ( .C (clk), .D (new_AGEMA_signal_2783), .Q (new_AGEMA_signal_14578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6757 ( .C (clk), .D (new_AGEMA_signal_2784), .Q (new_AGEMA_signal_14582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6761 ( .C (clk), .D (RoundKey[61]), .Q (new_AGEMA_signal_14586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6765 ( .C (clk), .D (new_AGEMA_signal_3106), .Q (new_AGEMA_signal_14590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6769 ( .C (clk), .D (new_AGEMA_signal_3107), .Q (new_AGEMA_signal_14594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6773 ( .C (clk), .D (new_AGEMA_signal_3108), .Q (new_AGEMA_signal_14598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6777 ( .C (clk), .D (RoundKey[93]), .Q (new_AGEMA_signal_14602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6781 ( .C (clk), .D (new_AGEMA_signal_3421), .Q (new_AGEMA_signal_14606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6785 ( .C (clk), .D (new_AGEMA_signal_3422), .Q (new_AGEMA_signal_14610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6789 ( .C (clk), .D (new_AGEMA_signal_3423), .Q (new_AGEMA_signal_14614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6793 ( .C (clk), .D (KSSubBytesInput[28]), .Q (new_AGEMA_signal_14618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6797 ( .C (clk), .D (new_AGEMA_signal_2773), .Q (new_AGEMA_signal_14622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6801 ( .C (clk), .D (new_AGEMA_signal_2774), .Q (new_AGEMA_signal_14626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6805 ( .C (clk), .D (new_AGEMA_signal_2775), .Q (new_AGEMA_signal_14630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6809 ( .C (clk), .D (RoundKey[60]), .Q (new_AGEMA_signal_14634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6813 ( .C (clk), .D (new_AGEMA_signal_3097), .Q (new_AGEMA_signal_14638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6817 ( .C (clk), .D (new_AGEMA_signal_3098), .Q (new_AGEMA_signal_14642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6821 ( .C (clk), .D (new_AGEMA_signal_3099), .Q (new_AGEMA_signal_14646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6825 ( .C (clk), .D (RoundKey[92]), .Q (new_AGEMA_signal_14650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6829 ( .C (clk), .D (new_AGEMA_signal_3412), .Q (new_AGEMA_signal_14654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6833 ( .C (clk), .D (new_AGEMA_signal_3413), .Q (new_AGEMA_signal_14658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6837 ( .C (clk), .D (new_AGEMA_signal_3414), .Q (new_AGEMA_signal_14662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6841 ( .C (clk), .D (KSSubBytesInput[27]), .Q (new_AGEMA_signal_14666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6845 ( .C (clk), .D (new_AGEMA_signal_2764), .Q (new_AGEMA_signal_14670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6849 ( .C (clk), .D (new_AGEMA_signal_2765), .Q (new_AGEMA_signal_14674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6853 ( .C (clk), .D (new_AGEMA_signal_2766), .Q (new_AGEMA_signal_14678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6857 ( .C (clk), .D (RoundKey[59]), .Q (new_AGEMA_signal_14682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6861 ( .C (clk), .D (new_AGEMA_signal_3079), .Q (new_AGEMA_signal_14686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6865 ( .C (clk), .D (new_AGEMA_signal_3080), .Q (new_AGEMA_signal_14690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6869 ( .C (clk), .D (new_AGEMA_signal_3081), .Q (new_AGEMA_signal_14694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6873 ( .C (clk), .D (RoundKey[91]), .Q (new_AGEMA_signal_14698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6877 ( .C (clk), .D (new_AGEMA_signal_3403), .Q (new_AGEMA_signal_14702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6881 ( .C (clk), .D (new_AGEMA_signal_3404), .Q (new_AGEMA_signal_14706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6885 ( .C (clk), .D (new_AGEMA_signal_3405), .Q (new_AGEMA_signal_14710) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6889 ( .C (clk), .D (KSSubBytesInput[26]), .Q (new_AGEMA_signal_14714) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6893 ( .C (clk), .D (new_AGEMA_signal_2755), .Q (new_AGEMA_signal_14718) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6897 ( .C (clk), .D (new_AGEMA_signal_2756), .Q (new_AGEMA_signal_14722) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6901 ( .C (clk), .D (new_AGEMA_signal_2757), .Q (new_AGEMA_signal_14726) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6905 ( .C (clk), .D (RoundKey[58]), .Q (new_AGEMA_signal_14730) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6909 ( .C (clk), .D (new_AGEMA_signal_3070), .Q (new_AGEMA_signal_14734) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6913 ( .C (clk), .D (new_AGEMA_signal_3071), .Q (new_AGEMA_signal_14738) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6917 ( .C (clk), .D (new_AGEMA_signal_3072), .Q (new_AGEMA_signal_14742) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6921 ( .C (clk), .D (RoundKey[90]), .Q (new_AGEMA_signal_14746) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6925 ( .C (clk), .D (new_AGEMA_signal_3394), .Q (new_AGEMA_signal_14750) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6929 ( .C (clk), .D (new_AGEMA_signal_3395), .Q (new_AGEMA_signal_14754) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6933 ( .C (clk), .D (new_AGEMA_signal_3396), .Q (new_AGEMA_signal_14758) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6937 ( .C (clk), .D (KSSubBytesInput[25]), .Q (new_AGEMA_signal_14762) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6941 ( .C (clk), .D (new_AGEMA_signal_2746), .Q (new_AGEMA_signal_14766) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6945 ( .C (clk), .D (new_AGEMA_signal_2747), .Q (new_AGEMA_signal_14770) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6949 ( .C (clk), .D (new_AGEMA_signal_2748), .Q (new_AGEMA_signal_14774) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6953 ( .C (clk), .D (RoundKey[57]), .Q (new_AGEMA_signal_14778) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6957 ( .C (clk), .D (new_AGEMA_signal_3061), .Q (new_AGEMA_signal_14782) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6961 ( .C (clk), .D (new_AGEMA_signal_3062), .Q (new_AGEMA_signal_14786) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6965 ( .C (clk), .D (new_AGEMA_signal_3063), .Q (new_AGEMA_signal_14790) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6969 ( .C (clk), .D (RoundKey[89]), .Q (new_AGEMA_signal_14794) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6973 ( .C (clk), .D (new_AGEMA_signal_3376), .Q (new_AGEMA_signal_14798) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6977 ( .C (clk), .D (new_AGEMA_signal_3377), .Q (new_AGEMA_signal_14802) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6981 ( .C (clk), .D (new_AGEMA_signal_3378), .Q (new_AGEMA_signal_14806) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6985 ( .C (clk), .D (KSSubBytesInput[24]), .Q (new_AGEMA_signal_14810) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6989 ( .C (clk), .D (new_AGEMA_signal_2737), .Q (new_AGEMA_signal_14814) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6993 ( .C (clk), .D (new_AGEMA_signal_2738), .Q (new_AGEMA_signal_14818) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6997 ( .C (clk), .D (new_AGEMA_signal_2739), .Q (new_AGEMA_signal_14822) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7001 ( .C (clk), .D (RoundKey[56]), .Q (new_AGEMA_signal_14826) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7005 ( .C (clk), .D (new_AGEMA_signal_3052), .Q (new_AGEMA_signal_14830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7009 ( .C (clk), .D (new_AGEMA_signal_3053), .Q (new_AGEMA_signal_14834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7013 ( .C (clk), .D (new_AGEMA_signal_3054), .Q (new_AGEMA_signal_14838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7017 ( .C (clk), .D (RoundKey[88]), .Q (new_AGEMA_signal_14842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7021 ( .C (clk), .D (new_AGEMA_signal_3367), .Q (new_AGEMA_signal_14846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7025 ( .C (clk), .D (new_AGEMA_signal_3368), .Q (new_AGEMA_signal_14850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7029 ( .C (clk), .D (new_AGEMA_signal_3369), .Q (new_AGEMA_signal_14854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7033 ( .C (clk), .D (KSSubBytesInput[7]), .Q (new_AGEMA_signal_14858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7037 ( .C (clk), .D (new_AGEMA_signal_2728), .Q (new_AGEMA_signal_14862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7041 ( .C (clk), .D (new_AGEMA_signal_2729), .Q (new_AGEMA_signal_14866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7045 ( .C (clk), .D (new_AGEMA_signal_2730), .Q (new_AGEMA_signal_14870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7049 ( .C (clk), .D (RoundKey[55]), .Q (new_AGEMA_signal_14874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7053 ( .C (clk), .D (new_AGEMA_signal_3043), .Q (new_AGEMA_signal_14878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7057 ( .C (clk), .D (new_AGEMA_signal_3044), .Q (new_AGEMA_signal_14882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7061 ( .C (clk), .D (new_AGEMA_signal_3045), .Q (new_AGEMA_signal_14886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7065 ( .C (clk), .D (RoundKey[87]), .Q (new_AGEMA_signal_14890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7069 ( .C (clk), .D (new_AGEMA_signal_3358), .Q (new_AGEMA_signal_14894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7073 ( .C (clk), .D (new_AGEMA_signal_3359), .Q (new_AGEMA_signal_14898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7077 ( .C (clk), .D (new_AGEMA_signal_3360), .Q (new_AGEMA_signal_14902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7081 ( .C (clk), .D (KSSubBytesInput[6]), .Q (new_AGEMA_signal_14906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7085 ( .C (clk), .D (new_AGEMA_signal_2719), .Q (new_AGEMA_signal_14910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7089 ( .C (clk), .D (new_AGEMA_signal_2720), .Q (new_AGEMA_signal_14914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7093 ( .C (clk), .D (new_AGEMA_signal_2721), .Q (new_AGEMA_signal_14918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7097 ( .C (clk), .D (RoundKey[54]), .Q (new_AGEMA_signal_14922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7101 ( .C (clk), .D (new_AGEMA_signal_3034), .Q (new_AGEMA_signal_14926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7105 ( .C (clk), .D (new_AGEMA_signal_3035), .Q (new_AGEMA_signal_14930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7109 ( .C (clk), .D (new_AGEMA_signal_3036), .Q (new_AGEMA_signal_14934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7113 ( .C (clk), .D (RoundKey[86]), .Q (new_AGEMA_signal_14938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7117 ( .C (clk), .D (new_AGEMA_signal_3349), .Q (new_AGEMA_signal_14942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7121 ( .C (clk), .D (new_AGEMA_signal_3350), .Q (new_AGEMA_signal_14946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7125 ( .C (clk), .D (new_AGEMA_signal_3351), .Q (new_AGEMA_signal_14950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7129 ( .C (clk), .D (KSSubBytesInput[5]), .Q (new_AGEMA_signal_14954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7133 ( .C (clk), .D (new_AGEMA_signal_2710), .Q (new_AGEMA_signal_14958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7137 ( .C (clk), .D (new_AGEMA_signal_2711), .Q (new_AGEMA_signal_14962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7141 ( .C (clk), .D (new_AGEMA_signal_2712), .Q (new_AGEMA_signal_14966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7145 ( .C (clk), .D (RoundKey[53]), .Q (new_AGEMA_signal_14970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7149 ( .C (clk), .D (new_AGEMA_signal_3025), .Q (new_AGEMA_signal_14974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7153 ( .C (clk), .D (new_AGEMA_signal_3026), .Q (new_AGEMA_signal_14978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7157 ( .C (clk), .D (new_AGEMA_signal_3027), .Q (new_AGEMA_signal_14982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7161 ( .C (clk), .D (RoundKey[85]), .Q (new_AGEMA_signal_14986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7165 ( .C (clk), .D (new_AGEMA_signal_3340), .Q (new_AGEMA_signal_14990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7169 ( .C (clk), .D (new_AGEMA_signal_3341), .Q (new_AGEMA_signal_14994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7173 ( .C (clk), .D (new_AGEMA_signal_3342), .Q (new_AGEMA_signal_14998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7177 ( .C (clk), .D (KSSubBytesInput[4]), .Q (new_AGEMA_signal_15002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7181 ( .C (clk), .D (new_AGEMA_signal_2701), .Q (new_AGEMA_signal_15006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7185 ( .C (clk), .D (new_AGEMA_signal_2702), .Q (new_AGEMA_signal_15010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7189 ( .C (clk), .D (new_AGEMA_signal_2703), .Q (new_AGEMA_signal_15014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7193 ( .C (clk), .D (RoundKey[52]), .Q (new_AGEMA_signal_15018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7197 ( .C (clk), .D (new_AGEMA_signal_3016), .Q (new_AGEMA_signal_15022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7201 ( .C (clk), .D (new_AGEMA_signal_3017), .Q (new_AGEMA_signal_15026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7205 ( .C (clk), .D (new_AGEMA_signal_3018), .Q (new_AGEMA_signal_15030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7209 ( .C (clk), .D (RoundKey[84]), .Q (new_AGEMA_signal_15034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7213 ( .C (clk), .D (new_AGEMA_signal_3331), .Q (new_AGEMA_signal_15038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7217 ( .C (clk), .D (new_AGEMA_signal_3332), .Q (new_AGEMA_signal_15042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7221 ( .C (clk), .D (new_AGEMA_signal_3333), .Q (new_AGEMA_signal_15046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7225 ( .C (clk), .D (KSSubBytesInput[17]), .Q (new_AGEMA_signal_15050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7229 ( .C (clk), .D (new_AGEMA_signal_2692), .Q (new_AGEMA_signal_15054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7233 ( .C (clk), .D (new_AGEMA_signal_2693), .Q (new_AGEMA_signal_15058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7237 ( .C (clk), .D (new_AGEMA_signal_2694), .Q (new_AGEMA_signal_15062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7241 ( .C (clk), .D (RoundKey[33]), .Q (new_AGEMA_signal_15066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7245 ( .C (clk), .D (new_AGEMA_signal_2827), .Q (new_AGEMA_signal_15070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7249 ( .C (clk), .D (new_AGEMA_signal_2828), .Q (new_AGEMA_signal_15074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7253 ( .C (clk), .D (new_AGEMA_signal_2829), .Q (new_AGEMA_signal_15078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7257 ( .C (clk), .D (RoundKey[65]), .Q (new_AGEMA_signal_15082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7261 ( .C (clk), .D (new_AGEMA_signal_3142), .Q (new_AGEMA_signal_15086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7265 ( .C (clk), .D (new_AGEMA_signal_3143), .Q (new_AGEMA_signal_15090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7269 ( .C (clk), .D (new_AGEMA_signal_3144), .Q (new_AGEMA_signal_15094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7273 ( .C (clk), .D (RoundKey[97]), .Q (new_AGEMA_signal_15098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7277 ( .C (clk), .D (new_AGEMA_signal_3457), .Q (new_AGEMA_signal_15102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7281 ( .C (clk), .D (new_AGEMA_signal_3458), .Q (new_AGEMA_signal_15106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7285 ( .C (clk), .D (new_AGEMA_signal_3459), .Q (new_AGEMA_signal_15110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7289 ( .C (clk), .D (KSSubBytesInput[3]), .Q (new_AGEMA_signal_15114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7293 ( .C (clk), .D (new_AGEMA_signal_2683), .Q (new_AGEMA_signal_15118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7297 ( .C (clk), .D (new_AGEMA_signal_2684), .Q (new_AGEMA_signal_15122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7301 ( .C (clk), .D (new_AGEMA_signal_2685), .Q (new_AGEMA_signal_15126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7305 ( .C (clk), .D (RoundKey[51]), .Q (new_AGEMA_signal_15130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7309 ( .C (clk), .D (new_AGEMA_signal_3007), .Q (new_AGEMA_signal_15134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7313 ( .C (clk), .D (new_AGEMA_signal_3008), .Q (new_AGEMA_signal_15138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7317 ( .C (clk), .D (new_AGEMA_signal_3009), .Q (new_AGEMA_signal_15142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7321 ( .C (clk), .D (RoundKey[83]), .Q (new_AGEMA_signal_15146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7325 ( .C (clk), .D (new_AGEMA_signal_3322), .Q (new_AGEMA_signal_15150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7329 ( .C (clk), .D (new_AGEMA_signal_3323), .Q (new_AGEMA_signal_15154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7333 ( .C (clk), .D (new_AGEMA_signal_3324), .Q (new_AGEMA_signal_15158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7337 ( .C (clk), .D (KSSubBytesInput[2]), .Q (new_AGEMA_signal_15162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7341 ( .C (clk), .D (new_AGEMA_signal_2674), .Q (new_AGEMA_signal_15166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7345 ( .C (clk), .D (new_AGEMA_signal_2675), .Q (new_AGEMA_signal_15170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7349 ( .C (clk), .D (new_AGEMA_signal_2676), .Q (new_AGEMA_signal_15174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7353 ( .C (clk), .D (RoundKey[50]), .Q (new_AGEMA_signal_15178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7357 ( .C (clk), .D (new_AGEMA_signal_2998), .Q (new_AGEMA_signal_15182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7361 ( .C (clk), .D (new_AGEMA_signal_2999), .Q (new_AGEMA_signal_15186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7365 ( .C (clk), .D (new_AGEMA_signal_3000), .Q (new_AGEMA_signal_15190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7369 ( .C (clk), .D (RoundKey[82]), .Q (new_AGEMA_signal_15194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7373 ( .C (clk), .D (new_AGEMA_signal_3313), .Q (new_AGEMA_signal_15198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7377 ( .C (clk), .D (new_AGEMA_signal_3314), .Q (new_AGEMA_signal_15202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7381 ( .C (clk), .D (new_AGEMA_signal_3315), .Q (new_AGEMA_signal_15206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7385 ( .C (clk), .D (KSSubBytesInput[1]), .Q (new_AGEMA_signal_15210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7389 ( .C (clk), .D (new_AGEMA_signal_2665), .Q (new_AGEMA_signal_15214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7393 ( .C (clk), .D (new_AGEMA_signal_2666), .Q (new_AGEMA_signal_15218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7397 ( .C (clk), .D (new_AGEMA_signal_2667), .Q (new_AGEMA_signal_15222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7401 ( .C (clk), .D (RoundKey[49]), .Q (new_AGEMA_signal_15226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7405 ( .C (clk), .D (new_AGEMA_signal_2980), .Q (new_AGEMA_signal_15230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7409 ( .C (clk), .D (new_AGEMA_signal_2981), .Q (new_AGEMA_signal_15234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7413 ( .C (clk), .D (new_AGEMA_signal_2982), .Q (new_AGEMA_signal_15238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7417 ( .C (clk), .D (RoundKey[81]), .Q (new_AGEMA_signal_15242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7421 ( .C (clk), .D (new_AGEMA_signal_3304), .Q (new_AGEMA_signal_15246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7425 ( .C (clk), .D (new_AGEMA_signal_3305), .Q (new_AGEMA_signal_15250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7429 ( .C (clk), .D (new_AGEMA_signal_3306), .Q (new_AGEMA_signal_15254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7433 ( .C (clk), .D (KSSubBytesInput[0]), .Q (new_AGEMA_signal_15258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7437 ( .C (clk), .D (new_AGEMA_signal_2656), .Q (new_AGEMA_signal_15262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7441 ( .C (clk), .D (new_AGEMA_signal_2657), .Q (new_AGEMA_signal_15266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7445 ( .C (clk), .D (new_AGEMA_signal_2658), .Q (new_AGEMA_signal_15270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7449 ( .C (clk), .D (RoundKey[48]), .Q (new_AGEMA_signal_15274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7453 ( .C (clk), .D (new_AGEMA_signal_2971), .Q (new_AGEMA_signal_15278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7457 ( .C (clk), .D (new_AGEMA_signal_2972), .Q (new_AGEMA_signal_15282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7461 ( .C (clk), .D (new_AGEMA_signal_2973), .Q (new_AGEMA_signal_15286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7465 ( .C (clk), .D (RoundKey[80]), .Q (new_AGEMA_signal_15290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7469 ( .C (clk), .D (new_AGEMA_signal_3295), .Q (new_AGEMA_signal_15294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7473 ( .C (clk), .D (new_AGEMA_signal_3296), .Q (new_AGEMA_signal_15298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7477 ( .C (clk), .D (new_AGEMA_signal_3297), .Q (new_AGEMA_signal_15302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7481 ( .C (clk), .D (KSSubBytesInput[15]), .Q (new_AGEMA_signal_15306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7485 ( .C (clk), .D (new_AGEMA_signal_2647), .Q (new_AGEMA_signal_15310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7489 ( .C (clk), .D (new_AGEMA_signal_2648), .Q (new_AGEMA_signal_15314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7493 ( .C (clk), .D (new_AGEMA_signal_2649), .Q (new_AGEMA_signal_15318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7497 ( .C (clk), .D (RoundKey[47]), .Q (new_AGEMA_signal_15322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7501 ( .C (clk), .D (new_AGEMA_signal_2962), .Q (new_AGEMA_signal_15326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7505 ( .C (clk), .D (new_AGEMA_signal_2963), .Q (new_AGEMA_signal_15330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7509 ( .C (clk), .D (new_AGEMA_signal_2964), .Q (new_AGEMA_signal_15334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7513 ( .C (clk), .D (RoundKey[79]), .Q (new_AGEMA_signal_15338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7517 ( .C (clk), .D (new_AGEMA_signal_3277), .Q (new_AGEMA_signal_15342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7521 ( .C (clk), .D (new_AGEMA_signal_3278), .Q (new_AGEMA_signal_15346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7525 ( .C (clk), .D (new_AGEMA_signal_3279), .Q (new_AGEMA_signal_15350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7529 ( .C (clk), .D (KSSubBytesInput[14]), .Q (new_AGEMA_signal_15354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7533 ( .C (clk), .D (new_AGEMA_signal_2638), .Q (new_AGEMA_signal_15358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7537 ( .C (clk), .D (new_AGEMA_signal_2639), .Q (new_AGEMA_signal_15362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7541 ( .C (clk), .D (new_AGEMA_signal_2640), .Q (new_AGEMA_signal_15366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7545 ( .C (clk), .D (RoundKey[46]), .Q (new_AGEMA_signal_15370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7549 ( .C (clk), .D (new_AGEMA_signal_2953), .Q (new_AGEMA_signal_15374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7553 ( .C (clk), .D (new_AGEMA_signal_2954), .Q (new_AGEMA_signal_15378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7557 ( .C (clk), .D (new_AGEMA_signal_2955), .Q (new_AGEMA_signal_15382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7561 ( .C (clk), .D (RoundKey[78]), .Q (new_AGEMA_signal_15386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7565 ( .C (clk), .D (new_AGEMA_signal_3268), .Q (new_AGEMA_signal_15390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7569 ( .C (clk), .D (new_AGEMA_signal_3269), .Q (new_AGEMA_signal_15394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7573 ( .C (clk), .D (new_AGEMA_signal_3270), .Q (new_AGEMA_signal_15398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7577 ( .C (clk), .D (KSSubBytesInput[13]), .Q (new_AGEMA_signal_15402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7581 ( .C (clk), .D (new_AGEMA_signal_2629), .Q (new_AGEMA_signal_15406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7585 ( .C (clk), .D (new_AGEMA_signal_2630), .Q (new_AGEMA_signal_15410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7589 ( .C (clk), .D (new_AGEMA_signal_2631), .Q (new_AGEMA_signal_15414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7593 ( .C (clk), .D (RoundKey[45]), .Q (new_AGEMA_signal_15418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7597 ( .C (clk), .D (new_AGEMA_signal_2944), .Q (new_AGEMA_signal_15422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7601 ( .C (clk), .D (new_AGEMA_signal_2945), .Q (new_AGEMA_signal_15426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7605 ( .C (clk), .D (new_AGEMA_signal_2946), .Q (new_AGEMA_signal_15430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7609 ( .C (clk), .D (RoundKey[77]), .Q (new_AGEMA_signal_15434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7613 ( .C (clk), .D (new_AGEMA_signal_3259), .Q (new_AGEMA_signal_15438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7617 ( .C (clk), .D (new_AGEMA_signal_3260), .Q (new_AGEMA_signal_15442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7621 ( .C (clk), .D (new_AGEMA_signal_3261), .Q (new_AGEMA_signal_15446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7625 ( .C (clk), .D (KSSubBytesInput[12]), .Q (new_AGEMA_signal_15450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7629 ( .C (clk), .D (new_AGEMA_signal_2620), .Q (new_AGEMA_signal_15454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7633 ( .C (clk), .D (new_AGEMA_signal_2621), .Q (new_AGEMA_signal_15458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7637 ( .C (clk), .D (new_AGEMA_signal_2622), .Q (new_AGEMA_signal_15462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7641 ( .C (clk), .D (RoundKey[44]), .Q (new_AGEMA_signal_15466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7645 ( .C (clk), .D (new_AGEMA_signal_2935), .Q (new_AGEMA_signal_15470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7649 ( .C (clk), .D (new_AGEMA_signal_2936), .Q (new_AGEMA_signal_15474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7653 ( .C (clk), .D (new_AGEMA_signal_2937), .Q (new_AGEMA_signal_15478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7657 ( .C (clk), .D (RoundKey[76]), .Q (new_AGEMA_signal_15482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7661 ( .C (clk), .D (new_AGEMA_signal_3250), .Q (new_AGEMA_signal_15486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7665 ( .C (clk), .D (new_AGEMA_signal_3251), .Q (new_AGEMA_signal_15490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7669 ( .C (clk), .D (new_AGEMA_signal_3252), .Q (new_AGEMA_signal_15494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7673 ( .C (clk), .D (RoundKey[127]), .Q (new_AGEMA_signal_15498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7677 ( .C (clk), .D (new_AGEMA_signal_2611), .Q (new_AGEMA_signal_15502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7681 ( .C (clk), .D (new_AGEMA_signal_2612), .Q (new_AGEMA_signal_15506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7685 ( .C (clk), .D (new_AGEMA_signal_2613), .Q (new_AGEMA_signal_15510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7689 ( .C (clk), .D (RoundKey[126]), .Q (new_AGEMA_signal_15514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7693 ( .C (clk), .D (new_AGEMA_signal_2602), .Q (new_AGEMA_signal_15518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7697 ( .C (clk), .D (new_AGEMA_signal_2603), .Q (new_AGEMA_signal_15522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7701 ( .C (clk), .D (new_AGEMA_signal_2604), .Q (new_AGEMA_signal_15526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7705 ( .C (clk), .D (RoundKey[125]), .Q (new_AGEMA_signal_15530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7709 ( .C (clk), .D (new_AGEMA_signal_2593), .Q (new_AGEMA_signal_15534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7713 ( .C (clk), .D (new_AGEMA_signal_2594), .Q (new_AGEMA_signal_15538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7717 ( .C (clk), .D (new_AGEMA_signal_2595), .Q (new_AGEMA_signal_15542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7721 ( .C (clk), .D (RoundKey[124]), .Q (new_AGEMA_signal_15546) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7725 ( .C (clk), .D (new_AGEMA_signal_2584), .Q (new_AGEMA_signal_15550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7729 ( .C (clk), .D (new_AGEMA_signal_2585), .Q (new_AGEMA_signal_15554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7733 ( .C (clk), .D (new_AGEMA_signal_2586), .Q (new_AGEMA_signal_15558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7737 ( .C (clk), .D (RoundKey[123]), .Q (new_AGEMA_signal_15562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7741 ( .C (clk), .D (new_AGEMA_signal_2575), .Q (new_AGEMA_signal_15566) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7745 ( .C (clk), .D (new_AGEMA_signal_2576), .Q (new_AGEMA_signal_15570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7749 ( .C (clk), .D (new_AGEMA_signal_2577), .Q (new_AGEMA_signal_15574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7753 ( .C (clk), .D (RoundKey[122]), .Q (new_AGEMA_signal_15578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7757 ( .C (clk), .D (new_AGEMA_signal_2566), .Q (new_AGEMA_signal_15582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7761 ( .C (clk), .D (new_AGEMA_signal_2567), .Q (new_AGEMA_signal_15586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7765 ( .C (clk), .D (new_AGEMA_signal_2568), .Q (new_AGEMA_signal_15590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7769 ( .C (clk), .D (RoundKey[121]), .Q (new_AGEMA_signal_15594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7773 ( .C (clk), .D (new_AGEMA_signal_2557), .Q (new_AGEMA_signal_15598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7777 ( .C (clk), .D (new_AGEMA_signal_2558), .Q (new_AGEMA_signal_15602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7781 ( .C (clk), .D (new_AGEMA_signal_2559), .Q (new_AGEMA_signal_15606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7785 ( .C (clk), .D (RoundKey[120]), .Q (new_AGEMA_signal_15610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7789 ( .C (clk), .D (new_AGEMA_signal_2548), .Q (new_AGEMA_signal_15614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7793 ( .C (clk), .D (new_AGEMA_signal_2549), .Q (new_AGEMA_signal_15618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7797 ( .C (clk), .D (new_AGEMA_signal_2550), .Q (new_AGEMA_signal_15622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7801 ( .C (clk), .D (KSSubBytesInput[11]), .Q (new_AGEMA_signal_15626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7805 ( .C (clk), .D (new_AGEMA_signal_2539), .Q (new_AGEMA_signal_15630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7809 ( .C (clk), .D (new_AGEMA_signal_2540), .Q (new_AGEMA_signal_15634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7813 ( .C (clk), .D (new_AGEMA_signal_2541), .Q (new_AGEMA_signal_15638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7817 ( .C (clk), .D (RoundKey[43]), .Q (new_AGEMA_signal_15642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7821 ( .C (clk), .D (new_AGEMA_signal_2926), .Q (new_AGEMA_signal_15646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7825 ( .C (clk), .D (new_AGEMA_signal_2927), .Q (new_AGEMA_signal_15650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7829 ( .C (clk), .D (new_AGEMA_signal_2928), .Q (new_AGEMA_signal_15654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7833 ( .C (clk), .D (RoundKey[75]), .Q (new_AGEMA_signal_15658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7837 ( .C (clk), .D (new_AGEMA_signal_3241), .Q (new_AGEMA_signal_15662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7841 ( .C (clk), .D (new_AGEMA_signal_3242), .Q (new_AGEMA_signal_15666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7845 ( .C (clk), .D (new_AGEMA_signal_3243), .Q (new_AGEMA_signal_15670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7849 ( .C (clk), .D (RoundKey[119]), .Q (new_AGEMA_signal_15674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7853 ( .C (clk), .D (new_AGEMA_signal_2530), .Q (new_AGEMA_signal_15678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7857 ( .C (clk), .D (new_AGEMA_signal_2531), .Q (new_AGEMA_signal_15682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7861 ( .C (clk), .D (new_AGEMA_signal_2532), .Q (new_AGEMA_signal_15686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7865 ( .C (clk), .D (RoundKey[118]), .Q (new_AGEMA_signal_15690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7869 ( .C (clk), .D (new_AGEMA_signal_2521), .Q (new_AGEMA_signal_15694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7873 ( .C (clk), .D (new_AGEMA_signal_2522), .Q (new_AGEMA_signal_15698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7877 ( .C (clk), .D (new_AGEMA_signal_2523), .Q (new_AGEMA_signal_15702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7881 ( .C (clk), .D (RoundKey[117]), .Q (new_AGEMA_signal_15706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7885 ( .C (clk), .D (new_AGEMA_signal_2512), .Q (new_AGEMA_signal_15710) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7889 ( .C (clk), .D (new_AGEMA_signal_2513), .Q (new_AGEMA_signal_15714) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7893 ( .C (clk), .D (new_AGEMA_signal_2514), .Q (new_AGEMA_signal_15718) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7897 ( .C (clk), .D (RoundKey[116]), .Q (new_AGEMA_signal_15722) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7901 ( .C (clk), .D (new_AGEMA_signal_2503), .Q (new_AGEMA_signal_15726) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7905 ( .C (clk), .D (new_AGEMA_signal_2504), .Q (new_AGEMA_signal_15730) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7909 ( .C (clk), .D (new_AGEMA_signal_2505), .Q (new_AGEMA_signal_15734) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7913 ( .C (clk), .D (RoundKey[115]), .Q (new_AGEMA_signal_15738) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7917 ( .C (clk), .D (new_AGEMA_signal_2494), .Q (new_AGEMA_signal_15742) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7921 ( .C (clk), .D (new_AGEMA_signal_2495), .Q (new_AGEMA_signal_15746) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7925 ( .C (clk), .D (new_AGEMA_signal_2496), .Q (new_AGEMA_signal_15750) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7929 ( .C (clk), .D (RoundKey[114]), .Q (new_AGEMA_signal_15754) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7933 ( .C (clk), .D (new_AGEMA_signal_2485), .Q (new_AGEMA_signal_15758) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7937 ( .C (clk), .D (new_AGEMA_signal_2486), .Q (new_AGEMA_signal_15762) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7941 ( .C (clk), .D (new_AGEMA_signal_2487), .Q (new_AGEMA_signal_15766) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7945 ( .C (clk), .D (RoundKey[113]), .Q (new_AGEMA_signal_15770) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7949 ( .C (clk), .D (new_AGEMA_signal_2476), .Q (new_AGEMA_signal_15774) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7953 ( .C (clk), .D (new_AGEMA_signal_2477), .Q (new_AGEMA_signal_15778) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7957 ( .C (clk), .D (new_AGEMA_signal_2478), .Q (new_AGEMA_signal_15782) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7961 ( .C (clk), .D (RoundKey[112]), .Q (new_AGEMA_signal_15786) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7965 ( .C (clk), .D (new_AGEMA_signal_2467), .Q (new_AGEMA_signal_15790) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7969 ( .C (clk), .D (new_AGEMA_signal_2468), .Q (new_AGEMA_signal_15794) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7973 ( .C (clk), .D (new_AGEMA_signal_2469), .Q (new_AGEMA_signal_15798) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7977 ( .C (clk), .D (RoundKey[111]), .Q (new_AGEMA_signal_15802) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7981 ( .C (clk), .D (new_AGEMA_signal_2458), .Q (new_AGEMA_signal_15806) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7985 ( .C (clk), .D (new_AGEMA_signal_2459), .Q (new_AGEMA_signal_15810) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7989 ( .C (clk), .D (new_AGEMA_signal_2460), .Q (new_AGEMA_signal_15814) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7993 ( .C (clk), .D (RoundKey[110]), .Q (new_AGEMA_signal_15818) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7997 ( .C (clk), .D (new_AGEMA_signal_2449), .Q (new_AGEMA_signal_15822) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8001 ( .C (clk), .D (new_AGEMA_signal_2450), .Q (new_AGEMA_signal_15826) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8005 ( .C (clk), .D (new_AGEMA_signal_2451), .Q (new_AGEMA_signal_15830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8009 ( .C (clk), .D (KSSubBytesInput[10]), .Q (new_AGEMA_signal_15834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8013 ( .C (clk), .D (new_AGEMA_signal_2440), .Q (new_AGEMA_signal_15838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8017 ( .C (clk), .D (new_AGEMA_signal_2441), .Q (new_AGEMA_signal_15842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8021 ( .C (clk), .D (new_AGEMA_signal_2442), .Q (new_AGEMA_signal_15846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8025 ( .C (clk), .D (RoundKey[42]), .Q (new_AGEMA_signal_15850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8029 ( .C (clk), .D (new_AGEMA_signal_2917), .Q (new_AGEMA_signal_15854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8033 ( .C (clk), .D (new_AGEMA_signal_2918), .Q (new_AGEMA_signal_15858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8037 ( .C (clk), .D (new_AGEMA_signal_2919), .Q (new_AGEMA_signal_15862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8041 ( .C (clk), .D (RoundKey[74]), .Q (new_AGEMA_signal_15866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8045 ( .C (clk), .D (new_AGEMA_signal_3232), .Q (new_AGEMA_signal_15870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8049 ( .C (clk), .D (new_AGEMA_signal_3233), .Q (new_AGEMA_signal_15874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8053 ( .C (clk), .D (new_AGEMA_signal_3234), .Q (new_AGEMA_signal_15878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8057 ( .C (clk), .D (RoundKey[109]), .Q (new_AGEMA_signal_15882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8061 ( .C (clk), .D (new_AGEMA_signal_2431), .Q (new_AGEMA_signal_15886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8065 ( .C (clk), .D (new_AGEMA_signal_2432), .Q (new_AGEMA_signal_15890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8069 ( .C (clk), .D (new_AGEMA_signal_2433), .Q (new_AGEMA_signal_15894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8073 ( .C (clk), .D (RoundKey[108]), .Q (new_AGEMA_signal_15898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8077 ( .C (clk), .D (new_AGEMA_signal_2422), .Q (new_AGEMA_signal_15902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8081 ( .C (clk), .D (new_AGEMA_signal_2423), .Q (new_AGEMA_signal_15906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8085 ( .C (clk), .D (new_AGEMA_signal_2424), .Q (new_AGEMA_signal_15910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8089 ( .C (clk), .D (RoundKey[107]), .Q (new_AGEMA_signal_15914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8093 ( .C (clk), .D (new_AGEMA_signal_2413), .Q (new_AGEMA_signal_15918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8097 ( .C (clk), .D (new_AGEMA_signal_2414), .Q (new_AGEMA_signal_15922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8101 ( .C (clk), .D (new_AGEMA_signal_2415), .Q (new_AGEMA_signal_15926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8105 ( .C (clk), .D (RoundKey[106]), .Q (new_AGEMA_signal_15930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8109 ( .C (clk), .D (new_AGEMA_signal_2404), .Q (new_AGEMA_signal_15934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8113 ( .C (clk), .D (new_AGEMA_signal_2405), .Q (new_AGEMA_signal_15938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8117 ( .C (clk), .D (new_AGEMA_signal_2406), .Q (new_AGEMA_signal_15942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8121 ( .C (clk), .D (RoundKey[105]), .Q (new_AGEMA_signal_15946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8125 ( .C (clk), .D (new_AGEMA_signal_2395), .Q (new_AGEMA_signal_15950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8129 ( .C (clk), .D (new_AGEMA_signal_2396), .Q (new_AGEMA_signal_15954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8133 ( .C (clk), .D (new_AGEMA_signal_2397), .Q (new_AGEMA_signal_15958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8137 ( .C (clk), .D (RoundKey[104]), .Q (new_AGEMA_signal_15962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8141 ( .C (clk), .D (new_AGEMA_signal_2386), .Q (new_AGEMA_signal_15966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8145 ( .C (clk), .D (new_AGEMA_signal_2387), .Q (new_AGEMA_signal_15970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8149 ( .C (clk), .D (new_AGEMA_signal_2388), .Q (new_AGEMA_signal_15974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8153 ( .C (clk), .D (RoundKey[103]), .Q (new_AGEMA_signal_15978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8157 ( .C (clk), .D (new_AGEMA_signal_2377), .Q (new_AGEMA_signal_15982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8161 ( .C (clk), .D (new_AGEMA_signal_2378), .Q (new_AGEMA_signal_15986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8165 ( .C (clk), .D (new_AGEMA_signal_2379), .Q (new_AGEMA_signal_15990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8169 ( .C (clk), .D (RoundKey[102]), .Q (new_AGEMA_signal_15994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8173 ( .C (clk), .D (new_AGEMA_signal_2368), .Q (new_AGEMA_signal_15998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8177 ( .C (clk), .D (new_AGEMA_signal_2369), .Q (new_AGEMA_signal_16002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8181 ( .C (clk), .D (new_AGEMA_signal_2370), .Q (new_AGEMA_signal_16006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8185 ( .C (clk), .D (RoundKey[101]), .Q (new_AGEMA_signal_16010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8189 ( .C (clk), .D (new_AGEMA_signal_2359), .Q (new_AGEMA_signal_16014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8193 ( .C (clk), .D (new_AGEMA_signal_2360), .Q (new_AGEMA_signal_16018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8197 ( .C (clk), .D (new_AGEMA_signal_2361), .Q (new_AGEMA_signal_16022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8201 ( .C (clk), .D (RoundKey[100]), .Q (new_AGEMA_signal_16026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8205 ( .C (clk), .D (new_AGEMA_signal_2350), .Q (new_AGEMA_signal_16030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8209 ( .C (clk), .D (new_AGEMA_signal_2351), .Q (new_AGEMA_signal_16034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8213 ( .C (clk), .D (new_AGEMA_signal_2352), .Q (new_AGEMA_signal_16038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8217 ( .C (clk), .D (KSSubBytesInput[16]), .Q (new_AGEMA_signal_16042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8221 ( .C (clk), .D (new_AGEMA_signal_2341), .Q (new_AGEMA_signal_16046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8225 ( .C (clk), .D (new_AGEMA_signal_2342), .Q (new_AGEMA_signal_16050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8229 ( .C (clk), .D (new_AGEMA_signal_2343), .Q (new_AGEMA_signal_16054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8233 ( .C (clk), .D (RoundKey[32]), .Q (new_AGEMA_signal_16058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8237 ( .C (clk), .D (new_AGEMA_signal_2818), .Q (new_AGEMA_signal_16062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8241 ( .C (clk), .D (new_AGEMA_signal_2819), .Q (new_AGEMA_signal_16066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8245 ( .C (clk), .D (new_AGEMA_signal_2820), .Q (new_AGEMA_signal_16070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8249 ( .C (clk), .D (RoundKey[64]), .Q (new_AGEMA_signal_16074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8253 ( .C (clk), .D (new_AGEMA_signal_3133), .Q (new_AGEMA_signal_16078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8257 ( .C (clk), .D (new_AGEMA_signal_3134), .Q (new_AGEMA_signal_16082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8261 ( .C (clk), .D (new_AGEMA_signal_3135), .Q (new_AGEMA_signal_16086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8265 ( .C (clk), .D (RoundKey[96]), .Q (new_AGEMA_signal_16090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8269 ( .C (clk), .D (new_AGEMA_signal_3448), .Q (new_AGEMA_signal_16094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8273 ( .C (clk), .D (new_AGEMA_signal_3449), .Q (new_AGEMA_signal_16098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8277 ( .C (clk), .D (new_AGEMA_signal_3450), .Q (new_AGEMA_signal_16102) ) ;
    buf_clk new_AGEMA_reg_buffer_8281 ( .C (clk), .D (Rcon[7]), .Q (new_AGEMA_signal_16106) ) ;
    buf_clk new_AGEMA_reg_buffer_8285 ( .C (clk), .D (Rcon[6]), .Q (new_AGEMA_signal_16110) ) ;
    buf_clk new_AGEMA_reg_buffer_8289 ( .C (clk), .D (Rcon[5]), .Q (new_AGEMA_signal_16114) ) ;
    buf_clk new_AGEMA_reg_buffer_8293 ( .C (clk), .D (Rcon[4]), .Q (new_AGEMA_signal_16118) ) ;
    buf_clk new_AGEMA_reg_buffer_8297 ( .C (clk), .D (Rcon[3]), .Q (new_AGEMA_signal_16122) ) ;
    buf_clk new_AGEMA_reg_buffer_8301 ( .C (clk), .D (Rcon[2]), .Q (new_AGEMA_signal_16126) ) ;
    buf_clk new_AGEMA_reg_buffer_8305 ( .C (clk), .D (Rcon[1]), .Q (new_AGEMA_signal_16130) ) ;
    buf_clk new_AGEMA_reg_buffer_8309 ( .C (clk), .D (Rcon[0]), .Q (new_AGEMA_signal_16134) ) ;
    buf_clk new_AGEMA_reg_buffer_8313 ( .C (clk), .D (MuxKeyExpansion_n15), .Q (new_AGEMA_signal_16138) ) ;
    buf_clk new_AGEMA_reg_buffer_8317 ( .C (clk), .D (MuxKeyExpansion_n16), .Q (new_AGEMA_signal_16142) ) ;
    buf_clk new_AGEMA_reg_buffer_8321 ( .C (clk), .D (MuxKeyExpansion_n17), .Q (new_AGEMA_signal_16146) ) ;
    buf_clk new_AGEMA_reg_buffer_8325 ( .C (clk), .D (MuxKeyExpansion_n18), .Q (new_AGEMA_signal_16150) ) ;
    buf_clk new_AGEMA_reg_buffer_8329 ( .C (clk), .D (MuxKeyExpansion_n19), .Q (new_AGEMA_signal_16154) ) ;
    buf_clk new_AGEMA_reg_buffer_8333 ( .C (clk), .D (MuxKeyExpansion_n20), .Q (new_AGEMA_signal_16158) ) ;
    buf_clk new_AGEMA_reg_buffer_8337 ( .C (clk), .D (MuxKeyExpansion_n14), .Q (new_AGEMA_signal_16162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8341 ( .C (clk), .D (RoundReg_Inst_ff_SDE_32_next_state), .Q (new_AGEMA_signal_16166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8345 ( .C (clk), .D (new_AGEMA_signal_3877), .Q (new_AGEMA_signal_16170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8349 ( .C (clk), .D (new_AGEMA_signal_3878), .Q (new_AGEMA_signal_16174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8353 ( .C (clk), .D (new_AGEMA_signal_3879), .Q (new_AGEMA_signal_16178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8357 ( .C (clk), .D (RoundReg_Inst_ff_SDE_33_next_state), .Q (new_AGEMA_signal_16182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8361 ( .C (clk), .D (new_AGEMA_signal_3883), .Q (new_AGEMA_signal_16186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8365 ( .C (clk), .D (new_AGEMA_signal_3884), .Q (new_AGEMA_signal_16190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8369 ( .C (clk), .D (new_AGEMA_signal_3885), .Q (new_AGEMA_signal_16194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8373 ( .C (clk), .D (RoundReg_Inst_ff_SDE_34_next_state), .Q (new_AGEMA_signal_16198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8377 ( .C (clk), .D (new_AGEMA_signal_3889), .Q (new_AGEMA_signal_16202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8381 ( .C (clk), .D (new_AGEMA_signal_3890), .Q (new_AGEMA_signal_16206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8385 ( .C (clk), .D (new_AGEMA_signal_3891), .Q (new_AGEMA_signal_16210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8389 ( .C (clk), .D (RoundReg_Inst_ff_SDE_35_next_state), .Q (new_AGEMA_signal_16214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8393 ( .C (clk), .D (new_AGEMA_signal_3895), .Q (new_AGEMA_signal_16218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8397 ( .C (clk), .D (new_AGEMA_signal_3896), .Q (new_AGEMA_signal_16222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8401 ( .C (clk), .D (new_AGEMA_signal_3897), .Q (new_AGEMA_signal_16226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8405 ( .C (clk), .D (RoundReg_Inst_ff_SDE_36_next_state), .Q (new_AGEMA_signal_16230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8409 ( .C (clk), .D (new_AGEMA_signal_3901), .Q (new_AGEMA_signal_16234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8413 ( .C (clk), .D (new_AGEMA_signal_3902), .Q (new_AGEMA_signal_16238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8417 ( .C (clk), .D (new_AGEMA_signal_3903), .Q (new_AGEMA_signal_16242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8421 ( .C (clk), .D (RoundReg_Inst_ff_SDE_37_next_state), .Q (new_AGEMA_signal_16246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8425 ( .C (clk), .D (new_AGEMA_signal_3907), .Q (new_AGEMA_signal_16250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8429 ( .C (clk), .D (new_AGEMA_signal_3908), .Q (new_AGEMA_signal_16254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8433 ( .C (clk), .D (new_AGEMA_signal_3909), .Q (new_AGEMA_signal_16258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8437 ( .C (clk), .D (RoundReg_Inst_ff_SDE_38_next_state), .Q (new_AGEMA_signal_16262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8441 ( .C (clk), .D (new_AGEMA_signal_3913), .Q (new_AGEMA_signal_16266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8445 ( .C (clk), .D (new_AGEMA_signal_3914), .Q (new_AGEMA_signal_16270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8449 ( .C (clk), .D (new_AGEMA_signal_3915), .Q (new_AGEMA_signal_16274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8453 ( .C (clk), .D (RoundReg_Inst_ff_SDE_39_next_state), .Q (new_AGEMA_signal_16278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8457 ( .C (clk), .D (new_AGEMA_signal_3919), .Q (new_AGEMA_signal_16282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8461 ( .C (clk), .D (new_AGEMA_signal_3920), .Q (new_AGEMA_signal_16286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8465 ( .C (clk), .D (new_AGEMA_signal_3921), .Q (new_AGEMA_signal_16290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8469 ( .C (clk), .D (RoundReg_Inst_ff_SDE_40_next_state), .Q (new_AGEMA_signal_16294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8473 ( .C (clk), .D (new_AGEMA_signal_3925), .Q (new_AGEMA_signal_16298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8477 ( .C (clk), .D (new_AGEMA_signal_3926), .Q (new_AGEMA_signal_16302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8481 ( .C (clk), .D (new_AGEMA_signal_3927), .Q (new_AGEMA_signal_16306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8485 ( .C (clk), .D (RoundReg_Inst_ff_SDE_41_next_state), .Q (new_AGEMA_signal_16310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8489 ( .C (clk), .D (new_AGEMA_signal_3931), .Q (new_AGEMA_signal_16314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8493 ( .C (clk), .D (new_AGEMA_signal_3932), .Q (new_AGEMA_signal_16318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8497 ( .C (clk), .D (new_AGEMA_signal_3933), .Q (new_AGEMA_signal_16322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8501 ( .C (clk), .D (RoundReg_Inst_ff_SDE_42_next_state), .Q (new_AGEMA_signal_16326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8505 ( .C (clk), .D (new_AGEMA_signal_3937), .Q (new_AGEMA_signal_16330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8509 ( .C (clk), .D (new_AGEMA_signal_3938), .Q (new_AGEMA_signal_16334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8513 ( .C (clk), .D (new_AGEMA_signal_3939), .Q (new_AGEMA_signal_16338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8517 ( .C (clk), .D (RoundReg_Inst_ff_SDE_43_next_state), .Q (new_AGEMA_signal_16342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8521 ( .C (clk), .D (new_AGEMA_signal_3943), .Q (new_AGEMA_signal_16346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8525 ( .C (clk), .D (new_AGEMA_signal_3944), .Q (new_AGEMA_signal_16350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8529 ( .C (clk), .D (new_AGEMA_signal_3945), .Q (new_AGEMA_signal_16354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8533 ( .C (clk), .D (RoundReg_Inst_ff_SDE_44_next_state), .Q (new_AGEMA_signal_16358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8537 ( .C (clk), .D (new_AGEMA_signal_3949), .Q (new_AGEMA_signal_16362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8541 ( .C (clk), .D (new_AGEMA_signal_3950), .Q (new_AGEMA_signal_16366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8545 ( .C (clk), .D (new_AGEMA_signal_3951), .Q (new_AGEMA_signal_16370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8549 ( .C (clk), .D (RoundReg_Inst_ff_SDE_45_next_state), .Q (new_AGEMA_signal_16374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8553 ( .C (clk), .D (new_AGEMA_signal_3955), .Q (new_AGEMA_signal_16378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8557 ( .C (clk), .D (new_AGEMA_signal_3956), .Q (new_AGEMA_signal_16382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8561 ( .C (clk), .D (new_AGEMA_signal_3957), .Q (new_AGEMA_signal_16386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8565 ( .C (clk), .D (RoundReg_Inst_ff_SDE_46_next_state), .Q (new_AGEMA_signal_16390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8569 ( .C (clk), .D (new_AGEMA_signal_3961), .Q (new_AGEMA_signal_16394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8573 ( .C (clk), .D (new_AGEMA_signal_3962), .Q (new_AGEMA_signal_16398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8577 ( .C (clk), .D (new_AGEMA_signal_3963), .Q (new_AGEMA_signal_16402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8581 ( .C (clk), .D (RoundReg_Inst_ff_SDE_47_next_state), .Q (new_AGEMA_signal_16406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8585 ( .C (clk), .D (new_AGEMA_signal_3967), .Q (new_AGEMA_signal_16410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8589 ( .C (clk), .D (new_AGEMA_signal_3968), .Q (new_AGEMA_signal_16414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8593 ( .C (clk), .D (new_AGEMA_signal_3969), .Q (new_AGEMA_signal_16418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8597 ( .C (clk), .D (RoundReg_Inst_ff_SDE_48_next_state), .Q (new_AGEMA_signal_16422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8601 ( .C (clk), .D (new_AGEMA_signal_3973), .Q (new_AGEMA_signal_16426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8605 ( .C (clk), .D (new_AGEMA_signal_3974), .Q (new_AGEMA_signal_16430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8609 ( .C (clk), .D (new_AGEMA_signal_3975), .Q (new_AGEMA_signal_16434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8613 ( .C (clk), .D (RoundReg_Inst_ff_SDE_49_next_state), .Q (new_AGEMA_signal_16438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8617 ( .C (clk), .D (new_AGEMA_signal_3979), .Q (new_AGEMA_signal_16442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8621 ( .C (clk), .D (new_AGEMA_signal_3980), .Q (new_AGEMA_signal_16446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8625 ( .C (clk), .D (new_AGEMA_signal_3981), .Q (new_AGEMA_signal_16450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8629 ( .C (clk), .D (RoundReg_Inst_ff_SDE_50_next_state), .Q (new_AGEMA_signal_16454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8633 ( .C (clk), .D (new_AGEMA_signal_3985), .Q (new_AGEMA_signal_16458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8637 ( .C (clk), .D (new_AGEMA_signal_3986), .Q (new_AGEMA_signal_16462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8641 ( .C (clk), .D (new_AGEMA_signal_3987), .Q (new_AGEMA_signal_16466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8645 ( .C (clk), .D (RoundReg_Inst_ff_SDE_51_next_state), .Q (new_AGEMA_signal_16470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8649 ( .C (clk), .D (new_AGEMA_signal_3991), .Q (new_AGEMA_signal_16474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8653 ( .C (clk), .D (new_AGEMA_signal_3992), .Q (new_AGEMA_signal_16478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8657 ( .C (clk), .D (new_AGEMA_signal_3993), .Q (new_AGEMA_signal_16482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8661 ( .C (clk), .D (RoundReg_Inst_ff_SDE_52_next_state), .Q (new_AGEMA_signal_16486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8665 ( .C (clk), .D (new_AGEMA_signal_3997), .Q (new_AGEMA_signal_16490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8669 ( .C (clk), .D (new_AGEMA_signal_3998), .Q (new_AGEMA_signal_16494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8673 ( .C (clk), .D (new_AGEMA_signal_3999), .Q (new_AGEMA_signal_16498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8677 ( .C (clk), .D (RoundReg_Inst_ff_SDE_53_next_state), .Q (new_AGEMA_signal_16502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8681 ( .C (clk), .D (new_AGEMA_signal_4003), .Q (new_AGEMA_signal_16506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8685 ( .C (clk), .D (new_AGEMA_signal_4004), .Q (new_AGEMA_signal_16510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8689 ( .C (clk), .D (new_AGEMA_signal_4005), .Q (new_AGEMA_signal_16514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8693 ( .C (clk), .D (RoundReg_Inst_ff_SDE_54_next_state), .Q (new_AGEMA_signal_16518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8697 ( .C (clk), .D (new_AGEMA_signal_4009), .Q (new_AGEMA_signal_16522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8701 ( .C (clk), .D (new_AGEMA_signal_4010), .Q (new_AGEMA_signal_16526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8705 ( .C (clk), .D (new_AGEMA_signal_4011), .Q (new_AGEMA_signal_16530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8709 ( .C (clk), .D (RoundReg_Inst_ff_SDE_55_next_state), .Q (new_AGEMA_signal_16534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8713 ( .C (clk), .D (new_AGEMA_signal_4015), .Q (new_AGEMA_signal_16538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8717 ( .C (clk), .D (new_AGEMA_signal_4016), .Q (new_AGEMA_signal_16542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8721 ( .C (clk), .D (new_AGEMA_signal_4017), .Q (new_AGEMA_signal_16546) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8725 ( .C (clk), .D (RoundReg_Inst_ff_SDE_56_next_state), .Q (new_AGEMA_signal_16550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8729 ( .C (clk), .D (new_AGEMA_signal_4021), .Q (new_AGEMA_signal_16554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8733 ( .C (clk), .D (new_AGEMA_signal_4022), .Q (new_AGEMA_signal_16558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8737 ( .C (clk), .D (new_AGEMA_signal_4023), .Q (new_AGEMA_signal_16562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8741 ( .C (clk), .D (RoundReg_Inst_ff_SDE_57_next_state), .Q (new_AGEMA_signal_16566) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8745 ( .C (clk), .D (new_AGEMA_signal_4027), .Q (new_AGEMA_signal_16570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8749 ( .C (clk), .D (new_AGEMA_signal_4028), .Q (new_AGEMA_signal_16574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8753 ( .C (clk), .D (new_AGEMA_signal_4029), .Q (new_AGEMA_signal_16578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8757 ( .C (clk), .D (RoundReg_Inst_ff_SDE_58_next_state), .Q (new_AGEMA_signal_16582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8761 ( .C (clk), .D (new_AGEMA_signal_4033), .Q (new_AGEMA_signal_16586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8765 ( .C (clk), .D (new_AGEMA_signal_4034), .Q (new_AGEMA_signal_16590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8769 ( .C (clk), .D (new_AGEMA_signal_4035), .Q (new_AGEMA_signal_16594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8773 ( .C (clk), .D (RoundReg_Inst_ff_SDE_59_next_state), .Q (new_AGEMA_signal_16598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8777 ( .C (clk), .D (new_AGEMA_signal_4039), .Q (new_AGEMA_signal_16602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8781 ( .C (clk), .D (new_AGEMA_signal_4040), .Q (new_AGEMA_signal_16606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8785 ( .C (clk), .D (new_AGEMA_signal_4041), .Q (new_AGEMA_signal_16610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8789 ( .C (clk), .D (RoundReg_Inst_ff_SDE_60_next_state), .Q (new_AGEMA_signal_16614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8793 ( .C (clk), .D (new_AGEMA_signal_4045), .Q (new_AGEMA_signal_16618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8797 ( .C (clk), .D (new_AGEMA_signal_4046), .Q (new_AGEMA_signal_16622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8801 ( .C (clk), .D (new_AGEMA_signal_4047), .Q (new_AGEMA_signal_16626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8805 ( .C (clk), .D (RoundReg_Inst_ff_SDE_61_next_state), .Q (new_AGEMA_signal_16630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8809 ( .C (clk), .D (new_AGEMA_signal_4051), .Q (new_AGEMA_signal_16634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8813 ( .C (clk), .D (new_AGEMA_signal_4052), .Q (new_AGEMA_signal_16638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8817 ( .C (clk), .D (new_AGEMA_signal_4053), .Q (new_AGEMA_signal_16642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8821 ( .C (clk), .D (RoundReg_Inst_ff_SDE_62_next_state), .Q (new_AGEMA_signal_16646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8825 ( .C (clk), .D (new_AGEMA_signal_4057), .Q (new_AGEMA_signal_16650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8829 ( .C (clk), .D (new_AGEMA_signal_4058), .Q (new_AGEMA_signal_16654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8833 ( .C (clk), .D (new_AGEMA_signal_4059), .Q (new_AGEMA_signal_16658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8837 ( .C (clk), .D (RoundReg_Inst_ff_SDE_63_next_state), .Q (new_AGEMA_signal_16662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8841 ( .C (clk), .D (new_AGEMA_signal_4063), .Q (new_AGEMA_signal_16666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8845 ( .C (clk), .D (new_AGEMA_signal_4064), .Q (new_AGEMA_signal_16670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8849 ( .C (clk), .D (new_AGEMA_signal_4065), .Q (new_AGEMA_signal_16674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8853 ( .C (clk), .D (RoundReg_Inst_ff_SDE_64_next_state), .Q (new_AGEMA_signal_16678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8857 ( .C (clk), .D (new_AGEMA_signal_4069), .Q (new_AGEMA_signal_16682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8861 ( .C (clk), .D (new_AGEMA_signal_4070), .Q (new_AGEMA_signal_16686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8865 ( .C (clk), .D (new_AGEMA_signal_4071), .Q (new_AGEMA_signal_16690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8869 ( .C (clk), .D (RoundReg_Inst_ff_SDE_65_next_state), .Q (new_AGEMA_signal_16694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8873 ( .C (clk), .D (new_AGEMA_signal_4075), .Q (new_AGEMA_signal_16698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8877 ( .C (clk), .D (new_AGEMA_signal_4076), .Q (new_AGEMA_signal_16702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8881 ( .C (clk), .D (new_AGEMA_signal_4077), .Q (new_AGEMA_signal_16706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8885 ( .C (clk), .D (RoundReg_Inst_ff_SDE_66_next_state), .Q (new_AGEMA_signal_16710) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8889 ( .C (clk), .D (new_AGEMA_signal_4081), .Q (new_AGEMA_signal_16714) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8893 ( .C (clk), .D (new_AGEMA_signal_4082), .Q (new_AGEMA_signal_16718) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8897 ( .C (clk), .D (new_AGEMA_signal_4083), .Q (new_AGEMA_signal_16722) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8901 ( .C (clk), .D (RoundReg_Inst_ff_SDE_67_next_state), .Q (new_AGEMA_signal_16726) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8905 ( .C (clk), .D (new_AGEMA_signal_4087), .Q (new_AGEMA_signal_16730) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8909 ( .C (clk), .D (new_AGEMA_signal_4088), .Q (new_AGEMA_signal_16734) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8913 ( .C (clk), .D (new_AGEMA_signal_4089), .Q (new_AGEMA_signal_16738) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8917 ( .C (clk), .D (RoundReg_Inst_ff_SDE_68_next_state), .Q (new_AGEMA_signal_16742) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8921 ( .C (clk), .D (new_AGEMA_signal_4093), .Q (new_AGEMA_signal_16746) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8925 ( .C (clk), .D (new_AGEMA_signal_4094), .Q (new_AGEMA_signal_16750) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8929 ( .C (clk), .D (new_AGEMA_signal_4095), .Q (new_AGEMA_signal_16754) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8933 ( .C (clk), .D (RoundReg_Inst_ff_SDE_69_next_state), .Q (new_AGEMA_signal_16758) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8937 ( .C (clk), .D (new_AGEMA_signal_4099), .Q (new_AGEMA_signal_16762) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8941 ( .C (clk), .D (new_AGEMA_signal_4100), .Q (new_AGEMA_signal_16766) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8945 ( .C (clk), .D (new_AGEMA_signal_4101), .Q (new_AGEMA_signal_16770) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8949 ( .C (clk), .D (RoundReg_Inst_ff_SDE_70_next_state), .Q (new_AGEMA_signal_16774) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8953 ( .C (clk), .D (new_AGEMA_signal_4105), .Q (new_AGEMA_signal_16778) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8957 ( .C (clk), .D (new_AGEMA_signal_4106), .Q (new_AGEMA_signal_16782) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8961 ( .C (clk), .D (new_AGEMA_signal_4107), .Q (new_AGEMA_signal_16786) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8965 ( .C (clk), .D (RoundReg_Inst_ff_SDE_71_next_state), .Q (new_AGEMA_signal_16790) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8969 ( .C (clk), .D (new_AGEMA_signal_4111), .Q (new_AGEMA_signal_16794) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8973 ( .C (clk), .D (new_AGEMA_signal_4112), .Q (new_AGEMA_signal_16798) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8977 ( .C (clk), .D (new_AGEMA_signal_4113), .Q (new_AGEMA_signal_16802) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8981 ( .C (clk), .D (RoundReg_Inst_ff_SDE_72_next_state), .Q (new_AGEMA_signal_16806) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8985 ( .C (clk), .D (new_AGEMA_signal_4117), .Q (new_AGEMA_signal_16810) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8989 ( .C (clk), .D (new_AGEMA_signal_4118), .Q (new_AGEMA_signal_16814) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8993 ( .C (clk), .D (new_AGEMA_signal_4119), .Q (new_AGEMA_signal_16818) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8997 ( .C (clk), .D (RoundReg_Inst_ff_SDE_73_next_state), .Q (new_AGEMA_signal_16822) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9001 ( .C (clk), .D (new_AGEMA_signal_4123), .Q (new_AGEMA_signal_16826) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9005 ( .C (clk), .D (new_AGEMA_signal_4124), .Q (new_AGEMA_signal_16830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9009 ( .C (clk), .D (new_AGEMA_signal_4125), .Q (new_AGEMA_signal_16834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9013 ( .C (clk), .D (RoundReg_Inst_ff_SDE_74_next_state), .Q (new_AGEMA_signal_16838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9017 ( .C (clk), .D (new_AGEMA_signal_4129), .Q (new_AGEMA_signal_16842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9021 ( .C (clk), .D (new_AGEMA_signal_4130), .Q (new_AGEMA_signal_16846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9025 ( .C (clk), .D (new_AGEMA_signal_4131), .Q (new_AGEMA_signal_16850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9029 ( .C (clk), .D (RoundReg_Inst_ff_SDE_75_next_state), .Q (new_AGEMA_signal_16854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9033 ( .C (clk), .D (new_AGEMA_signal_4135), .Q (new_AGEMA_signal_16858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9037 ( .C (clk), .D (new_AGEMA_signal_4136), .Q (new_AGEMA_signal_16862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9041 ( .C (clk), .D (new_AGEMA_signal_4137), .Q (new_AGEMA_signal_16866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9045 ( .C (clk), .D (RoundReg_Inst_ff_SDE_76_next_state), .Q (new_AGEMA_signal_16870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9049 ( .C (clk), .D (new_AGEMA_signal_4141), .Q (new_AGEMA_signal_16874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9053 ( .C (clk), .D (new_AGEMA_signal_4142), .Q (new_AGEMA_signal_16878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9057 ( .C (clk), .D (new_AGEMA_signal_4143), .Q (new_AGEMA_signal_16882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9061 ( .C (clk), .D (RoundReg_Inst_ff_SDE_77_next_state), .Q (new_AGEMA_signal_16886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9065 ( .C (clk), .D (new_AGEMA_signal_4147), .Q (new_AGEMA_signal_16890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9069 ( .C (clk), .D (new_AGEMA_signal_4148), .Q (new_AGEMA_signal_16894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9073 ( .C (clk), .D (new_AGEMA_signal_4149), .Q (new_AGEMA_signal_16898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9077 ( .C (clk), .D (RoundReg_Inst_ff_SDE_78_next_state), .Q (new_AGEMA_signal_16902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9081 ( .C (clk), .D (new_AGEMA_signal_4153), .Q (new_AGEMA_signal_16906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9085 ( .C (clk), .D (new_AGEMA_signal_4154), .Q (new_AGEMA_signal_16910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9089 ( .C (clk), .D (new_AGEMA_signal_4155), .Q (new_AGEMA_signal_16914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9093 ( .C (clk), .D (RoundReg_Inst_ff_SDE_79_next_state), .Q (new_AGEMA_signal_16918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9097 ( .C (clk), .D (new_AGEMA_signal_4159), .Q (new_AGEMA_signal_16922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9101 ( .C (clk), .D (new_AGEMA_signal_4160), .Q (new_AGEMA_signal_16926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9105 ( .C (clk), .D (new_AGEMA_signal_4161), .Q (new_AGEMA_signal_16930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9109 ( .C (clk), .D (RoundReg_Inst_ff_SDE_80_next_state), .Q (new_AGEMA_signal_16934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9113 ( .C (clk), .D (new_AGEMA_signal_4165), .Q (new_AGEMA_signal_16938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9117 ( .C (clk), .D (new_AGEMA_signal_4166), .Q (new_AGEMA_signal_16942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9121 ( .C (clk), .D (new_AGEMA_signal_4167), .Q (new_AGEMA_signal_16946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9125 ( .C (clk), .D (RoundReg_Inst_ff_SDE_81_next_state), .Q (new_AGEMA_signal_16950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9129 ( .C (clk), .D (new_AGEMA_signal_4171), .Q (new_AGEMA_signal_16954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9133 ( .C (clk), .D (new_AGEMA_signal_4172), .Q (new_AGEMA_signal_16958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9137 ( .C (clk), .D (new_AGEMA_signal_4173), .Q (new_AGEMA_signal_16962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9141 ( .C (clk), .D (RoundReg_Inst_ff_SDE_82_next_state), .Q (new_AGEMA_signal_16966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9145 ( .C (clk), .D (new_AGEMA_signal_4177), .Q (new_AGEMA_signal_16970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9149 ( .C (clk), .D (new_AGEMA_signal_4178), .Q (new_AGEMA_signal_16974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9153 ( .C (clk), .D (new_AGEMA_signal_4179), .Q (new_AGEMA_signal_16978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9157 ( .C (clk), .D (RoundReg_Inst_ff_SDE_83_next_state), .Q (new_AGEMA_signal_16982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9161 ( .C (clk), .D (new_AGEMA_signal_4183), .Q (new_AGEMA_signal_16986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9165 ( .C (clk), .D (new_AGEMA_signal_4184), .Q (new_AGEMA_signal_16990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9169 ( .C (clk), .D (new_AGEMA_signal_4185), .Q (new_AGEMA_signal_16994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9173 ( .C (clk), .D (RoundReg_Inst_ff_SDE_84_next_state), .Q (new_AGEMA_signal_16998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9177 ( .C (clk), .D (new_AGEMA_signal_4189), .Q (new_AGEMA_signal_17002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9181 ( .C (clk), .D (new_AGEMA_signal_4190), .Q (new_AGEMA_signal_17006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9185 ( .C (clk), .D (new_AGEMA_signal_4191), .Q (new_AGEMA_signal_17010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9189 ( .C (clk), .D (RoundReg_Inst_ff_SDE_85_next_state), .Q (new_AGEMA_signal_17014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9193 ( .C (clk), .D (new_AGEMA_signal_4195), .Q (new_AGEMA_signal_17018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9197 ( .C (clk), .D (new_AGEMA_signal_4196), .Q (new_AGEMA_signal_17022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9201 ( .C (clk), .D (new_AGEMA_signal_4197), .Q (new_AGEMA_signal_17026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9205 ( .C (clk), .D (RoundReg_Inst_ff_SDE_86_next_state), .Q (new_AGEMA_signal_17030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9209 ( .C (clk), .D (new_AGEMA_signal_4201), .Q (new_AGEMA_signal_17034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9213 ( .C (clk), .D (new_AGEMA_signal_4202), .Q (new_AGEMA_signal_17038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9217 ( .C (clk), .D (new_AGEMA_signal_4203), .Q (new_AGEMA_signal_17042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9221 ( .C (clk), .D (RoundReg_Inst_ff_SDE_87_next_state), .Q (new_AGEMA_signal_17046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9225 ( .C (clk), .D (new_AGEMA_signal_4207), .Q (new_AGEMA_signal_17050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9229 ( .C (clk), .D (new_AGEMA_signal_4208), .Q (new_AGEMA_signal_17054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9233 ( .C (clk), .D (new_AGEMA_signal_4209), .Q (new_AGEMA_signal_17058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9237 ( .C (clk), .D (RoundReg_Inst_ff_SDE_88_next_state), .Q (new_AGEMA_signal_17062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9241 ( .C (clk), .D (new_AGEMA_signal_4213), .Q (new_AGEMA_signal_17066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9245 ( .C (clk), .D (new_AGEMA_signal_4214), .Q (new_AGEMA_signal_17070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9249 ( .C (clk), .D (new_AGEMA_signal_4215), .Q (new_AGEMA_signal_17074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9253 ( .C (clk), .D (RoundReg_Inst_ff_SDE_89_next_state), .Q (new_AGEMA_signal_17078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9257 ( .C (clk), .D (new_AGEMA_signal_4219), .Q (new_AGEMA_signal_17082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9261 ( .C (clk), .D (new_AGEMA_signal_4220), .Q (new_AGEMA_signal_17086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9265 ( .C (clk), .D (new_AGEMA_signal_4221), .Q (new_AGEMA_signal_17090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9269 ( .C (clk), .D (RoundReg_Inst_ff_SDE_90_next_state), .Q (new_AGEMA_signal_17094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9273 ( .C (clk), .D (new_AGEMA_signal_4225), .Q (new_AGEMA_signal_17098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9277 ( .C (clk), .D (new_AGEMA_signal_4226), .Q (new_AGEMA_signal_17102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9281 ( .C (clk), .D (new_AGEMA_signal_4227), .Q (new_AGEMA_signal_17106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9285 ( .C (clk), .D (RoundReg_Inst_ff_SDE_91_next_state), .Q (new_AGEMA_signal_17110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9289 ( .C (clk), .D (new_AGEMA_signal_4231), .Q (new_AGEMA_signal_17114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9293 ( .C (clk), .D (new_AGEMA_signal_4232), .Q (new_AGEMA_signal_17118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9297 ( .C (clk), .D (new_AGEMA_signal_4233), .Q (new_AGEMA_signal_17122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9301 ( .C (clk), .D (RoundReg_Inst_ff_SDE_92_next_state), .Q (new_AGEMA_signal_17126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9305 ( .C (clk), .D (new_AGEMA_signal_4237), .Q (new_AGEMA_signal_17130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9309 ( .C (clk), .D (new_AGEMA_signal_4238), .Q (new_AGEMA_signal_17134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9313 ( .C (clk), .D (new_AGEMA_signal_4239), .Q (new_AGEMA_signal_17138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9317 ( .C (clk), .D (RoundReg_Inst_ff_SDE_93_next_state), .Q (new_AGEMA_signal_17142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9321 ( .C (clk), .D (new_AGEMA_signal_4243), .Q (new_AGEMA_signal_17146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9325 ( .C (clk), .D (new_AGEMA_signal_4244), .Q (new_AGEMA_signal_17150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9329 ( .C (clk), .D (new_AGEMA_signal_4245), .Q (new_AGEMA_signal_17154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9333 ( .C (clk), .D (RoundReg_Inst_ff_SDE_94_next_state), .Q (new_AGEMA_signal_17158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9337 ( .C (clk), .D (new_AGEMA_signal_4249), .Q (new_AGEMA_signal_17162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9341 ( .C (clk), .D (new_AGEMA_signal_4250), .Q (new_AGEMA_signal_17166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9345 ( .C (clk), .D (new_AGEMA_signal_4251), .Q (new_AGEMA_signal_17170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9349 ( .C (clk), .D (RoundReg_Inst_ff_SDE_95_next_state), .Q (new_AGEMA_signal_17174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9353 ( .C (clk), .D (new_AGEMA_signal_4255), .Q (new_AGEMA_signal_17178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9357 ( .C (clk), .D (new_AGEMA_signal_4256), .Q (new_AGEMA_signal_17182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9361 ( .C (clk), .D (new_AGEMA_signal_4257), .Q (new_AGEMA_signal_17186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9365 ( .C (clk), .D (RoundReg_Inst_ff_SDE_96_next_state), .Q (new_AGEMA_signal_17190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9369 ( .C (clk), .D (new_AGEMA_signal_4261), .Q (new_AGEMA_signal_17194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9373 ( .C (clk), .D (new_AGEMA_signal_4262), .Q (new_AGEMA_signal_17198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9377 ( .C (clk), .D (new_AGEMA_signal_4263), .Q (new_AGEMA_signal_17202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9381 ( .C (clk), .D (RoundReg_Inst_ff_SDE_97_next_state), .Q (new_AGEMA_signal_17206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9385 ( .C (clk), .D (new_AGEMA_signal_4267), .Q (new_AGEMA_signal_17210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9389 ( .C (clk), .D (new_AGEMA_signal_4268), .Q (new_AGEMA_signal_17214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9393 ( .C (clk), .D (new_AGEMA_signal_4269), .Q (new_AGEMA_signal_17218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9397 ( .C (clk), .D (RoundReg_Inst_ff_SDE_98_next_state), .Q (new_AGEMA_signal_17222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9401 ( .C (clk), .D (new_AGEMA_signal_4273), .Q (new_AGEMA_signal_17226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9405 ( .C (clk), .D (new_AGEMA_signal_4274), .Q (new_AGEMA_signal_17230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9409 ( .C (clk), .D (new_AGEMA_signal_4275), .Q (new_AGEMA_signal_17234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9413 ( .C (clk), .D (RoundReg_Inst_ff_SDE_99_next_state), .Q (new_AGEMA_signal_17238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9417 ( .C (clk), .D (new_AGEMA_signal_4279), .Q (new_AGEMA_signal_17242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9421 ( .C (clk), .D (new_AGEMA_signal_4280), .Q (new_AGEMA_signal_17246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9425 ( .C (clk), .D (new_AGEMA_signal_4281), .Q (new_AGEMA_signal_17250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9429 ( .C (clk), .D (RoundReg_Inst_ff_SDE_100_next_state), .Q (new_AGEMA_signal_17254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9433 ( .C (clk), .D (new_AGEMA_signal_4285), .Q (new_AGEMA_signal_17258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9437 ( .C (clk), .D (new_AGEMA_signal_4286), .Q (new_AGEMA_signal_17262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9441 ( .C (clk), .D (new_AGEMA_signal_4287), .Q (new_AGEMA_signal_17266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9445 ( .C (clk), .D (RoundReg_Inst_ff_SDE_101_next_state), .Q (new_AGEMA_signal_17270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9449 ( .C (clk), .D (new_AGEMA_signal_4291), .Q (new_AGEMA_signal_17274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9453 ( .C (clk), .D (new_AGEMA_signal_4292), .Q (new_AGEMA_signal_17278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9457 ( .C (clk), .D (new_AGEMA_signal_4293), .Q (new_AGEMA_signal_17282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9461 ( .C (clk), .D (RoundReg_Inst_ff_SDE_102_next_state), .Q (new_AGEMA_signal_17286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9465 ( .C (clk), .D (new_AGEMA_signal_4297), .Q (new_AGEMA_signal_17290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9469 ( .C (clk), .D (new_AGEMA_signal_4298), .Q (new_AGEMA_signal_17294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9473 ( .C (clk), .D (new_AGEMA_signal_4299), .Q (new_AGEMA_signal_17298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9477 ( .C (clk), .D (RoundReg_Inst_ff_SDE_103_next_state), .Q (new_AGEMA_signal_17302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9481 ( .C (clk), .D (new_AGEMA_signal_4303), .Q (new_AGEMA_signal_17306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9485 ( .C (clk), .D (new_AGEMA_signal_4304), .Q (new_AGEMA_signal_17310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9489 ( .C (clk), .D (new_AGEMA_signal_4305), .Q (new_AGEMA_signal_17314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9493 ( .C (clk), .D (RoundReg_Inst_ff_SDE_104_next_state), .Q (new_AGEMA_signal_17318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9497 ( .C (clk), .D (new_AGEMA_signal_4309), .Q (new_AGEMA_signal_17322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9501 ( .C (clk), .D (new_AGEMA_signal_4310), .Q (new_AGEMA_signal_17326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9505 ( .C (clk), .D (new_AGEMA_signal_4311), .Q (new_AGEMA_signal_17330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9509 ( .C (clk), .D (RoundReg_Inst_ff_SDE_105_next_state), .Q (new_AGEMA_signal_17334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9513 ( .C (clk), .D (new_AGEMA_signal_4315), .Q (new_AGEMA_signal_17338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9517 ( .C (clk), .D (new_AGEMA_signal_4316), .Q (new_AGEMA_signal_17342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9521 ( .C (clk), .D (new_AGEMA_signal_4317), .Q (new_AGEMA_signal_17346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9525 ( .C (clk), .D (RoundReg_Inst_ff_SDE_106_next_state), .Q (new_AGEMA_signal_17350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9529 ( .C (clk), .D (new_AGEMA_signal_4321), .Q (new_AGEMA_signal_17354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9533 ( .C (clk), .D (new_AGEMA_signal_4322), .Q (new_AGEMA_signal_17358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9537 ( .C (clk), .D (new_AGEMA_signal_4323), .Q (new_AGEMA_signal_17362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9541 ( .C (clk), .D (RoundReg_Inst_ff_SDE_107_next_state), .Q (new_AGEMA_signal_17366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9545 ( .C (clk), .D (new_AGEMA_signal_4327), .Q (new_AGEMA_signal_17370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9549 ( .C (clk), .D (new_AGEMA_signal_4328), .Q (new_AGEMA_signal_17374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9553 ( .C (clk), .D (new_AGEMA_signal_4329), .Q (new_AGEMA_signal_17378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9557 ( .C (clk), .D (RoundReg_Inst_ff_SDE_108_next_state), .Q (new_AGEMA_signal_17382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9561 ( .C (clk), .D (new_AGEMA_signal_4333), .Q (new_AGEMA_signal_17386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9565 ( .C (clk), .D (new_AGEMA_signal_4334), .Q (new_AGEMA_signal_17390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9569 ( .C (clk), .D (new_AGEMA_signal_4335), .Q (new_AGEMA_signal_17394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9573 ( .C (clk), .D (RoundReg_Inst_ff_SDE_109_next_state), .Q (new_AGEMA_signal_17398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9577 ( .C (clk), .D (new_AGEMA_signal_4339), .Q (new_AGEMA_signal_17402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9581 ( .C (clk), .D (new_AGEMA_signal_4340), .Q (new_AGEMA_signal_17406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9585 ( .C (clk), .D (new_AGEMA_signal_4341), .Q (new_AGEMA_signal_17410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9589 ( .C (clk), .D (RoundReg_Inst_ff_SDE_110_next_state), .Q (new_AGEMA_signal_17414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9593 ( .C (clk), .D (new_AGEMA_signal_4345), .Q (new_AGEMA_signal_17418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9597 ( .C (clk), .D (new_AGEMA_signal_4346), .Q (new_AGEMA_signal_17422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9601 ( .C (clk), .D (new_AGEMA_signal_4347), .Q (new_AGEMA_signal_17426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9605 ( .C (clk), .D (RoundReg_Inst_ff_SDE_111_next_state), .Q (new_AGEMA_signal_17430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9609 ( .C (clk), .D (new_AGEMA_signal_4351), .Q (new_AGEMA_signal_17434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9613 ( .C (clk), .D (new_AGEMA_signal_4352), .Q (new_AGEMA_signal_17438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9617 ( .C (clk), .D (new_AGEMA_signal_4353), .Q (new_AGEMA_signal_17442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9621 ( .C (clk), .D (RoundReg_Inst_ff_SDE_112_next_state), .Q (new_AGEMA_signal_17446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9625 ( .C (clk), .D (new_AGEMA_signal_4357), .Q (new_AGEMA_signal_17450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9629 ( .C (clk), .D (new_AGEMA_signal_4358), .Q (new_AGEMA_signal_17454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9633 ( .C (clk), .D (new_AGEMA_signal_4359), .Q (new_AGEMA_signal_17458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9637 ( .C (clk), .D (RoundReg_Inst_ff_SDE_113_next_state), .Q (new_AGEMA_signal_17462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9641 ( .C (clk), .D (new_AGEMA_signal_4363), .Q (new_AGEMA_signal_17466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9645 ( .C (clk), .D (new_AGEMA_signal_4364), .Q (new_AGEMA_signal_17470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9649 ( .C (clk), .D (new_AGEMA_signal_4365), .Q (new_AGEMA_signal_17474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9653 ( .C (clk), .D (RoundReg_Inst_ff_SDE_114_next_state), .Q (new_AGEMA_signal_17478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9657 ( .C (clk), .D (new_AGEMA_signal_4369), .Q (new_AGEMA_signal_17482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9661 ( .C (clk), .D (new_AGEMA_signal_4370), .Q (new_AGEMA_signal_17486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9665 ( .C (clk), .D (new_AGEMA_signal_4371), .Q (new_AGEMA_signal_17490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9669 ( .C (clk), .D (RoundReg_Inst_ff_SDE_115_next_state), .Q (new_AGEMA_signal_17494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9673 ( .C (clk), .D (new_AGEMA_signal_4375), .Q (new_AGEMA_signal_17498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9677 ( .C (clk), .D (new_AGEMA_signal_4376), .Q (new_AGEMA_signal_17502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9681 ( .C (clk), .D (new_AGEMA_signal_4377), .Q (new_AGEMA_signal_17506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9685 ( .C (clk), .D (RoundReg_Inst_ff_SDE_116_next_state), .Q (new_AGEMA_signal_17510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9689 ( .C (clk), .D (new_AGEMA_signal_4381), .Q (new_AGEMA_signal_17514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9693 ( .C (clk), .D (new_AGEMA_signal_4382), .Q (new_AGEMA_signal_17518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9697 ( .C (clk), .D (new_AGEMA_signal_4383), .Q (new_AGEMA_signal_17522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9701 ( .C (clk), .D (RoundReg_Inst_ff_SDE_117_next_state), .Q (new_AGEMA_signal_17526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9705 ( .C (clk), .D (new_AGEMA_signal_4387), .Q (new_AGEMA_signal_17530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9709 ( .C (clk), .D (new_AGEMA_signal_4388), .Q (new_AGEMA_signal_17534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9713 ( .C (clk), .D (new_AGEMA_signal_4389), .Q (new_AGEMA_signal_17538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9717 ( .C (clk), .D (RoundReg_Inst_ff_SDE_118_next_state), .Q (new_AGEMA_signal_17542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9721 ( .C (clk), .D (new_AGEMA_signal_4393), .Q (new_AGEMA_signal_17546) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9725 ( .C (clk), .D (new_AGEMA_signal_4394), .Q (new_AGEMA_signal_17550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9729 ( .C (clk), .D (new_AGEMA_signal_4395), .Q (new_AGEMA_signal_17554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9733 ( .C (clk), .D (RoundReg_Inst_ff_SDE_119_next_state), .Q (new_AGEMA_signal_17558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9737 ( .C (clk), .D (new_AGEMA_signal_4399), .Q (new_AGEMA_signal_17562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9741 ( .C (clk), .D (new_AGEMA_signal_4400), .Q (new_AGEMA_signal_17566) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9745 ( .C (clk), .D (new_AGEMA_signal_4401), .Q (new_AGEMA_signal_17570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9749 ( .C (clk), .D (RoundReg_Inst_ff_SDE_120_next_state), .Q (new_AGEMA_signal_17574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9753 ( .C (clk), .D (new_AGEMA_signal_4405), .Q (new_AGEMA_signal_17578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9757 ( .C (clk), .D (new_AGEMA_signal_4406), .Q (new_AGEMA_signal_17582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9761 ( .C (clk), .D (new_AGEMA_signal_4407), .Q (new_AGEMA_signal_17586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9765 ( .C (clk), .D (RoundReg_Inst_ff_SDE_121_next_state), .Q (new_AGEMA_signal_17590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9769 ( .C (clk), .D (new_AGEMA_signal_4411), .Q (new_AGEMA_signal_17594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9773 ( .C (clk), .D (new_AGEMA_signal_4412), .Q (new_AGEMA_signal_17598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9777 ( .C (clk), .D (new_AGEMA_signal_4413), .Q (new_AGEMA_signal_17602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9781 ( .C (clk), .D (RoundReg_Inst_ff_SDE_122_next_state), .Q (new_AGEMA_signal_17606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9785 ( .C (clk), .D (new_AGEMA_signal_4417), .Q (new_AGEMA_signal_17610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9789 ( .C (clk), .D (new_AGEMA_signal_4418), .Q (new_AGEMA_signal_17614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9793 ( .C (clk), .D (new_AGEMA_signal_4419), .Q (new_AGEMA_signal_17618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9797 ( .C (clk), .D (RoundReg_Inst_ff_SDE_123_next_state), .Q (new_AGEMA_signal_17622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9801 ( .C (clk), .D (new_AGEMA_signal_4423), .Q (new_AGEMA_signal_17626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9805 ( .C (clk), .D (new_AGEMA_signal_4424), .Q (new_AGEMA_signal_17630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9809 ( .C (clk), .D (new_AGEMA_signal_4425), .Q (new_AGEMA_signal_17634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9813 ( .C (clk), .D (RoundReg_Inst_ff_SDE_124_next_state), .Q (new_AGEMA_signal_17638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9817 ( .C (clk), .D (new_AGEMA_signal_4429), .Q (new_AGEMA_signal_17642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9821 ( .C (clk), .D (new_AGEMA_signal_4430), .Q (new_AGEMA_signal_17646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9825 ( .C (clk), .D (new_AGEMA_signal_4431), .Q (new_AGEMA_signal_17650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9829 ( .C (clk), .D (RoundReg_Inst_ff_SDE_125_next_state), .Q (new_AGEMA_signal_17654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9833 ( .C (clk), .D (new_AGEMA_signal_4435), .Q (new_AGEMA_signal_17658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9837 ( .C (clk), .D (new_AGEMA_signal_4436), .Q (new_AGEMA_signal_17662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9841 ( .C (clk), .D (new_AGEMA_signal_4437), .Q (new_AGEMA_signal_17666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9845 ( .C (clk), .D (RoundReg_Inst_ff_SDE_126_next_state), .Q (new_AGEMA_signal_17670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9849 ( .C (clk), .D (new_AGEMA_signal_4441), .Q (new_AGEMA_signal_17674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9853 ( .C (clk), .D (new_AGEMA_signal_4442), .Q (new_AGEMA_signal_17678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9857 ( .C (clk), .D (new_AGEMA_signal_4443), .Q (new_AGEMA_signal_17682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9861 ( .C (clk), .D (RoundReg_Inst_ff_SDE_127_next_state), .Q (new_AGEMA_signal_17686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9865 ( .C (clk), .D (new_AGEMA_signal_4447), .Q (new_AGEMA_signal_17690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9869 ( .C (clk), .D (new_AGEMA_signal_4448), .Q (new_AGEMA_signal_17694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9873 ( .C (clk), .D (new_AGEMA_signal_4449), .Q (new_AGEMA_signal_17698) ) ;
    buf_clk new_AGEMA_reg_buffer_9877 ( .C (clk), .D (RoundCounterIns_n45), .Q (new_AGEMA_signal_17702) ) ;
    buf_clk new_AGEMA_reg_buffer_9881 ( .C (clk), .D (RoundCounterIns_n44), .Q (new_AGEMA_signal_17706) ) ;
    buf_clk new_AGEMA_reg_buffer_9885 ( .C (clk), .D (RoundCounterIns_n1), .Q (new_AGEMA_signal_17710) ) ;
    buf_clk new_AGEMA_reg_buffer_9889 ( .C (clk), .D (RoundCounterIns_n42), .Q (new_AGEMA_signal_17714) ) ;
    buf_clk new_AGEMA_reg_buffer_9893 ( .C (clk), .D (InRoundCounterIns_n41), .Q (new_AGEMA_signal_17718) ) ;
    buf_clk new_AGEMA_reg_buffer_9897 ( .C (clk), .D (InRoundCounterIns_n40), .Q (new_AGEMA_signal_17722) ) ;
    buf_clk new_AGEMA_reg_buffer_9901 ( .C (clk), .D (InRoundCounterIns_n39), .Q (new_AGEMA_signal_17726) ) ;

    /* cells in depth 2 */
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, new_AGEMA_signal_4999, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, new_AGEMA_signal_4993, SubBytesIns_Inst_Sbox_0_M20}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_5043, new_AGEMA_signal_5042, new_AGEMA_signal_5041, SubBytesIns_Inst_Sbox_0_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_9953, new_AGEMA_signal_9952, new_AGEMA_signal_9951, new_AGEMA_signal_9950}), .b ({new_AGEMA_signal_5043, new_AGEMA_signal_5042, new_AGEMA_signal_5041, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_5091, new_AGEMA_signal_5090, new_AGEMA_signal_5089, SubBytesIns_Inst_Sbox_0_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_9957, new_AGEMA_signal_9956, new_AGEMA_signal_9955, new_AGEMA_signal_9954}), .b ({new_AGEMA_signal_5043, new_AGEMA_signal_5042, new_AGEMA_signal_5041, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_5094, new_AGEMA_signal_5093, new_AGEMA_signal_5092, SubBytesIns_Inst_Sbox_0_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, new_AGEMA_signal_4993, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_5040, new_AGEMA_signal_5039, new_AGEMA_signal_5038, SubBytesIns_Inst_Sbox_0_M23}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450], Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_5097, new_AGEMA_signal_5096, new_AGEMA_signal_5095, SubBytesIns_Inst_Sbox_0_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_9961, new_AGEMA_signal_9960, new_AGEMA_signal_9959, new_AGEMA_signal_9958}), .b ({new_AGEMA_signal_5043, new_AGEMA_signal_5042, new_AGEMA_signal_5041, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_5100, new_AGEMA_signal_5099, new_AGEMA_signal_5098, SubBytesIns_Inst_Sbox_0_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_4998, new_AGEMA_signal_4997, new_AGEMA_signal_4996, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, new_AGEMA_signal_4999, SubBytesIns_Inst_Sbox_0_M22}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462], Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, new_AGEMA_signal_5047, SubBytesIns_Inst_Sbox_0_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_9965, new_AGEMA_signal_9964, new_AGEMA_signal_9963, new_AGEMA_signal_9962}), .b ({new_AGEMA_signal_5043, new_AGEMA_signal_5042, new_AGEMA_signal_5041, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_5160, new_AGEMA_signal_5159, new_AGEMA_signal_5158, SubBytesIns_Inst_Sbox_0_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, new_AGEMA_signal_5011, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_5007, new_AGEMA_signal_5006, new_AGEMA_signal_5005, SubBytesIns_Inst_Sbox_1_M20}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, new_AGEMA_signal_5053, SubBytesIns_Inst_Sbox_1_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_9969, new_AGEMA_signal_9968, new_AGEMA_signal_9967, new_AGEMA_signal_9966}), .b ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, new_AGEMA_signal_5053, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_5106, new_AGEMA_signal_5105, new_AGEMA_signal_5104, SubBytesIns_Inst_Sbox_1_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_9973, new_AGEMA_signal_9972, new_AGEMA_signal_9971, new_AGEMA_signal_9970}), .b ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, new_AGEMA_signal_5053, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_5109, new_AGEMA_signal_5108, new_AGEMA_signal_5107, SubBytesIns_Inst_Sbox_1_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_5007, new_AGEMA_signal_5006, new_AGEMA_signal_5005, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_5052, new_AGEMA_signal_5051, new_AGEMA_signal_5050, SubBytesIns_Inst_Sbox_1_M23}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_5112, new_AGEMA_signal_5111, new_AGEMA_signal_5110, SubBytesIns_Inst_Sbox_1_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_9977, new_AGEMA_signal_9976, new_AGEMA_signal_9975, new_AGEMA_signal_9974}), .b ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, new_AGEMA_signal_5053, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_5115, new_AGEMA_signal_5114, new_AGEMA_signal_5113, SubBytesIns_Inst_Sbox_1_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_5010, new_AGEMA_signal_5009, new_AGEMA_signal_5008, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, new_AGEMA_signal_5011, SubBytesIns_Inst_Sbox_1_M22}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498], Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_5061, new_AGEMA_signal_5060, new_AGEMA_signal_5059, SubBytesIns_Inst_Sbox_1_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_9981, new_AGEMA_signal_9980, new_AGEMA_signal_9979, new_AGEMA_signal_9978}), .b ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, new_AGEMA_signal_5053, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_5175, new_AGEMA_signal_5174, new_AGEMA_signal_5173, SubBytesIns_Inst_Sbox_1_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_5025, new_AGEMA_signal_5024, new_AGEMA_signal_5023, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, new_AGEMA_signal_5017, SubBytesIns_Inst_Sbox_2_M20}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510], Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, new_AGEMA_signal_5065, SubBytesIns_Inst_Sbox_2_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_9985, new_AGEMA_signal_9984, new_AGEMA_signal_9983, new_AGEMA_signal_9982}), .b ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, new_AGEMA_signal_5065, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_5121, new_AGEMA_signal_5120, new_AGEMA_signal_5119, SubBytesIns_Inst_Sbox_2_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_9989, new_AGEMA_signal_9988, new_AGEMA_signal_9987, new_AGEMA_signal_9986}), .b ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, new_AGEMA_signal_5065, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_5124, new_AGEMA_signal_5123, new_AGEMA_signal_5122, SubBytesIns_Inst_Sbox_2_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, new_AGEMA_signal_5017, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_5064, new_AGEMA_signal_5063, new_AGEMA_signal_5062, SubBytesIns_Inst_Sbox_2_M23}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_5127, new_AGEMA_signal_5126, new_AGEMA_signal_5125, SubBytesIns_Inst_Sbox_2_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_9993, new_AGEMA_signal_9992, new_AGEMA_signal_9991, new_AGEMA_signal_9990}), .b ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, new_AGEMA_signal_5065, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_5130, new_AGEMA_signal_5129, new_AGEMA_signal_5128, SubBytesIns_Inst_Sbox_2_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_5025, new_AGEMA_signal_5024, new_AGEMA_signal_5023, SubBytesIns_Inst_Sbox_2_M22}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_5073, new_AGEMA_signal_5072, new_AGEMA_signal_5071, SubBytesIns_Inst_Sbox_2_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_9997, new_AGEMA_signal_9996, new_AGEMA_signal_9995, new_AGEMA_signal_9994}), .b ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, new_AGEMA_signal_5065, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_5190, new_AGEMA_signal_5189, new_AGEMA_signal_5188, SubBytesIns_Inst_Sbox_2_M36}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, new_AGEMA_signal_5035, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, new_AGEMA_signal_5029, SubBytesIns_Inst_Sbox_3_M20}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_5079, new_AGEMA_signal_5078, new_AGEMA_signal_5077, SubBytesIns_Inst_Sbox_3_M25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_10001, new_AGEMA_signal_10000, new_AGEMA_signal_9999, new_AGEMA_signal_9998}), .b ({new_AGEMA_signal_5079, new_AGEMA_signal_5078, new_AGEMA_signal_5077, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_5136, new_AGEMA_signal_5135, new_AGEMA_signal_5134, SubBytesIns_Inst_Sbox_3_M26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_10005, new_AGEMA_signal_10004, new_AGEMA_signal_10003, new_AGEMA_signal_10002}), .b ({new_AGEMA_signal_5079, new_AGEMA_signal_5078, new_AGEMA_signal_5077, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_5139, new_AGEMA_signal_5138, new_AGEMA_signal_5137, SubBytesIns_Inst_Sbox_3_M28}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, new_AGEMA_signal_5029, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_5076, new_AGEMA_signal_5075, new_AGEMA_signal_5074, SubBytesIns_Inst_Sbox_3_M23}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_5142, new_AGEMA_signal_5141, new_AGEMA_signal_5140, SubBytesIns_Inst_Sbox_3_M31}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_10009, new_AGEMA_signal_10008, new_AGEMA_signal_10007, new_AGEMA_signal_10006}), .b ({new_AGEMA_signal_5079, new_AGEMA_signal_5078, new_AGEMA_signal_5077, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_5145, new_AGEMA_signal_5144, new_AGEMA_signal_5143, SubBytesIns_Inst_Sbox_3_M33}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_5034, new_AGEMA_signal_5033, new_AGEMA_signal_5032, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, new_AGEMA_signal_5035, SubBytesIns_Inst_Sbox_3_M22}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570], Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_5085, new_AGEMA_signal_5084, new_AGEMA_signal_5083, SubBytesIns_Inst_Sbox_3_M34}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_10013, new_AGEMA_signal_10012, new_AGEMA_signal_10011, new_AGEMA_signal_10010}), .b ({new_AGEMA_signal_5079, new_AGEMA_signal_5078, new_AGEMA_signal_5077, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_5205, new_AGEMA_signal_5204, new_AGEMA_signal_5203, SubBytesIns_Inst_Sbox_3_M36}) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2125 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M21), .Q (new_AGEMA_signal_9950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2126 ( .C (clk), .D (new_AGEMA_signal_4996), .Q (new_AGEMA_signal_9951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2127 ( .C (clk), .D (new_AGEMA_signal_4997), .Q (new_AGEMA_signal_9952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2128 ( .C (clk), .D (new_AGEMA_signal_4998), .Q (new_AGEMA_signal_9953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2129 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M23), .Q (new_AGEMA_signal_9954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2130 ( .C (clk), .D (new_AGEMA_signal_5038), .Q (new_AGEMA_signal_9955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2131 ( .C (clk), .D (new_AGEMA_signal_5039), .Q (new_AGEMA_signal_9956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2132 ( .C (clk), .D (new_AGEMA_signal_5040), .Q (new_AGEMA_signal_9957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2133 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M27), .Q (new_AGEMA_signal_9958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2134 ( .C (clk), .D (new_AGEMA_signal_5044), .Q (new_AGEMA_signal_9959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2135 ( .C (clk), .D (new_AGEMA_signal_5045), .Q (new_AGEMA_signal_9960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2136 ( .C (clk), .D (new_AGEMA_signal_5046), .Q (new_AGEMA_signal_9961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2137 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M24), .Q (new_AGEMA_signal_9962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2138 ( .C (clk), .D (new_AGEMA_signal_5086), .Q (new_AGEMA_signal_9963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2139 ( .C (clk), .D (new_AGEMA_signal_5087), .Q (new_AGEMA_signal_9964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2140 ( .C (clk), .D (new_AGEMA_signal_5088), .Q (new_AGEMA_signal_9965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2141 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M21), .Q (new_AGEMA_signal_9966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2142 ( .C (clk), .D (new_AGEMA_signal_5008), .Q (new_AGEMA_signal_9967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2143 ( .C (clk), .D (new_AGEMA_signal_5009), .Q (new_AGEMA_signal_9968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2144 ( .C (clk), .D (new_AGEMA_signal_5010), .Q (new_AGEMA_signal_9969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2145 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M23), .Q (new_AGEMA_signal_9970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2146 ( .C (clk), .D (new_AGEMA_signal_5050), .Q (new_AGEMA_signal_9971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2147 ( .C (clk), .D (new_AGEMA_signal_5051), .Q (new_AGEMA_signal_9972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2148 ( .C (clk), .D (new_AGEMA_signal_5052), .Q (new_AGEMA_signal_9973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2149 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M27), .Q (new_AGEMA_signal_9974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2150 ( .C (clk), .D (new_AGEMA_signal_5056), .Q (new_AGEMA_signal_9975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2151 ( .C (clk), .D (new_AGEMA_signal_5057), .Q (new_AGEMA_signal_9976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2152 ( .C (clk), .D (new_AGEMA_signal_5058), .Q (new_AGEMA_signal_9977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2153 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M24), .Q (new_AGEMA_signal_9978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2154 ( .C (clk), .D (new_AGEMA_signal_5101), .Q (new_AGEMA_signal_9979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2155 ( .C (clk), .D (new_AGEMA_signal_5102), .Q (new_AGEMA_signal_9980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2156 ( .C (clk), .D (new_AGEMA_signal_5103), .Q (new_AGEMA_signal_9981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2157 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M21), .Q (new_AGEMA_signal_9982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2158 ( .C (clk), .D (new_AGEMA_signal_5020), .Q (new_AGEMA_signal_9983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2159 ( .C (clk), .D (new_AGEMA_signal_5021), .Q (new_AGEMA_signal_9984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2160 ( .C (clk), .D (new_AGEMA_signal_5022), .Q (new_AGEMA_signal_9985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2161 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M23), .Q (new_AGEMA_signal_9986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2162 ( .C (clk), .D (new_AGEMA_signal_5062), .Q (new_AGEMA_signal_9987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2163 ( .C (clk), .D (new_AGEMA_signal_5063), .Q (new_AGEMA_signal_9988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2164 ( .C (clk), .D (new_AGEMA_signal_5064), .Q (new_AGEMA_signal_9989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2165 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M27), .Q (new_AGEMA_signal_9990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2166 ( .C (clk), .D (new_AGEMA_signal_5068), .Q (new_AGEMA_signal_9991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2167 ( .C (clk), .D (new_AGEMA_signal_5069), .Q (new_AGEMA_signal_9992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2168 ( .C (clk), .D (new_AGEMA_signal_5070), .Q (new_AGEMA_signal_9993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2169 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M24), .Q (new_AGEMA_signal_9994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2170 ( .C (clk), .D (new_AGEMA_signal_5116), .Q (new_AGEMA_signal_9995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2171 ( .C (clk), .D (new_AGEMA_signal_5117), .Q (new_AGEMA_signal_9996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2172 ( .C (clk), .D (new_AGEMA_signal_5118), .Q (new_AGEMA_signal_9997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2173 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M21), .Q (new_AGEMA_signal_9998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2174 ( .C (clk), .D (new_AGEMA_signal_5032), .Q (new_AGEMA_signal_9999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2175 ( .C (clk), .D (new_AGEMA_signal_5033), .Q (new_AGEMA_signal_10000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2176 ( .C (clk), .D (new_AGEMA_signal_5034), .Q (new_AGEMA_signal_10001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2177 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M23), .Q (new_AGEMA_signal_10002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2178 ( .C (clk), .D (new_AGEMA_signal_5074), .Q (new_AGEMA_signal_10003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2179 ( .C (clk), .D (new_AGEMA_signal_5075), .Q (new_AGEMA_signal_10004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2180 ( .C (clk), .D (new_AGEMA_signal_5076), .Q (new_AGEMA_signal_10005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2181 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M27), .Q (new_AGEMA_signal_10006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2182 ( .C (clk), .D (new_AGEMA_signal_5080), .Q (new_AGEMA_signal_10007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2183 ( .C (clk), .D (new_AGEMA_signal_5081), .Q (new_AGEMA_signal_10008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2184 ( .C (clk), .D (new_AGEMA_signal_5082), .Q (new_AGEMA_signal_10009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2185 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M24), .Q (new_AGEMA_signal_10010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2186 ( .C (clk), .D (new_AGEMA_signal_5131), .Q (new_AGEMA_signal_10011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2187 ( .C (clk), .D (new_AGEMA_signal_5132), .Q (new_AGEMA_signal_10012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2188 ( .C (clk), .D (new_AGEMA_signal_5133), .Q (new_AGEMA_signal_10013) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C (clk), .D (new_AGEMA_signal_10078), .Q (new_AGEMA_signal_10079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2258 ( .C (clk), .D (new_AGEMA_signal_10082), .Q (new_AGEMA_signal_10083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2262 ( .C (clk), .D (new_AGEMA_signal_10086), .Q (new_AGEMA_signal_10087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2266 ( .C (clk), .D (new_AGEMA_signal_10090), .Q (new_AGEMA_signal_10091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2270 ( .C (clk), .D (new_AGEMA_signal_10094), .Q (new_AGEMA_signal_10095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2274 ( .C (clk), .D (new_AGEMA_signal_10098), .Q (new_AGEMA_signal_10099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2278 ( .C (clk), .D (new_AGEMA_signal_10102), .Q (new_AGEMA_signal_10103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2282 ( .C (clk), .D (new_AGEMA_signal_10106), .Q (new_AGEMA_signal_10107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2286 ( .C (clk), .D (new_AGEMA_signal_10110), .Q (new_AGEMA_signal_10111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2290 ( .C (clk), .D (new_AGEMA_signal_10114), .Q (new_AGEMA_signal_10115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2294 ( .C (clk), .D (new_AGEMA_signal_10118), .Q (new_AGEMA_signal_10119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2298 ( .C (clk), .D (new_AGEMA_signal_10122), .Q (new_AGEMA_signal_10123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2302 ( .C (clk), .D (new_AGEMA_signal_10126), .Q (new_AGEMA_signal_10127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2306 ( .C (clk), .D (new_AGEMA_signal_10130), .Q (new_AGEMA_signal_10131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2310 ( .C (clk), .D (new_AGEMA_signal_10134), .Q (new_AGEMA_signal_10135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2314 ( .C (clk), .D (new_AGEMA_signal_10138), .Q (new_AGEMA_signal_10139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2318 ( .C (clk), .D (new_AGEMA_signal_10142), .Q (new_AGEMA_signal_10143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2322 ( .C (clk), .D (new_AGEMA_signal_10146), .Q (new_AGEMA_signal_10147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2326 ( .C (clk), .D (new_AGEMA_signal_10150), .Q (new_AGEMA_signal_10151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2330 ( .C (clk), .D (new_AGEMA_signal_10154), .Q (new_AGEMA_signal_10155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2334 ( .C (clk), .D (new_AGEMA_signal_10158), .Q (new_AGEMA_signal_10159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2338 ( .C (clk), .D (new_AGEMA_signal_10162), .Q (new_AGEMA_signal_10163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2342 ( .C (clk), .D (new_AGEMA_signal_10166), .Q (new_AGEMA_signal_10167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2346 ( .C (clk), .D (new_AGEMA_signal_10170), .Q (new_AGEMA_signal_10171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2350 ( .C (clk), .D (new_AGEMA_signal_10174), .Q (new_AGEMA_signal_10175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2354 ( .C (clk), .D (new_AGEMA_signal_10178), .Q (new_AGEMA_signal_10179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2358 ( .C (clk), .D (new_AGEMA_signal_10182), .Q (new_AGEMA_signal_10183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2362 ( .C (clk), .D (new_AGEMA_signal_10186), .Q (new_AGEMA_signal_10187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2366 ( .C (clk), .D (new_AGEMA_signal_10190), .Q (new_AGEMA_signal_10191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2370 ( .C (clk), .D (new_AGEMA_signal_10194), .Q (new_AGEMA_signal_10195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2374 ( .C (clk), .D (new_AGEMA_signal_10198), .Q (new_AGEMA_signal_10199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2378 ( .C (clk), .D (new_AGEMA_signal_10202), .Q (new_AGEMA_signal_10203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2382 ( .C (clk), .D (new_AGEMA_signal_10206), .Q (new_AGEMA_signal_10207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2386 ( .C (clk), .D (new_AGEMA_signal_10210), .Q (new_AGEMA_signal_10211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2390 ( .C (clk), .D (new_AGEMA_signal_10214), .Q (new_AGEMA_signal_10215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2394 ( .C (clk), .D (new_AGEMA_signal_10218), .Q (new_AGEMA_signal_10219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2398 ( .C (clk), .D (new_AGEMA_signal_10222), .Q (new_AGEMA_signal_10223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2402 ( .C (clk), .D (new_AGEMA_signal_10226), .Q (new_AGEMA_signal_10227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2406 ( .C (clk), .D (new_AGEMA_signal_10230), .Q (new_AGEMA_signal_10231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2410 ( .C (clk), .D (new_AGEMA_signal_10234), .Q (new_AGEMA_signal_10235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2414 ( .C (clk), .D (new_AGEMA_signal_10238), .Q (new_AGEMA_signal_10239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2418 ( .C (clk), .D (new_AGEMA_signal_10242), .Q (new_AGEMA_signal_10243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2422 ( .C (clk), .D (new_AGEMA_signal_10246), .Q (new_AGEMA_signal_10247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2426 ( .C (clk), .D (new_AGEMA_signal_10250), .Q (new_AGEMA_signal_10251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2430 ( .C (clk), .D (new_AGEMA_signal_10254), .Q (new_AGEMA_signal_10255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2434 ( .C (clk), .D (new_AGEMA_signal_10258), .Q (new_AGEMA_signal_10259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2438 ( .C (clk), .D (new_AGEMA_signal_10262), .Q (new_AGEMA_signal_10263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2442 ( .C (clk), .D (new_AGEMA_signal_10266), .Q (new_AGEMA_signal_10267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2446 ( .C (clk), .D (new_AGEMA_signal_10270), .Q (new_AGEMA_signal_10271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2450 ( .C (clk), .D (new_AGEMA_signal_10274), .Q (new_AGEMA_signal_10275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2454 ( .C (clk), .D (new_AGEMA_signal_10278), .Q (new_AGEMA_signal_10279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2458 ( .C (clk), .D (new_AGEMA_signal_10282), .Q (new_AGEMA_signal_10283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2462 ( .C (clk), .D (new_AGEMA_signal_10286), .Q (new_AGEMA_signal_10287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2466 ( .C (clk), .D (new_AGEMA_signal_10290), .Q (new_AGEMA_signal_10291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2470 ( .C (clk), .D (new_AGEMA_signal_10294), .Q (new_AGEMA_signal_10295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2474 ( .C (clk), .D (new_AGEMA_signal_10298), .Q (new_AGEMA_signal_10299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2478 ( .C (clk), .D (new_AGEMA_signal_10302), .Q (new_AGEMA_signal_10303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2482 ( .C (clk), .D (new_AGEMA_signal_10306), .Q (new_AGEMA_signal_10307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2486 ( .C (clk), .D (new_AGEMA_signal_10310), .Q (new_AGEMA_signal_10311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2490 ( .C (clk), .D (new_AGEMA_signal_10314), .Q (new_AGEMA_signal_10315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2494 ( .C (clk), .D (new_AGEMA_signal_10318), .Q (new_AGEMA_signal_10319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2498 ( .C (clk), .D (new_AGEMA_signal_10322), .Q (new_AGEMA_signal_10323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2502 ( .C (clk), .D (new_AGEMA_signal_10326), .Q (new_AGEMA_signal_10327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2506 ( .C (clk), .D (new_AGEMA_signal_10330), .Q (new_AGEMA_signal_10331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2510 ( .C (clk), .D (new_AGEMA_signal_10334), .Q (new_AGEMA_signal_10335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2514 ( .C (clk), .D (new_AGEMA_signal_10338), .Q (new_AGEMA_signal_10339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2518 ( .C (clk), .D (new_AGEMA_signal_10342), .Q (new_AGEMA_signal_10343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2522 ( .C (clk), .D (new_AGEMA_signal_10346), .Q (new_AGEMA_signal_10347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2526 ( .C (clk), .D (new_AGEMA_signal_10350), .Q (new_AGEMA_signal_10351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2530 ( .C (clk), .D (new_AGEMA_signal_10354), .Q (new_AGEMA_signal_10355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2534 ( .C (clk), .D (new_AGEMA_signal_10358), .Q (new_AGEMA_signal_10359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2538 ( .C (clk), .D (new_AGEMA_signal_10362), .Q (new_AGEMA_signal_10363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2542 ( .C (clk), .D (new_AGEMA_signal_10366), .Q (new_AGEMA_signal_10367) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2546 ( .C (clk), .D (new_AGEMA_signal_10370), .Q (new_AGEMA_signal_10371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2550 ( .C (clk), .D (new_AGEMA_signal_10374), .Q (new_AGEMA_signal_10375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2554 ( .C (clk), .D (new_AGEMA_signal_10378), .Q (new_AGEMA_signal_10379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2558 ( .C (clk), .D (new_AGEMA_signal_10382), .Q (new_AGEMA_signal_10383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2562 ( .C (clk), .D (new_AGEMA_signal_10386), .Q (new_AGEMA_signal_10387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2566 ( .C (clk), .D (new_AGEMA_signal_10390), .Q (new_AGEMA_signal_10391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2570 ( .C (clk), .D (new_AGEMA_signal_10394), .Q (new_AGEMA_signal_10395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2574 ( .C (clk), .D (new_AGEMA_signal_10398), .Q (new_AGEMA_signal_10399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2578 ( .C (clk), .D (new_AGEMA_signal_10402), .Q (new_AGEMA_signal_10403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2582 ( .C (clk), .D (new_AGEMA_signal_10406), .Q (new_AGEMA_signal_10407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2586 ( .C (clk), .D (new_AGEMA_signal_10410), .Q (new_AGEMA_signal_10411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2590 ( .C (clk), .D (new_AGEMA_signal_10414), .Q (new_AGEMA_signal_10415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2594 ( .C (clk), .D (new_AGEMA_signal_10418), .Q (new_AGEMA_signal_10419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2598 ( .C (clk), .D (new_AGEMA_signal_10422), .Q (new_AGEMA_signal_10423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2602 ( .C (clk), .D (new_AGEMA_signal_10426), .Q (new_AGEMA_signal_10427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2606 ( .C (clk), .D (new_AGEMA_signal_10430), .Q (new_AGEMA_signal_10431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2610 ( .C (clk), .D (new_AGEMA_signal_10434), .Q (new_AGEMA_signal_10435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2614 ( .C (clk), .D (new_AGEMA_signal_10438), .Q (new_AGEMA_signal_10439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2618 ( .C (clk), .D (new_AGEMA_signal_10442), .Q (new_AGEMA_signal_10443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2622 ( .C (clk), .D (new_AGEMA_signal_10446), .Q (new_AGEMA_signal_10447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2626 ( .C (clk), .D (new_AGEMA_signal_10450), .Q (new_AGEMA_signal_10451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2630 ( .C (clk), .D (new_AGEMA_signal_10454), .Q (new_AGEMA_signal_10455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2634 ( .C (clk), .D (new_AGEMA_signal_10458), .Q (new_AGEMA_signal_10459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2638 ( .C (clk), .D (new_AGEMA_signal_10462), .Q (new_AGEMA_signal_10463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2642 ( .C (clk), .D (new_AGEMA_signal_10466), .Q (new_AGEMA_signal_10467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2646 ( .C (clk), .D (new_AGEMA_signal_10470), .Q (new_AGEMA_signal_10471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2650 ( .C (clk), .D (new_AGEMA_signal_10474), .Q (new_AGEMA_signal_10475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2654 ( .C (clk), .D (new_AGEMA_signal_10478), .Q (new_AGEMA_signal_10479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2658 ( .C (clk), .D (new_AGEMA_signal_10482), .Q (new_AGEMA_signal_10483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2662 ( .C (clk), .D (new_AGEMA_signal_10486), .Q (new_AGEMA_signal_10487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2666 ( .C (clk), .D (new_AGEMA_signal_10490), .Q (new_AGEMA_signal_10491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2670 ( .C (clk), .D (new_AGEMA_signal_10494), .Q (new_AGEMA_signal_10495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2674 ( .C (clk), .D (new_AGEMA_signal_10498), .Q (new_AGEMA_signal_10499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2678 ( .C (clk), .D (new_AGEMA_signal_10502), .Q (new_AGEMA_signal_10503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2682 ( .C (clk), .D (new_AGEMA_signal_10506), .Q (new_AGEMA_signal_10507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2686 ( .C (clk), .D (new_AGEMA_signal_10510), .Q (new_AGEMA_signal_10511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2690 ( .C (clk), .D (new_AGEMA_signal_10514), .Q (new_AGEMA_signal_10515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2694 ( .C (clk), .D (new_AGEMA_signal_10518), .Q (new_AGEMA_signal_10519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2698 ( .C (clk), .D (new_AGEMA_signal_10522), .Q (new_AGEMA_signal_10523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2702 ( .C (clk), .D (new_AGEMA_signal_10526), .Q (new_AGEMA_signal_10527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2706 ( .C (clk), .D (new_AGEMA_signal_10530), .Q (new_AGEMA_signal_10531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2710 ( .C (clk), .D (new_AGEMA_signal_10534), .Q (new_AGEMA_signal_10535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2714 ( .C (clk), .D (new_AGEMA_signal_10538), .Q (new_AGEMA_signal_10539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2718 ( .C (clk), .D (new_AGEMA_signal_10542), .Q (new_AGEMA_signal_10543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2722 ( .C (clk), .D (new_AGEMA_signal_10546), .Q (new_AGEMA_signal_10547) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2726 ( .C (clk), .D (new_AGEMA_signal_10550), .Q (new_AGEMA_signal_10551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2730 ( .C (clk), .D (new_AGEMA_signal_10554), .Q (new_AGEMA_signal_10555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2734 ( .C (clk), .D (new_AGEMA_signal_10558), .Q (new_AGEMA_signal_10559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2738 ( .C (clk), .D (new_AGEMA_signal_10562), .Q (new_AGEMA_signal_10563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2742 ( .C (clk), .D (new_AGEMA_signal_10566), .Q (new_AGEMA_signal_10567) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2746 ( .C (clk), .D (new_AGEMA_signal_10570), .Q (new_AGEMA_signal_10571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2750 ( .C (clk), .D (new_AGEMA_signal_10574), .Q (new_AGEMA_signal_10575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2754 ( .C (clk), .D (new_AGEMA_signal_10578), .Q (new_AGEMA_signal_10579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2758 ( .C (clk), .D (new_AGEMA_signal_10582), .Q (new_AGEMA_signal_10583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2762 ( .C (clk), .D (new_AGEMA_signal_10586), .Q (new_AGEMA_signal_10587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2766 ( .C (clk), .D (new_AGEMA_signal_10590), .Q (new_AGEMA_signal_10591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2770 ( .C (clk), .D (new_AGEMA_signal_10594), .Q (new_AGEMA_signal_10595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2773 ( .C (clk), .D (new_AGEMA_signal_10597), .Q (new_AGEMA_signal_10598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2776 ( .C (clk), .D (new_AGEMA_signal_10600), .Q (new_AGEMA_signal_10601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2779 ( .C (clk), .D (new_AGEMA_signal_10603), .Q (new_AGEMA_signal_10604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2782 ( .C (clk), .D (new_AGEMA_signal_10606), .Q (new_AGEMA_signal_10607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2785 ( .C (clk), .D (new_AGEMA_signal_10609), .Q (new_AGEMA_signal_10610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2788 ( .C (clk), .D (new_AGEMA_signal_10612), .Q (new_AGEMA_signal_10613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2791 ( .C (clk), .D (new_AGEMA_signal_10615), .Q (new_AGEMA_signal_10616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2794 ( .C (clk), .D (new_AGEMA_signal_10618), .Q (new_AGEMA_signal_10619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2797 ( .C (clk), .D (new_AGEMA_signal_10621), .Q (new_AGEMA_signal_10622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2800 ( .C (clk), .D (new_AGEMA_signal_10624), .Q (new_AGEMA_signal_10625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2803 ( .C (clk), .D (new_AGEMA_signal_10627), .Q (new_AGEMA_signal_10628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2806 ( .C (clk), .D (new_AGEMA_signal_10630), .Q (new_AGEMA_signal_10631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2809 ( .C (clk), .D (new_AGEMA_signal_10633), .Q (new_AGEMA_signal_10634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2812 ( .C (clk), .D (new_AGEMA_signal_10636), .Q (new_AGEMA_signal_10637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2815 ( .C (clk), .D (new_AGEMA_signal_10639), .Q (new_AGEMA_signal_10640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2818 ( .C (clk), .D (new_AGEMA_signal_10642), .Q (new_AGEMA_signal_10643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2821 ( .C (clk), .D (new_AGEMA_signal_10645), .Q (new_AGEMA_signal_10646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2824 ( .C (clk), .D (new_AGEMA_signal_10648), .Q (new_AGEMA_signal_10649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2827 ( .C (clk), .D (new_AGEMA_signal_10651), .Q (new_AGEMA_signal_10652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2830 ( .C (clk), .D (new_AGEMA_signal_10654), .Q (new_AGEMA_signal_10655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2833 ( .C (clk), .D (new_AGEMA_signal_10657), .Q (new_AGEMA_signal_10658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2836 ( .C (clk), .D (new_AGEMA_signal_10660), .Q (new_AGEMA_signal_10661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2839 ( .C (clk), .D (new_AGEMA_signal_10663), .Q (new_AGEMA_signal_10664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2842 ( .C (clk), .D (new_AGEMA_signal_10666), .Q (new_AGEMA_signal_10667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2845 ( .C (clk), .D (new_AGEMA_signal_10669), .Q (new_AGEMA_signal_10670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2848 ( .C (clk), .D (new_AGEMA_signal_10672), .Q (new_AGEMA_signal_10673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2851 ( .C (clk), .D (new_AGEMA_signal_10675), .Q (new_AGEMA_signal_10676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2854 ( .C (clk), .D (new_AGEMA_signal_10678), .Q (new_AGEMA_signal_10679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2857 ( .C (clk), .D (new_AGEMA_signal_10681), .Q (new_AGEMA_signal_10682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2860 ( .C (clk), .D (new_AGEMA_signal_10684), .Q (new_AGEMA_signal_10685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2863 ( .C (clk), .D (new_AGEMA_signal_10687), .Q (new_AGEMA_signal_10688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2866 ( .C (clk), .D (new_AGEMA_signal_10690), .Q (new_AGEMA_signal_10691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2869 ( .C (clk), .D (new_AGEMA_signal_10693), .Q (new_AGEMA_signal_10694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2872 ( .C (clk), .D (new_AGEMA_signal_10696), .Q (new_AGEMA_signal_10697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2875 ( .C (clk), .D (new_AGEMA_signal_10699), .Q (new_AGEMA_signal_10700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2878 ( .C (clk), .D (new_AGEMA_signal_10702), .Q (new_AGEMA_signal_10703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2881 ( .C (clk), .D (new_AGEMA_signal_10705), .Q (new_AGEMA_signal_10706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2884 ( .C (clk), .D (new_AGEMA_signal_10708), .Q (new_AGEMA_signal_10709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2887 ( .C (clk), .D (new_AGEMA_signal_10711), .Q (new_AGEMA_signal_10712) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2890 ( .C (clk), .D (new_AGEMA_signal_10714), .Q (new_AGEMA_signal_10715) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2893 ( .C (clk), .D (new_AGEMA_signal_10717), .Q (new_AGEMA_signal_10718) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2896 ( .C (clk), .D (new_AGEMA_signal_10720), .Q (new_AGEMA_signal_10721) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2899 ( .C (clk), .D (new_AGEMA_signal_10723), .Q (new_AGEMA_signal_10724) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2902 ( .C (clk), .D (new_AGEMA_signal_10726), .Q (new_AGEMA_signal_10727) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2905 ( .C (clk), .D (new_AGEMA_signal_10729), .Q (new_AGEMA_signal_10730) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2908 ( .C (clk), .D (new_AGEMA_signal_10732), .Q (new_AGEMA_signal_10733) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2911 ( .C (clk), .D (new_AGEMA_signal_10735), .Q (new_AGEMA_signal_10736) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2914 ( .C (clk), .D (new_AGEMA_signal_10738), .Q (new_AGEMA_signal_10739) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2917 ( .C (clk), .D (new_AGEMA_signal_10741), .Q (new_AGEMA_signal_10742) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2920 ( .C (clk), .D (new_AGEMA_signal_10744), .Q (new_AGEMA_signal_10745) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2923 ( .C (clk), .D (new_AGEMA_signal_10747), .Q (new_AGEMA_signal_10748) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2926 ( .C (clk), .D (new_AGEMA_signal_10750), .Q (new_AGEMA_signal_10751) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2929 ( .C (clk), .D (new_AGEMA_signal_10753), .Q (new_AGEMA_signal_10754) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2932 ( .C (clk), .D (new_AGEMA_signal_10756), .Q (new_AGEMA_signal_10757) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2935 ( .C (clk), .D (new_AGEMA_signal_10759), .Q (new_AGEMA_signal_10760) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2938 ( .C (clk), .D (new_AGEMA_signal_10762), .Q (new_AGEMA_signal_10763) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2941 ( .C (clk), .D (new_AGEMA_signal_10765), .Q (new_AGEMA_signal_10766) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2944 ( .C (clk), .D (new_AGEMA_signal_10768), .Q (new_AGEMA_signal_10769) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2947 ( .C (clk), .D (new_AGEMA_signal_10771), .Q (new_AGEMA_signal_10772) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2950 ( .C (clk), .D (new_AGEMA_signal_10774), .Q (new_AGEMA_signal_10775) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2953 ( .C (clk), .D (new_AGEMA_signal_10777), .Q (new_AGEMA_signal_10778) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2956 ( .C (clk), .D (new_AGEMA_signal_10780), .Q (new_AGEMA_signal_10781) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2959 ( .C (clk), .D (new_AGEMA_signal_10783), .Q (new_AGEMA_signal_10784) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2962 ( .C (clk), .D (new_AGEMA_signal_10786), .Q (new_AGEMA_signal_10787) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2965 ( .C (clk), .D (new_AGEMA_signal_10789), .Q (new_AGEMA_signal_10790) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2968 ( .C (clk), .D (new_AGEMA_signal_10792), .Q (new_AGEMA_signal_10793) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2971 ( .C (clk), .D (new_AGEMA_signal_10795), .Q (new_AGEMA_signal_10796) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2974 ( .C (clk), .D (new_AGEMA_signal_10798), .Q (new_AGEMA_signal_10799) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2977 ( .C (clk), .D (new_AGEMA_signal_10801), .Q (new_AGEMA_signal_10802) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2980 ( .C (clk), .D (new_AGEMA_signal_10804), .Q (new_AGEMA_signal_10805) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2983 ( .C (clk), .D (new_AGEMA_signal_10807), .Q (new_AGEMA_signal_10808) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2986 ( .C (clk), .D (new_AGEMA_signal_10810), .Q (new_AGEMA_signal_10811) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2989 ( .C (clk), .D (new_AGEMA_signal_10813), .Q (new_AGEMA_signal_10814) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2992 ( .C (clk), .D (new_AGEMA_signal_10816), .Q (new_AGEMA_signal_10817) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2995 ( .C (clk), .D (new_AGEMA_signal_10819), .Q (new_AGEMA_signal_10820) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2998 ( .C (clk), .D (new_AGEMA_signal_10822), .Q (new_AGEMA_signal_10823) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3001 ( .C (clk), .D (new_AGEMA_signal_10825), .Q (new_AGEMA_signal_10826) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3004 ( .C (clk), .D (new_AGEMA_signal_10828), .Q (new_AGEMA_signal_10829) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3007 ( .C (clk), .D (new_AGEMA_signal_10831), .Q (new_AGEMA_signal_10832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3010 ( .C (clk), .D (new_AGEMA_signal_10834), .Q (new_AGEMA_signal_10835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3013 ( .C (clk), .D (new_AGEMA_signal_10837), .Q (new_AGEMA_signal_10838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3016 ( .C (clk), .D (new_AGEMA_signal_10840), .Q (new_AGEMA_signal_10841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3019 ( .C (clk), .D (new_AGEMA_signal_10843), .Q (new_AGEMA_signal_10844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3022 ( .C (clk), .D (new_AGEMA_signal_10846), .Q (new_AGEMA_signal_10847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3025 ( .C (clk), .D (new_AGEMA_signal_10849), .Q (new_AGEMA_signal_10850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3028 ( .C (clk), .D (new_AGEMA_signal_10852), .Q (new_AGEMA_signal_10853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3031 ( .C (clk), .D (new_AGEMA_signal_10855), .Q (new_AGEMA_signal_10856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3034 ( .C (clk), .D (new_AGEMA_signal_10858), .Q (new_AGEMA_signal_10859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3037 ( .C (clk), .D (new_AGEMA_signal_10861), .Q (new_AGEMA_signal_10862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3040 ( .C (clk), .D (new_AGEMA_signal_10864), .Q (new_AGEMA_signal_10865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3043 ( .C (clk), .D (new_AGEMA_signal_10867), .Q (new_AGEMA_signal_10868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3046 ( .C (clk), .D (new_AGEMA_signal_10870), .Q (new_AGEMA_signal_10871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3049 ( .C (clk), .D (new_AGEMA_signal_10873), .Q (new_AGEMA_signal_10874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3052 ( .C (clk), .D (new_AGEMA_signal_10876), .Q (new_AGEMA_signal_10877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3055 ( .C (clk), .D (new_AGEMA_signal_10879), .Q (new_AGEMA_signal_10880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3058 ( .C (clk), .D (new_AGEMA_signal_10882), .Q (new_AGEMA_signal_10883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3061 ( .C (clk), .D (new_AGEMA_signal_10885), .Q (new_AGEMA_signal_10886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3064 ( .C (clk), .D (new_AGEMA_signal_10888), .Q (new_AGEMA_signal_10889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3067 ( .C (clk), .D (new_AGEMA_signal_10891), .Q (new_AGEMA_signal_10892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3070 ( .C (clk), .D (new_AGEMA_signal_10894), .Q (new_AGEMA_signal_10895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3073 ( .C (clk), .D (new_AGEMA_signal_10897), .Q (new_AGEMA_signal_10898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3076 ( .C (clk), .D (new_AGEMA_signal_10900), .Q (new_AGEMA_signal_10901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3079 ( .C (clk), .D (new_AGEMA_signal_10903), .Q (new_AGEMA_signal_10904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3082 ( .C (clk), .D (new_AGEMA_signal_10906), .Q (new_AGEMA_signal_10907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3085 ( .C (clk), .D (new_AGEMA_signal_10909), .Q (new_AGEMA_signal_10910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3088 ( .C (clk), .D (new_AGEMA_signal_10912), .Q (new_AGEMA_signal_10913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3091 ( .C (clk), .D (new_AGEMA_signal_10915), .Q (new_AGEMA_signal_10916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3094 ( .C (clk), .D (new_AGEMA_signal_10918), .Q (new_AGEMA_signal_10919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3097 ( .C (clk), .D (new_AGEMA_signal_10921), .Q (new_AGEMA_signal_10922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3100 ( .C (clk), .D (new_AGEMA_signal_10924), .Q (new_AGEMA_signal_10925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3103 ( .C (clk), .D (new_AGEMA_signal_10927), .Q (new_AGEMA_signal_10928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3106 ( .C (clk), .D (new_AGEMA_signal_10930), .Q (new_AGEMA_signal_10931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3109 ( .C (clk), .D (new_AGEMA_signal_10933), .Q (new_AGEMA_signal_10934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3112 ( .C (clk), .D (new_AGEMA_signal_10936), .Q (new_AGEMA_signal_10937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3115 ( .C (clk), .D (new_AGEMA_signal_10939), .Q (new_AGEMA_signal_10940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3118 ( .C (clk), .D (new_AGEMA_signal_10942), .Q (new_AGEMA_signal_10943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3121 ( .C (clk), .D (new_AGEMA_signal_10945), .Q (new_AGEMA_signal_10946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3124 ( .C (clk), .D (new_AGEMA_signal_10948), .Q (new_AGEMA_signal_10949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3127 ( .C (clk), .D (new_AGEMA_signal_10951), .Q (new_AGEMA_signal_10952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3130 ( .C (clk), .D (new_AGEMA_signal_10954), .Q (new_AGEMA_signal_10955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3133 ( .C (clk), .D (new_AGEMA_signal_10957), .Q (new_AGEMA_signal_10958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3136 ( .C (clk), .D (new_AGEMA_signal_10960), .Q (new_AGEMA_signal_10961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3139 ( .C (clk), .D (new_AGEMA_signal_10963), .Q (new_AGEMA_signal_10964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3142 ( .C (clk), .D (new_AGEMA_signal_10966), .Q (new_AGEMA_signal_10967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3145 ( .C (clk), .D (new_AGEMA_signal_10969), .Q (new_AGEMA_signal_10970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3148 ( .C (clk), .D (new_AGEMA_signal_10972), .Q (new_AGEMA_signal_10973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3151 ( .C (clk), .D (new_AGEMA_signal_10975), .Q (new_AGEMA_signal_10976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3154 ( .C (clk), .D (new_AGEMA_signal_10978), .Q (new_AGEMA_signal_10979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3157 ( .C (clk), .D (new_AGEMA_signal_10981), .Q (new_AGEMA_signal_10982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3160 ( .C (clk), .D (new_AGEMA_signal_10984), .Q (new_AGEMA_signal_10985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3163 ( .C (clk), .D (new_AGEMA_signal_10987), .Q (new_AGEMA_signal_10988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3166 ( .C (clk), .D (new_AGEMA_signal_10990), .Q (new_AGEMA_signal_10991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3169 ( .C (clk), .D (new_AGEMA_signal_10993), .Q (new_AGEMA_signal_10994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3172 ( .C (clk), .D (new_AGEMA_signal_10996), .Q (new_AGEMA_signal_10997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3175 ( .C (clk), .D (new_AGEMA_signal_10999), .Q (new_AGEMA_signal_11000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3178 ( .C (clk), .D (new_AGEMA_signal_11002), .Q (new_AGEMA_signal_11003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3181 ( .C (clk), .D (new_AGEMA_signal_11005), .Q (new_AGEMA_signal_11006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3184 ( .C (clk), .D (new_AGEMA_signal_11008), .Q (new_AGEMA_signal_11009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3187 ( .C (clk), .D (new_AGEMA_signal_11011), .Q (new_AGEMA_signal_11012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3190 ( .C (clk), .D (new_AGEMA_signal_11014), .Q (new_AGEMA_signal_11015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3193 ( .C (clk), .D (new_AGEMA_signal_11017), .Q (new_AGEMA_signal_11018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3196 ( .C (clk), .D (new_AGEMA_signal_11020), .Q (new_AGEMA_signal_11021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3199 ( .C (clk), .D (new_AGEMA_signal_11023), .Q (new_AGEMA_signal_11024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3202 ( .C (clk), .D (new_AGEMA_signal_11026), .Q (new_AGEMA_signal_11027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3205 ( .C (clk), .D (new_AGEMA_signal_11029), .Q (new_AGEMA_signal_11030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3208 ( .C (clk), .D (new_AGEMA_signal_11032), .Q (new_AGEMA_signal_11033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3211 ( .C (clk), .D (new_AGEMA_signal_11035), .Q (new_AGEMA_signal_11036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3214 ( .C (clk), .D (new_AGEMA_signal_11038), .Q (new_AGEMA_signal_11039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3217 ( .C (clk), .D (new_AGEMA_signal_11041), .Q (new_AGEMA_signal_11042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3220 ( .C (clk), .D (new_AGEMA_signal_11044), .Q (new_AGEMA_signal_11045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3223 ( .C (clk), .D (new_AGEMA_signal_11047), .Q (new_AGEMA_signal_11048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3226 ( .C (clk), .D (new_AGEMA_signal_11050), .Q (new_AGEMA_signal_11051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3229 ( .C (clk), .D (new_AGEMA_signal_11053), .Q (new_AGEMA_signal_11054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3232 ( .C (clk), .D (new_AGEMA_signal_11056), .Q (new_AGEMA_signal_11057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3235 ( .C (clk), .D (new_AGEMA_signal_11059), .Q (new_AGEMA_signal_11060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3238 ( .C (clk), .D (new_AGEMA_signal_11062), .Q (new_AGEMA_signal_11063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3241 ( .C (clk), .D (new_AGEMA_signal_11065), .Q (new_AGEMA_signal_11066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3244 ( .C (clk), .D (new_AGEMA_signal_11068), .Q (new_AGEMA_signal_11069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3247 ( .C (clk), .D (new_AGEMA_signal_11071), .Q (new_AGEMA_signal_11072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3250 ( .C (clk), .D (new_AGEMA_signal_11074), .Q (new_AGEMA_signal_11075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3253 ( .C (clk), .D (new_AGEMA_signal_11077), .Q (new_AGEMA_signal_11078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3256 ( .C (clk), .D (new_AGEMA_signal_11080), .Q (new_AGEMA_signal_11081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3259 ( .C (clk), .D (new_AGEMA_signal_11083), .Q (new_AGEMA_signal_11084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3262 ( .C (clk), .D (new_AGEMA_signal_11086), .Q (new_AGEMA_signal_11087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3265 ( .C (clk), .D (new_AGEMA_signal_11089), .Q (new_AGEMA_signal_11090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3268 ( .C (clk), .D (new_AGEMA_signal_11092), .Q (new_AGEMA_signal_11093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3271 ( .C (clk), .D (new_AGEMA_signal_11095), .Q (new_AGEMA_signal_11096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3274 ( .C (clk), .D (new_AGEMA_signal_11098), .Q (new_AGEMA_signal_11099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3277 ( .C (clk), .D (new_AGEMA_signal_11101), .Q (new_AGEMA_signal_11102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3280 ( .C (clk), .D (new_AGEMA_signal_11104), .Q (new_AGEMA_signal_11105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3283 ( .C (clk), .D (new_AGEMA_signal_11107), .Q (new_AGEMA_signal_11108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3286 ( .C (clk), .D (new_AGEMA_signal_11110), .Q (new_AGEMA_signal_11111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3289 ( .C (clk), .D (new_AGEMA_signal_11113), .Q (new_AGEMA_signal_11114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3292 ( .C (clk), .D (new_AGEMA_signal_11116), .Q (new_AGEMA_signal_11117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3295 ( .C (clk), .D (new_AGEMA_signal_11119), .Q (new_AGEMA_signal_11120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3298 ( .C (clk), .D (new_AGEMA_signal_11122), .Q (new_AGEMA_signal_11123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3301 ( .C (clk), .D (new_AGEMA_signal_11125), .Q (new_AGEMA_signal_11126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3304 ( .C (clk), .D (new_AGEMA_signal_11128), .Q (new_AGEMA_signal_11129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3307 ( .C (clk), .D (new_AGEMA_signal_11131), .Q (new_AGEMA_signal_11132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3310 ( .C (clk), .D (new_AGEMA_signal_11134), .Q (new_AGEMA_signal_11135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3313 ( .C (clk), .D (new_AGEMA_signal_11137), .Q (new_AGEMA_signal_11138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3316 ( .C (clk), .D (new_AGEMA_signal_11140), .Q (new_AGEMA_signal_11141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3319 ( .C (clk), .D (new_AGEMA_signal_11143), .Q (new_AGEMA_signal_11144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3322 ( .C (clk), .D (new_AGEMA_signal_11146), .Q (new_AGEMA_signal_11147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3325 ( .C (clk), .D (new_AGEMA_signal_11149), .Q (new_AGEMA_signal_11150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3328 ( .C (clk), .D (new_AGEMA_signal_11152), .Q (new_AGEMA_signal_11153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3331 ( .C (clk), .D (new_AGEMA_signal_11155), .Q (new_AGEMA_signal_11156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3334 ( .C (clk), .D (new_AGEMA_signal_11158), .Q (new_AGEMA_signal_11159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3337 ( .C (clk), .D (new_AGEMA_signal_11161), .Q (new_AGEMA_signal_11162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3340 ( .C (clk), .D (new_AGEMA_signal_11164), .Q (new_AGEMA_signal_11165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3343 ( .C (clk), .D (new_AGEMA_signal_11167), .Q (new_AGEMA_signal_11168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3346 ( .C (clk), .D (new_AGEMA_signal_11170), .Q (new_AGEMA_signal_11171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3349 ( .C (clk), .D (new_AGEMA_signal_11173), .Q (new_AGEMA_signal_11174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3352 ( .C (clk), .D (new_AGEMA_signal_11176), .Q (new_AGEMA_signal_11177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3355 ( .C (clk), .D (new_AGEMA_signal_11179), .Q (new_AGEMA_signal_11180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3358 ( .C (clk), .D (new_AGEMA_signal_11182), .Q (new_AGEMA_signal_11183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3361 ( .C (clk), .D (new_AGEMA_signal_11185), .Q (new_AGEMA_signal_11186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3364 ( .C (clk), .D (new_AGEMA_signal_11188), .Q (new_AGEMA_signal_11189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3367 ( .C (clk), .D (new_AGEMA_signal_11191), .Q (new_AGEMA_signal_11192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3370 ( .C (clk), .D (new_AGEMA_signal_11194), .Q (new_AGEMA_signal_11195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3373 ( .C (clk), .D (new_AGEMA_signal_11197), .Q (new_AGEMA_signal_11198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3376 ( .C (clk), .D (new_AGEMA_signal_11200), .Q (new_AGEMA_signal_11201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3379 ( .C (clk), .D (new_AGEMA_signal_11203), .Q (new_AGEMA_signal_11204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3382 ( .C (clk), .D (new_AGEMA_signal_11206), .Q (new_AGEMA_signal_11207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3385 ( .C (clk), .D (new_AGEMA_signal_11209), .Q (new_AGEMA_signal_11210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3388 ( .C (clk), .D (new_AGEMA_signal_11212), .Q (new_AGEMA_signal_11213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3391 ( .C (clk), .D (new_AGEMA_signal_11215), .Q (new_AGEMA_signal_11216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3394 ( .C (clk), .D (new_AGEMA_signal_11218), .Q (new_AGEMA_signal_11219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3397 ( .C (clk), .D (new_AGEMA_signal_11221), .Q (new_AGEMA_signal_11222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3400 ( .C (clk), .D (new_AGEMA_signal_11224), .Q (new_AGEMA_signal_11225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3403 ( .C (clk), .D (new_AGEMA_signal_11227), .Q (new_AGEMA_signal_11228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3406 ( .C (clk), .D (new_AGEMA_signal_11230), .Q (new_AGEMA_signal_11231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3409 ( .C (clk), .D (new_AGEMA_signal_11233), .Q (new_AGEMA_signal_11234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3412 ( .C (clk), .D (new_AGEMA_signal_11236), .Q (new_AGEMA_signal_11237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3415 ( .C (clk), .D (new_AGEMA_signal_11239), .Q (new_AGEMA_signal_11240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3418 ( .C (clk), .D (new_AGEMA_signal_11242), .Q (new_AGEMA_signal_11243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3421 ( .C (clk), .D (new_AGEMA_signal_11245), .Q (new_AGEMA_signal_11246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3424 ( .C (clk), .D (new_AGEMA_signal_11248), .Q (new_AGEMA_signal_11249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3427 ( .C (clk), .D (new_AGEMA_signal_11251), .Q (new_AGEMA_signal_11252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3430 ( .C (clk), .D (new_AGEMA_signal_11254), .Q (new_AGEMA_signal_11255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3433 ( .C (clk), .D (new_AGEMA_signal_11257), .Q (new_AGEMA_signal_11258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3436 ( .C (clk), .D (new_AGEMA_signal_11260), .Q (new_AGEMA_signal_11261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3439 ( .C (clk), .D (new_AGEMA_signal_11263), .Q (new_AGEMA_signal_11264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3442 ( .C (clk), .D (new_AGEMA_signal_11266), .Q (new_AGEMA_signal_11267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3445 ( .C (clk), .D (new_AGEMA_signal_11269), .Q (new_AGEMA_signal_11270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3448 ( .C (clk), .D (new_AGEMA_signal_11272), .Q (new_AGEMA_signal_11273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3451 ( .C (clk), .D (new_AGEMA_signal_11275), .Q (new_AGEMA_signal_11276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3454 ( .C (clk), .D (new_AGEMA_signal_11278), .Q (new_AGEMA_signal_11279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3457 ( .C (clk), .D (new_AGEMA_signal_11281), .Q (new_AGEMA_signal_11282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3460 ( .C (clk), .D (new_AGEMA_signal_11284), .Q (new_AGEMA_signal_11285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3463 ( .C (clk), .D (new_AGEMA_signal_11287), .Q (new_AGEMA_signal_11288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3466 ( .C (clk), .D (new_AGEMA_signal_11290), .Q (new_AGEMA_signal_11291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3469 ( .C (clk), .D (new_AGEMA_signal_11293), .Q (new_AGEMA_signal_11294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3472 ( .C (clk), .D (new_AGEMA_signal_11296), .Q (new_AGEMA_signal_11297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3475 ( .C (clk), .D (new_AGEMA_signal_11299), .Q (new_AGEMA_signal_11300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3478 ( .C (clk), .D (new_AGEMA_signal_11302), .Q (new_AGEMA_signal_11303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3481 ( .C (clk), .D (new_AGEMA_signal_11305), .Q (new_AGEMA_signal_11306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3484 ( .C (clk), .D (new_AGEMA_signal_11308), .Q (new_AGEMA_signal_11309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3487 ( .C (clk), .D (new_AGEMA_signal_11311), .Q (new_AGEMA_signal_11312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3490 ( .C (clk), .D (new_AGEMA_signal_11314), .Q (new_AGEMA_signal_11315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3493 ( .C (clk), .D (new_AGEMA_signal_11317), .Q (new_AGEMA_signal_11318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3496 ( .C (clk), .D (new_AGEMA_signal_11320), .Q (new_AGEMA_signal_11321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3499 ( .C (clk), .D (new_AGEMA_signal_11323), .Q (new_AGEMA_signal_11324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3502 ( .C (clk), .D (new_AGEMA_signal_11326), .Q (new_AGEMA_signal_11327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3505 ( .C (clk), .D (new_AGEMA_signal_11329), .Q (new_AGEMA_signal_11330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3508 ( .C (clk), .D (new_AGEMA_signal_11332), .Q (new_AGEMA_signal_11333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3511 ( .C (clk), .D (new_AGEMA_signal_11335), .Q (new_AGEMA_signal_11336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3514 ( .C (clk), .D (new_AGEMA_signal_11338), .Q (new_AGEMA_signal_11339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3517 ( .C (clk), .D (new_AGEMA_signal_11341), .Q (new_AGEMA_signal_11342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3520 ( .C (clk), .D (new_AGEMA_signal_11344), .Q (new_AGEMA_signal_11345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3523 ( .C (clk), .D (new_AGEMA_signal_11347), .Q (new_AGEMA_signal_11348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3526 ( .C (clk), .D (new_AGEMA_signal_11350), .Q (new_AGEMA_signal_11351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3529 ( .C (clk), .D (new_AGEMA_signal_11353), .Q (new_AGEMA_signal_11354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3532 ( .C (clk), .D (new_AGEMA_signal_11356), .Q (new_AGEMA_signal_11357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3535 ( .C (clk), .D (new_AGEMA_signal_11359), .Q (new_AGEMA_signal_11360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3538 ( .C (clk), .D (new_AGEMA_signal_11362), .Q (new_AGEMA_signal_11363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3541 ( .C (clk), .D (new_AGEMA_signal_11365), .Q (new_AGEMA_signal_11366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3544 ( .C (clk), .D (new_AGEMA_signal_11368), .Q (new_AGEMA_signal_11369) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3547 ( .C (clk), .D (new_AGEMA_signal_11371), .Q (new_AGEMA_signal_11372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3550 ( .C (clk), .D (new_AGEMA_signal_11374), .Q (new_AGEMA_signal_11375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3553 ( .C (clk), .D (new_AGEMA_signal_11377), .Q (new_AGEMA_signal_11378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3556 ( .C (clk), .D (new_AGEMA_signal_11380), .Q (new_AGEMA_signal_11381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3559 ( .C (clk), .D (new_AGEMA_signal_11383), .Q (new_AGEMA_signal_11384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3562 ( .C (clk), .D (new_AGEMA_signal_11386), .Q (new_AGEMA_signal_11387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3565 ( .C (clk), .D (new_AGEMA_signal_11389), .Q (new_AGEMA_signal_11390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3568 ( .C (clk), .D (new_AGEMA_signal_11392), .Q (new_AGEMA_signal_11393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3571 ( .C (clk), .D (new_AGEMA_signal_11395), .Q (new_AGEMA_signal_11396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3574 ( .C (clk), .D (new_AGEMA_signal_11398), .Q (new_AGEMA_signal_11399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3577 ( .C (clk), .D (new_AGEMA_signal_11401), .Q (new_AGEMA_signal_11402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3580 ( .C (clk), .D (new_AGEMA_signal_11404), .Q (new_AGEMA_signal_11405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3583 ( .C (clk), .D (new_AGEMA_signal_11407), .Q (new_AGEMA_signal_11408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3586 ( .C (clk), .D (new_AGEMA_signal_11410), .Q (new_AGEMA_signal_11411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3589 ( .C (clk), .D (new_AGEMA_signal_11413), .Q (new_AGEMA_signal_11414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3592 ( .C (clk), .D (new_AGEMA_signal_11416), .Q (new_AGEMA_signal_11417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3595 ( .C (clk), .D (new_AGEMA_signal_11419), .Q (new_AGEMA_signal_11420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3598 ( .C (clk), .D (new_AGEMA_signal_11422), .Q (new_AGEMA_signal_11423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3601 ( .C (clk), .D (new_AGEMA_signal_11425), .Q (new_AGEMA_signal_11426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3604 ( .C (clk), .D (new_AGEMA_signal_11428), .Q (new_AGEMA_signal_11429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3607 ( .C (clk), .D (new_AGEMA_signal_11431), .Q (new_AGEMA_signal_11432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3610 ( .C (clk), .D (new_AGEMA_signal_11434), .Q (new_AGEMA_signal_11435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3613 ( .C (clk), .D (new_AGEMA_signal_11437), .Q (new_AGEMA_signal_11438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3616 ( .C (clk), .D (new_AGEMA_signal_11440), .Q (new_AGEMA_signal_11441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3619 ( .C (clk), .D (new_AGEMA_signal_11443), .Q (new_AGEMA_signal_11444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3622 ( .C (clk), .D (new_AGEMA_signal_11446), .Q (new_AGEMA_signal_11447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3625 ( .C (clk), .D (new_AGEMA_signal_11449), .Q (new_AGEMA_signal_11450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3628 ( .C (clk), .D (new_AGEMA_signal_11452), .Q (new_AGEMA_signal_11453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3631 ( .C (clk), .D (new_AGEMA_signal_11455), .Q (new_AGEMA_signal_11456) ) ;
    buf_clk new_AGEMA_reg_buffer_3634 ( .C (clk), .D (new_AGEMA_signal_11458), .Q (new_AGEMA_signal_11459) ) ;
    buf_clk new_AGEMA_reg_buffer_3638 ( .C (clk), .D (new_AGEMA_signal_11462), .Q (new_AGEMA_signal_11463) ) ;
    buf_clk new_AGEMA_reg_buffer_3642 ( .C (clk), .D (new_AGEMA_signal_11466), .Q (new_AGEMA_signal_11467) ) ;
    buf_clk new_AGEMA_reg_buffer_3646 ( .C (clk), .D (new_AGEMA_signal_11470), .Q (new_AGEMA_signal_11471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3650 ( .C (clk), .D (new_AGEMA_signal_11474), .Q (new_AGEMA_signal_11475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3654 ( .C (clk), .D (new_AGEMA_signal_11478), .Q (new_AGEMA_signal_11479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3658 ( .C (clk), .D (new_AGEMA_signal_11482), .Q (new_AGEMA_signal_11483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3662 ( .C (clk), .D (new_AGEMA_signal_11486), .Q (new_AGEMA_signal_11487) ) ;
    buf_clk new_AGEMA_reg_buffer_3666 ( .C (clk), .D (new_AGEMA_signal_11490), .Q (new_AGEMA_signal_11491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3670 ( .C (clk), .D (new_AGEMA_signal_11494), .Q (new_AGEMA_signal_11495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3674 ( .C (clk), .D (new_AGEMA_signal_11498), .Q (new_AGEMA_signal_11499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3678 ( .C (clk), .D (new_AGEMA_signal_11502), .Q (new_AGEMA_signal_11503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3682 ( .C (clk), .D (new_AGEMA_signal_11506), .Q (new_AGEMA_signal_11507) ) ;
    buf_clk new_AGEMA_reg_buffer_3686 ( .C (clk), .D (new_AGEMA_signal_11510), .Q (new_AGEMA_signal_11511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3690 ( .C (clk), .D (new_AGEMA_signal_11514), .Q (new_AGEMA_signal_11515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3694 ( .C (clk), .D (new_AGEMA_signal_11518), .Q (new_AGEMA_signal_11519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3698 ( .C (clk), .D (new_AGEMA_signal_11522), .Q (new_AGEMA_signal_11523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3702 ( .C (clk), .D (new_AGEMA_signal_11526), .Q (new_AGEMA_signal_11527) ) ;
    buf_clk new_AGEMA_reg_buffer_3706 ( .C (clk), .D (new_AGEMA_signal_11530), .Q (new_AGEMA_signal_11531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3710 ( .C (clk), .D (new_AGEMA_signal_11534), .Q (new_AGEMA_signal_11535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3714 ( .C (clk), .D (new_AGEMA_signal_11538), .Q (new_AGEMA_signal_11539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3718 ( .C (clk), .D (new_AGEMA_signal_11542), .Q (new_AGEMA_signal_11543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3722 ( .C (clk), .D (new_AGEMA_signal_11546), .Q (new_AGEMA_signal_11547) ) ;
    buf_clk new_AGEMA_reg_buffer_3726 ( .C (clk), .D (new_AGEMA_signal_11550), .Q (new_AGEMA_signal_11551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3730 ( .C (clk), .D (new_AGEMA_signal_11554), .Q (new_AGEMA_signal_11555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3734 ( .C (clk), .D (new_AGEMA_signal_11558), .Q (new_AGEMA_signal_11559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3738 ( .C (clk), .D (new_AGEMA_signal_11562), .Q (new_AGEMA_signal_11563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3742 ( .C (clk), .D (new_AGEMA_signal_11566), .Q (new_AGEMA_signal_11567) ) ;
    buf_clk new_AGEMA_reg_buffer_3746 ( .C (clk), .D (new_AGEMA_signal_11570), .Q (new_AGEMA_signal_11571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3750 ( .C (clk), .D (new_AGEMA_signal_11574), .Q (new_AGEMA_signal_11575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3754 ( .C (clk), .D (new_AGEMA_signal_11578), .Q (new_AGEMA_signal_11579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3758 ( .C (clk), .D (new_AGEMA_signal_11582), .Q (new_AGEMA_signal_11583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3762 ( .C (clk), .D (new_AGEMA_signal_11586), .Q (new_AGEMA_signal_11587) ) ;
    buf_clk new_AGEMA_reg_buffer_3766 ( .C (clk), .D (new_AGEMA_signal_11590), .Q (new_AGEMA_signal_11591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3770 ( .C (clk), .D (new_AGEMA_signal_11594), .Q (new_AGEMA_signal_11595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3774 ( .C (clk), .D (new_AGEMA_signal_11598), .Q (new_AGEMA_signal_11599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3778 ( .C (clk), .D (new_AGEMA_signal_11602), .Q (new_AGEMA_signal_11603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3782 ( .C (clk), .D (new_AGEMA_signal_11606), .Q (new_AGEMA_signal_11607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3786 ( .C (clk), .D (new_AGEMA_signal_11610), .Q (new_AGEMA_signal_11611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3790 ( .C (clk), .D (new_AGEMA_signal_11614), .Q (new_AGEMA_signal_11615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3794 ( .C (clk), .D (new_AGEMA_signal_11618), .Q (new_AGEMA_signal_11619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3798 ( .C (clk), .D (new_AGEMA_signal_11622), .Q (new_AGEMA_signal_11623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3802 ( .C (clk), .D (new_AGEMA_signal_11626), .Q (new_AGEMA_signal_11627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3806 ( .C (clk), .D (new_AGEMA_signal_11630), .Q (new_AGEMA_signal_11631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3810 ( .C (clk), .D (new_AGEMA_signal_11634), .Q (new_AGEMA_signal_11635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3814 ( .C (clk), .D (new_AGEMA_signal_11638), .Q (new_AGEMA_signal_11639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3818 ( .C (clk), .D (new_AGEMA_signal_11642), .Q (new_AGEMA_signal_11643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3822 ( .C (clk), .D (new_AGEMA_signal_11646), .Q (new_AGEMA_signal_11647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3826 ( .C (clk), .D (new_AGEMA_signal_11650), .Q (new_AGEMA_signal_11651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3830 ( .C (clk), .D (new_AGEMA_signal_11654), .Q (new_AGEMA_signal_11655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3834 ( .C (clk), .D (new_AGEMA_signal_11658), .Q (new_AGEMA_signal_11659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3838 ( .C (clk), .D (new_AGEMA_signal_11662), .Q (new_AGEMA_signal_11663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3842 ( .C (clk), .D (new_AGEMA_signal_11666), .Q (new_AGEMA_signal_11667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3846 ( .C (clk), .D (new_AGEMA_signal_11670), .Q (new_AGEMA_signal_11671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3850 ( .C (clk), .D (new_AGEMA_signal_11674), .Q (new_AGEMA_signal_11675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3854 ( .C (clk), .D (new_AGEMA_signal_11678), .Q (new_AGEMA_signal_11679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3858 ( .C (clk), .D (new_AGEMA_signal_11682), .Q (new_AGEMA_signal_11683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3862 ( .C (clk), .D (new_AGEMA_signal_11686), .Q (new_AGEMA_signal_11687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3866 ( .C (clk), .D (new_AGEMA_signal_11690), .Q (new_AGEMA_signal_11691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3870 ( .C (clk), .D (new_AGEMA_signal_11694), .Q (new_AGEMA_signal_11695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3874 ( .C (clk), .D (new_AGEMA_signal_11698), .Q (new_AGEMA_signal_11699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3878 ( .C (clk), .D (new_AGEMA_signal_11702), .Q (new_AGEMA_signal_11703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3882 ( .C (clk), .D (new_AGEMA_signal_11706), .Q (new_AGEMA_signal_11707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3886 ( .C (clk), .D (new_AGEMA_signal_11710), .Q (new_AGEMA_signal_11711) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3890 ( .C (clk), .D (new_AGEMA_signal_11714), .Q (new_AGEMA_signal_11715) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3894 ( .C (clk), .D (new_AGEMA_signal_11718), .Q (new_AGEMA_signal_11719) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3898 ( .C (clk), .D (new_AGEMA_signal_11722), .Q (new_AGEMA_signal_11723) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3902 ( .C (clk), .D (new_AGEMA_signal_11726), .Q (new_AGEMA_signal_11727) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3906 ( .C (clk), .D (new_AGEMA_signal_11730), .Q (new_AGEMA_signal_11731) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3910 ( .C (clk), .D (new_AGEMA_signal_11734), .Q (new_AGEMA_signal_11735) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3914 ( .C (clk), .D (new_AGEMA_signal_11738), .Q (new_AGEMA_signal_11739) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3918 ( .C (clk), .D (new_AGEMA_signal_11742), .Q (new_AGEMA_signal_11743) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3922 ( .C (clk), .D (new_AGEMA_signal_11746), .Q (new_AGEMA_signal_11747) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3926 ( .C (clk), .D (new_AGEMA_signal_11750), .Q (new_AGEMA_signal_11751) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3930 ( .C (clk), .D (new_AGEMA_signal_11754), .Q (new_AGEMA_signal_11755) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3934 ( .C (clk), .D (new_AGEMA_signal_11758), .Q (new_AGEMA_signal_11759) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3938 ( .C (clk), .D (new_AGEMA_signal_11762), .Q (new_AGEMA_signal_11763) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3942 ( .C (clk), .D (new_AGEMA_signal_11766), .Q (new_AGEMA_signal_11767) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3946 ( .C (clk), .D (new_AGEMA_signal_11770), .Q (new_AGEMA_signal_11771) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3950 ( .C (clk), .D (new_AGEMA_signal_11774), .Q (new_AGEMA_signal_11775) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3954 ( .C (clk), .D (new_AGEMA_signal_11778), .Q (new_AGEMA_signal_11779) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3958 ( .C (clk), .D (new_AGEMA_signal_11782), .Q (new_AGEMA_signal_11783) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3962 ( .C (clk), .D (new_AGEMA_signal_11786), .Q (new_AGEMA_signal_11787) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3966 ( .C (clk), .D (new_AGEMA_signal_11790), .Q (new_AGEMA_signal_11791) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3970 ( .C (clk), .D (new_AGEMA_signal_11794), .Q (new_AGEMA_signal_11795) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3974 ( .C (clk), .D (new_AGEMA_signal_11798), .Q (new_AGEMA_signal_11799) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3978 ( .C (clk), .D (new_AGEMA_signal_11802), .Q (new_AGEMA_signal_11803) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3982 ( .C (clk), .D (new_AGEMA_signal_11806), .Q (new_AGEMA_signal_11807) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3986 ( .C (clk), .D (new_AGEMA_signal_11810), .Q (new_AGEMA_signal_11811) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3990 ( .C (clk), .D (new_AGEMA_signal_11814), .Q (new_AGEMA_signal_11815) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3994 ( .C (clk), .D (new_AGEMA_signal_11818), .Q (new_AGEMA_signal_11819) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3998 ( .C (clk), .D (new_AGEMA_signal_11822), .Q (new_AGEMA_signal_11823) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4002 ( .C (clk), .D (new_AGEMA_signal_11826), .Q (new_AGEMA_signal_11827) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4006 ( .C (clk), .D (new_AGEMA_signal_11830), .Q (new_AGEMA_signal_11831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4010 ( .C (clk), .D (new_AGEMA_signal_11834), .Q (new_AGEMA_signal_11835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4014 ( .C (clk), .D (new_AGEMA_signal_11838), .Q (new_AGEMA_signal_11839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4018 ( .C (clk), .D (new_AGEMA_signal_11842), .Q (new_AGEMA_signal_11843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4022 ( .C (clk), .D (new_AGEMA_signal_11846), .Q (new_AGEMA_signal_11847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4026 ( .C (clk), .D (new_AGEMA_signal_11850), .Q (new_AGEMA_signal_11851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4030 ( .C (clk), .D (new_AGEMA_signal_11854), .Q (new_AGEMA_signal_11855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4034 ( .C (clk), .D (new_AGEMA_signal_11858), .Q (new_AGEMA_signal_11859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4038 ( .C (clk), .D (new_AGEMA_signal_11862), .Q (new_AGEMA_signal_11863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4042 ( .C (clk), .D (new_AGEMA_signal_11866), .Q (new_AGEMA_signal_11867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4046 ( .C (clk), .D (new_AGEMA_signal_11870), .Q (new_AGEMA_signal_11871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4050 ( .C (clk), .D (new_AGEMA_signal_11874), .Q (new_AGEMA_signal_11875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4054 ( .C (clk), .D (new_AGEMA_signal_11878), .Q (new_AGEMA_signal_11879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4058 ( .C (clk), .D (new_AGEMA_signal_11882), .Q (new_AGEMA_signal_11883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4062 ( .C (clk), .D (new_AGEMA_signal_11886), .Q (new_AGEMA_signal_11887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4066 ( .C (clk), .D (new_AGEMA_signal_11890), .Q (new_AGEMA_signal_11891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4070 ( .C (clk), .D (new_AGEMA_signal_11894), .Q (new_AGEMA_signal_11895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4074 ( .C (clk), .D (new_AGEMA_signal_11898), .Q (new_AGEMA_signal_11899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4078 ( .C (clk), .D (new_AGEMA_signal_11902), .Q (new_AGEMA_signal_11903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4082 ( .C (clk), .D (new_AGEMA_signal_11906), .Q (new_AGEMA_signal_11907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4086 ( .C (clk), .D (new_AGEMA_signal_11910), .Q (new_AGEMA_signal_11911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4090 ( .C (clk), .D (new_AGEMA_signal_11914), .Q (new_AGEMA_signal_11915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4094 ( .C (clk), .D (new_AGEMA_signal_11918), .Q (new_AGEMA_signal_11919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4098 ( .C (clk), .D (new_AGEMA_signal_11922), .Q (new_AGEMA_signal_11923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4102 ( .C (clk), .D (new_AGEMA_signal_11926), .Q (new_AGEMA_signal_11927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4106 ( .C (clk), .D (new_AGEMA_signal_11930), .Q (new_AGEMA_signal_11931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4110 ( .C (clk), .D (new_AGEMA_signal_11934), .Q (new_AGEMA_signal_11935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4114 ( .C (clk), .D (new_AGEMA_signal_11938), .Q (new_AGEMA_signal_11939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4118 ( .C (clk), .D (new_AGEMA_signal_11942), .Q (new_AGEMA_signal_11943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4122 ( .C (clk), .D (new_AGEMA_signal_11946), .Q (new_AGEMA_signal_11947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4126 ( .C (clk), .D (new_AGEMA_signal_11950), .Q (new_AGEMA_signal_11951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4130 ( .C (clk), .D (new_AGEMA_signal_11954), .Q (new_AGEMA_signal_11955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4134 ( .C (clk), .D (new_AGEMA_signal_11958), .Q (new_AGEMA_signal_11959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4138 ( .C (clk), .D (new_AGEMA_signal_11962), .Q (new_AGEMA_signal_11963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4142 ( .C (clk), .D (new_AGEMA_signal_11966), .Q (new_AGEMA_signal_11967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4146 ( .C (clk), .D (new_AGEMA_signal_11970), .Q (new_AGEMA_signal_11971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4150 ( .C (clk), .D (new_AGEMA_signal_11974), .Q (new_AGEMA_signal_11975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4154 ( .C (clk), .D (new_AGEMA_signal_11978), .Q (new_AGEMA_signal_11979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4158 ( .C (clk), .D (new_AGEMA_signal_11982), .Q (new_AGEMA_signal_11983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4162 ( .C (clk), .D (new_AGEMA_signal_11986), .Q (new_AGEMA_signal_11987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4166 ( .C (clk), .D (new_AGEMA_signal_11990), .Q (new_AGEMA_signal_11991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4170 ( .C (clk), .D (new_AGEMA_signal_11994), .Q (new_AGEMA_signal_11995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4174 ( .C (clk), .D (new_AGEMA_signal_11998), .Q (new_AGEMA_signal_11999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4178 ( .C (clk), .D (new_AGEMA_signal_12002), .Q (new_AGEMA_signal_12003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4182 ( .C (clk), .D (new_AGEMA_signal_12006), .Q (new_AGEMA_signal_12007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4186 ( .C (clk), .D (new_AGEMA_signal_12010), .Q (new_AGEMA_signal_12011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4190 ( .C (clk), .D (new_AGEMA_signal_12014), .Q (new_AGEMA_signal_12015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4194 ( .C (clk), .D (new_AGEMA_signal_12018), .Q (new_AGEMA_signal_12019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4198 ( .C (clk), .D (new_AGEMA_signal_12022), .Q (new_AGEMA_signal_12023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4202 ( .C (clk), .D (new_AGEMA_signal_12026), .Q (new_AGEMA_signal_12027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4206 ( .C (clk), .D (new_AGEMA_signal_12030), .Q (new_AGEMA_signal_12031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4210 ( .C (clk), .D (new_AGEMA_signal_12034), .Q (new_AGEMA_signal_12035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4214 ( .C (clk), .D (new_AGEMA_signal_12038), .Q (new_AGEMA_signal_12039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4218 ( .C (clk), .D (new_AGEMA_signal_12042), .Q (new_AGEMA_signal_12043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4222 ( .C (clk), .D (new_AGEMA_signal_12046), .Q (new_AGEMA_signal_12047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4226 ( .C (clk), .D (new_AGEMA_signal_12050), .Q (new_AGEMA_signal_12051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4230 ( .C (clk), .D (new_AGEMA_signal_12054), .Q (new_AGEMA_signal_12055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4234 ( .C (clk), .D (new_AGEMA_signal_12058), .Q (new_AGEMA_signal_12059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4238 ( .C (clk), .D (new_AGEMA_signal_12062), .Q (new_AGEMA_signal_12063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4242 ( .C (clk), .D (new_AGEMA_signal_12066), .Q (new_AGEMA_signal_12067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4246 ( .C (clk), .D (new_AGEMA_signal_12070), .Q (new_AGEMA_signal_12071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4250 ( .C (clk), .D (new_AGEMA_signal_12074), .Q (new_AGEMA_signal_12075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4254 ( .C (clk), .D (new_AGEMA_signal_12078), .Q (new_AGEMA_signal_12079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4258 ( .C (clk), .D (new_AGEMA_signal_12082), .Q (new_AGEMA_signal_12083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4262 ( .C (clk), .D (new_AGEMA_signal_12086), .Q (new_AGEMA_signal_12087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4266 ( .C (clk), .D (new_AGEMA_signal_12090), .Q (new_AGEMA_signal_12091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4270 ( .C (clk), .D (new_AGEMA_signal_12094), .Q (new_AGEMA_signal_12095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4274 ( .C (clk), .D (new_AGEMA_signal_12098), .Q (new_AGEMA_signal_12099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4278 ( .C (clk), .D (new_AGEMA_signal_12102), .Q (new_AGEMA_signal_12103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4282 ( .C (clk), .D (new_AGEMA_signal_12106), .Q (new_AGEMA_signal_12107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4286 ( .C (clk), .D (new_AGEMA_signal_12110), .Q (new_AGEMA_signal_12111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4290 ( .C (clk), .D (new_AGEMA_signal_12114), .Q (new_AGEMA_signal_12115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4294 ( .C (clk), .D (new_AGEMA_signal_12118), .Q (new_AGEMA_signal_12119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4298 ( .C (clk), .D (new_AGEMA_signal_12122), .Q (new_AGEMA_signal_12123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4302 ( .C (clk), .D (new_AGEMA_signal_12126), .Q (new_AGEMA_signal_12127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4306 ( .C (clk), .D (new_AGEMA_signal_12130), .Q (new_AGEMA_signal_12131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4310 ( .C (clk), .D (new_AGEMA_signal_12134), .Q (new_AGEMA_signal_12135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4314 ( .C (clk), .D (new_AGEMA_signal_12138), .Q (new_AGEMA_signal_12139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4318 ( .C (clk), .D (new_AGEMA_signal_12142), .Q (new_AGEMA_signal_12143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4322 ( .C (clk), .D (new_AGEMA_signal_12146), .Q (new_AGEMA_signal_12147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4326 ( .C (clk), .D (new_AGEMA_signal_12150), .Q (new_AGEMA_signal_12151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4330 ( .C (clk), .D (new_AGEMA_signal_12154), .Q (new_AGEMA_signal_12155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4334 ( .C (clk), .D (new_AGEMA_signal_12158), .Q (new_AGEMA_signal_12159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4338 ( .C (clk), .D (new_AGEMA_signal_12162), .Q (new_AGEMA_signal_12163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4342 ( .C (clk), .D (new_AGEMA_signal_12166), .Q (new_AGEMA_signal_12167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4346 ( .C (clk), .D (new_AGEMA_signal_12170), .Q (new_AGEMA_signal_12171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4350 ( .C (clk), .D (new_AGEMA_signal_12174), .Q (new_AGEMA_signal_12175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4354 ( .C (clk), .D (new_AGEMA_signal_12178), .Q (new_AGEMA_signal_12179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4358 ( .C (clk), .D (new_AGEMA_signal_12182), .Q (new_AGEMA_signal_12183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4362 ( .C (clk), .D (new_AGEMA_signal_12186), .Q (new_AGEMA_signal_12187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4366 ( .C (clk), .D (new_AGEMA_signal_12190), .Q (new_AGEMA_signal_12191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4370 ( .C (clk), .D (new_AGEMA_signal_12194), .Q (new_AGEMA_signal_12195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4374 ( .C (clk), .D (new_AGEMA_signal_12198), .Q (new_AGEMA_signal_12199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4378 ( .C (clk), .D (new_AGEMA_signal_12202), .Q (new_AGEMA_signal_12203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4382 ( .C (clk), .D (new_AGEMA_signal_12206), .Q (new_AGEMA_signal_12207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4386 ( .C (clk), .D (new_AGEMA_signal_12210), .Q (new_AGEMA_signal_12211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4390 ( .C (clk), .D (new_AGEMA_signal_12214), .Q (new_AGEMA_signal_12215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4394 ( .C (clk), .D (new_AGEMA_signal_12218), .Q (new_AGEMA_signal_12219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4398 ( .C (clk), .D (new_AGEMA_signal_12222), .Q (new_AGEMA_signal_12223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4402 ( .C (clk), .D (new_AGEMA_signal_12226), .Q (new_AGEMA_signal_12227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4406 ( .C (clk), .D (new_AGEMA_signal_12230), .Q (new_AGEMA_signal_12231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4410 ( .C (clk), .D (new_AGEMA_signal_12234), .Q (new_AGEMA_signal_12235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4414 ( .C (clk), .D (new_AGEMA_signal_12238), .Q (new_AGEMA_signal_12239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4418 ( .C (clk), .D (new_AGEMA_signal_12242), .Q (new_AGEMA_signal_12243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4422 ( .C (clk), .D (new_AGEMA_signal_12246), .Q (new_AGEMA_signal_12247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4426 ( .C (clk), .D (new_AGEMA_signal_12250), .Q (new_AGEMA_signal_12251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4430 ( .C (clk), .D (new_AGEMA_signal_12254), .Q (new_AGEMA_signal_12255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4434 ( .C (clk), .D (new_AGEMA_signal_12258), .Q (new_AGEMA_signal_12259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4438 ( .C (clk), .D (new_AGEMA_signal_12262), .Q (new_AGEMA_signal_12263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4442 ( .C (clk), .D (new_AGEMA_signal_12266), .Q (new_AGEMA_signal_12267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4446 ( .C (clk), .D (new_AGEMA_signal_12270), .Q (new_AGEMA_signal_12271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4450 ( .C (clk), .D (new_AGEMA_signal_12274), .Q (new_AGEMA_signal_12275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4454 ( .C (clk), .D (new_AGEMA_signal_12278), .Q (new_AGEMA_signal_12279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4458 ( .C (clk), .D (new_AGEMA_signal_12282), .Q (new_AGEMA_signal_12283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4462 ( .C (clk), .D (new_AGEMA_signal_12286), .Q (new_AGEMA_signal_12287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4466 ( .C (clk), .D (new_AGEMA_signal_12290), .Q (new_AGEMA_signal_12291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4470 ( .C (clk), .D (new_AGEMA_signal_12294), .Q (new_AGEMA_signal_12295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4474 ( .C (clk), .D (new_AGEMA_signal_12298), .Q (new_AGEMA_signal_12299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4478 ( .C (clk), .D (new_AGEMA_signal_12302), .Q (new_AGEMA_signal_12303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4482 ( .C (clk), .D (new_AGEMA_signal_12306), .Q (new_AGEMA_signal_12307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4486 ( .C (clk), .D (new_AGEMA_signal_12310), .Q (new_AGEMA_signal_12311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4490 ( .C (clk), .D (new_AGEMA_signal_12314), .Q (new_AGEMA_signal_12315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4494 ( .C (clk), .D (new_AGEMA_signal_12318), .Q (new_AGEMA_signal_12319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4498 ( .C (clk), .D (new_AGEMA_signal_12322), .Q (new_AGEMA_signal_12323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4502 ( .C (clk), .D (new_AGEMA_signal_12326), .Q (new_AGEMA_signal_12327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4506 ( .C (clk), .D (new_AGEMA_signal_12330), .Q (new_AGEMA_signal_12331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4510 ( .C (clk), .D (new_AGEMA_signal_12334), .Q (new_AGEMA_signal_12335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4514 ( .C (clk), .D (new_AGEMA_signal_12338), .Q (new_AGEMA_signal_12339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4518 ( .C (clk), .D (new_AGEMA_signal_12342), .Q (new_AGEMA_signal_12343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4522 ( .C (clk), .D (new_AGEMA_signal_12346), .Q (new_AGEMA_signal_12347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4526 ( .C (clk), .D (new_AGEMA_signal_12350), .Q (new_AGEMA_signal_12351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4530 ( .C (clk), .D (new_AGEMA_signal_12354), .Q (new_AGEMA_signal_12355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4534 ( .C (clk), .D (new_AGEMA_signal_12358), .Q (new_AGEMA_signal_12359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4538 ( .C (clk), .D (new_AGEMA_signal_12362), .Q (new_AGEMA_signal_12363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4542 ( .C (clk), .D (new_AGEMA_signal_12366), .Q (new_AGEMA_signal_12367) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4546 ( .C (clk), .D (new_AGEMA_signal_12370), .Q (new_AGEMA_signal_12371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4550 ( .C (clk), .D (new_AGEMA_signal_12374), .Q (new_AGEMA_signal_12375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4554 ( .C (clk), .D (new_AGEMA_signal_12378), .Q (new_AGEMA_signal_12379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4558 ( .C (clk), .D (new_AGEMA_signal_12382), .Q (new_AGEMA_signal_12383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4562 ( .C (clk), .D (new_AGEMA_signal_12386), .Q (new_AGEMA_signal_12387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4566 ( .C (clk), .D (new_AGEMA_signal_12390), .Q (new_AGEMA_signal_12391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4570 ( .C (clk), .D (new_AGEMA_signal_12394), .Q (new_AGEMA_signal_12395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4574 ( .C (clk), .D (new_AGEMA_signal_12398), .Q (new_AGEMA_signal_12399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4578 ( .C (clk), .D (new_AGEMA_signal_12402), .Q (new_AGEMA_signal_12403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4582 ( .C (clk), .D (new_AGEMA_signal_12406), .Q (new_AGEMA_signal_12407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4586 ( .C (clk), .D (new_AGEMA_signal_12410), .Q (new_AGEMA_signal_12411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4590 ( .C (clk), .D (new_AGEMA_signal_12414), .Q (new_AGEMA_signal_12415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4594 ( .C (clk), .D (new_AGEMA_signal_12418), .Q (new_AGEMA_signal_12419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4598 ( .C (clk), .D (new_AGEMA_signal_12422), .Q (new_AGEMA_signal_12423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4602 ( .C (clk), .D (new_AGEMA_signal_12426), .Q (new_AGEMA_signal_12427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4606 ( .C (clk), .D (new_AGEMA_signal_12430), .Q (new_AGEMA_signal_12431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4610 ( .C (clk), .D (new_AGEMA_signal_12434), .Q (new_AGEMA_signal_12435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4614 ( .C (clk), .D (new_AGEMA_signal_12438), .Q (new_AGEMA_signal_12439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4618 ( .C (clk), .D (new_AGEMA_signal_12442), .Q (new_AGEMA_signal_12443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4622 ( .C (clk), .D (new_AGEMA_signal_12446), .Q (new_AGEMA_signal_12447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4626 ( .C (clk), .D (new_AGEMA_signal_12450), .Q (new_AGEMA_signal_12451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4630 ( .C (clk), .D (new_AGEMA_signal_12454), .Q (new_AGEMA_signal_12455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4634 ( .C (clk), .D (new_AGEMA_signal_12458), .Q (new_AGEMA_signal_12459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4638 ( .C (clk), .D (new_AGEMA_signal_12462), .Q (new_AGEMA_signal_12463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4642 ( .C (clk), .D (new_AGEMA_signal_12466), .Q (new_AGEMA_signal_12467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4646 ( .C (clk), .D (new_AGEMA_signal_12470), .Q (new_AGEMA_signal_12471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4650 ( .C (clk), .D (new_AGEMA_signal_12474), .Q (new_AGEMA_signal_12475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4654 ( .C (clk), .D (new_AGEMA_signal_12478), .Q (new_AGEMA_signal_12479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4658 ( .C (clk), .D (new_AGEMA_signal_12482), .Q (new_AGEMA_signal_12483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4662 ( .C (clk), .D (new_AGEMA_signal_12486), .Q (new_AGEMA_signal_12487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4666 ( .C (clk), .D (new_AGEMA_signal_12490), .Q (new_AGEMA_signal_12491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4670 ( .C (clk), .D (new_AGEMA_signal_12494), .Q (new_AGEMA_signal_12495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4674 ( .C (clk), .D (new_AGEMA_signal_12498), .Q (new_AGEMA_signal_12499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4678 ( .C (clk), .D (new_AGEMA_signal_12502), .Q (new_AGEMA_signal_12503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4682 ( .C (clk), .D (new_AGEMA_signal_12506), .Q (new_AGEMA_signal_12507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4686 ( .C (clk), .D (new_AGEMA_signal_12510), .Q (new_AGEMA_signal_12511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4690 ( .C (clk), .D (new_AGEMA_signal_12514), .Q (new_AGEMA_signal_12515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4694 ( .C (clk), .D (new_AGEMA_signal_12518), .Q (new_AGEMA_signal_12519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4698 ( .C (clk), .D (new_AGEMA_signal_12522), .Q (new_AGEMA_signal_12523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4702 ( .C (clk), .D (new_AGEMA_signal_12526), .Q (new_AGEMA_signal_12527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4706 ( .C (clk), .D (new_AGEMA_signal_12530), .Q (new_AGEMA_signal_12531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4710 ( .C (clk), .D (new_AGEMA_signal_12534), .Q (new_AGEMA_signal_12535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4714 ( .C (clk), .D (new_AGEMA_signal_12538), .Q (new_AGEMA_signal_12539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4718 ( .C (clk), .D (new_AGEMA_signal_12542), .Q (new_AGEMA_signal_12543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4722 ( .C (clk), .D (new_AGEMA_signal_12546), .Q (new_AGEMA_signal_12547) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4726 ( .C (clk), .D (new_AGEMA_signal_12550), .Q (new_AGEMA_signal_12551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4730 ( .C (clk), .D (new_AGEMA_signal_12554), .Q (new_AGEMA_signal_12555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4734 ( .C (clk), .D (new_AGEMA_signal_12558), .Q (new_AGEMA_signal_12559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4738 ( .C (clk), .D (new_AGEMA_signal_12562), .Q (new_AGEMA_signal_12563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4742 ( .C (clk), .D (new_AGEMA_signal_12566), .Q (new_AGEMA_signal_12567) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4746 ( .C (clk), .D (new_AGEMA_signal_12570), .Q (new_AGEMA_signal_12571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4750 ( .C (clk), .D (new_AGEMA_signal_12574), .Q (new_AGEMA_signal_12575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4754 ( .C (clk), .D (new_AGEMA_signal_12578), .Q (new_AGEMA_signal_12579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4758 ( .C (clk), .D (new_AGEMA_signal_12582), .Q (new_AGEMA_signal_12583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4762 ( .C (clk), .D (new_AGEMA_signal_12586), .Q (new_AGEMA_signal_12587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4766 ( .C (clk), .D (new_AGEMA_signal_12590), .Q (new_AGEMA_signal_12591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4770 ( .C (clk), .D (new_AGEMA_signal_12594), .Q (new_AGEMA_signal_12595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4774 ( .C (clk), .D (new_AGEMA_signal_12598), .Q (new_AGEMA_signal_12599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4778 ( .C (clk), .D (new_AGEMA_signal_12602), .Q (new_AGEMA_signal_12603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4782 ( .C (clk), .D (new_AGEMA_signal_12606), .Q (new_AGEMA_signal_12607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4786 ( .C (clk), .D (new_AGEMA_signal_12610), .Q (new_AGEMA_signal_12611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4790 ( .C (clk), .D (new_AGEMA_signal_12614), .Q (new_AGEMA_signal_12615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4794 ( .C (clk), .D (new_AGEMA_signal_12618), .Q (new_AGEMA_signal_12619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4798 ( .C (clk), .D (new_AGEMA_signal_12622), .Q (new_AGEMA_signal_12623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4802 ( .C (clk), .D (new_AGEMA_signal_12626), .Q (new_AGEMA_signal_12627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4806 ( .C (clk), .D (new_AGEMA_signal_12630), .Q (new_AGEMA_signal_12631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4810 ( .C (clk), .D (new_AGEMA_signal_12634), .Q (new_AGEMA_signal_12635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4814 ( .C (clk), .D (new_AGEMA_signal_12638), .Q (new_AGEMA_signal_12639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4818 ( .C (clk), .D (new_AGEMA_signal_12642), .Q (new_AGEMA_signal_12643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4822 ( .C (clk), .D (new_AGEMA_signal_12646), .Q (new_AGEMA_signal_12647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4826 ( .C (clk), .D (new_AGEMA_signal_12650), .Q (new_AGEMA_signal_12651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4830 ( .C (clk), .D (new_AGEMA_signal_12654), .Q (new_AGEMA_signal_12655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4834 ( .C (clk), .D (new_AGEMA_signal_12658), .Q (new_AGEMA_signal_12659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4838 ( .C (clk), .D (new_AGEMA_signal_12662), .Q (new_AGEMA_signal_12663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4842 ( .C (clk), .D (new_AGEMA_signal_12666), .Q (new_AGEMA_signal_12667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4846 ( .C (clk), .D (new_AGEMA_signal_12670), .Q (new_AGEMA_signal_12671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4850 ( .C (clk), .D (new_AGEMA_signal_12674), .Q (new_AGEMA_signal_12675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4854 ( .C (clk), .D (new_AGEMA_signal_12678), .Q (new_AGEMA_signal_12679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4858 ( .C (clk), .D (new_AGEMA_signal_12682), .Q (new_AGEMA_signal_12683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4862 ( .C (clk), .D (new_AGEMA_signal_12686), .Q (new_AGEMA_signal_12687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4866 ( .C (clk), .D (new_AGEMA_signal_12690), .Q (new_AGEMA_signal_12691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4870 ( .C (clk), .D (new_AGEMA_signal_12694), .Q (new_AGEMA_signal_12695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4874 ( .C (clk), .D (new_AGEMA_signal_12698), .Q (new_AGEMA_signal_12699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4878 ( .C (clk), .D (new_AGEMA_signal_12702), .Q (new_AGEMA_signal_12703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4882 ( .C (clk), .D (new_AGEMA_signal_12706), .Q (new_AGEMA_signal_12707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4886 ( .C (clk), .D (new_AGEMA_signal_12710), .Q (new_AGEMA_signal_12711) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4890 ( .C (clk), .D (new_AGEMA_signal_12714), .Q (new_AGEMA_signal_12715) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4894 ( .C (clk), .D (new_AGEMA_signal_12718), .Q (new_AGEMA_signal_12719) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4898 ( .C (clk), .D (new_AGEMA_signal_12722), .Q (new_AGEMA_signal_12723) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4902 ( .C (clk), .D (new_AGEMA_signal_12726), .Q (new_AGEMA_signal_12727) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4906 ( .C (clk), .D (new_AGEMA_signal_12730), .Q (new_AGEMA_signal_12731) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4910 ( .C (clk), .D (new_AGEMA_signal_12734), .Q (new_AGEMA_signal_12735) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4914 ( .C (clk), .D (new_AGEMA_signal_12738), .Q (new_AGEMA_signal_12739) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4918 ( .C (clk), .D (new_AGEMA_signal_12742), .Q (new_AGEMA_signal_12743) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4922 ( .C (clk), .D (new_AGEMA_signal_12746), .Q (new_AGEMA_signal_12747) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4926 ( .C (clk), .D (new_AGEMA_signal_12750), .Q (new_AGEMA_signal_12751) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4930 ( .C (clk), .D (new_AGEMA_signal_12754), .Q (new_AGEMA_signal_12755) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4934 ( .C (clk), .D (new_AGEMA_signal_12758), .Q (new_AGEMA_signal_12759) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4938 ( .C (clk), .D (new_AGEMA_signal_12762), .Q (new_AGEMA_signal_12763) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4942 ( .C (clk), .D (new_AGEMA_signal_12766), .Q (new_AGEMA_signal_12767) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4946 ( .C (clk), .D (new_AGEMA_signal_12770), .Q (new_AGEMA_signal_12771) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4950 ( .C (clk), .D (new_AGEMA_signal_12774), .Q (new_AGEMA_signal_12775) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4954 ( .C (clk), .D (new_AGEMA_signal_12778), .Q (new_AGEMA_signal_12779) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4958 ( .C (clk), .D (new_AGEMA_signal_12782), .Q (new_AGEMA_signal_12783) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4962 ( .C (clk), .D (new_AGEMA_signal_12786), .Q (new_AGEMA_signal_12787) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4966 ( .C (clk), .D (new_AGEMA_signal_12790), .Q (new_AGEMA_signal_12791) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4970 ( .C (clk), .D (new_AGEMA_signal_12794), .Q (new_AGEMA_signal_12795) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4974 ( .C (clk), .D (new_AGEMA_signal_12798), .Q (new_AGEMA_signal_12799) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4978 ( .C (clk), .D (new_AGEMA_signal_12802), .Q (new_AGEMA_signal_12803) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4982 ( .C (clk), .D (new_AGEMA_signal_12806), .Q (new_AGEMA_signal_12807) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4986 ( .C (clk), .D (new_AGEMA_signal_12810), .Q (new_AGEMA_signal_12811) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4990 ( .C (clk), .D (new_AGEMA_signal_12814), .Q (new_AGEMA_signal_12815) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4994 ( .C (clk), .D (new_AGEMA_signal_12818), .Q (new_AGEMA_signal_12819) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4998 ( .C (clk), .D (new_AGEMA_signal_12822), .Q (new_AGEMA_signal_12823) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5002 ( .C (clk), .D (new_AGEMA_signal_12826), .Q (new_AGEMA_signal_12827) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5006 ( .C (clk), .D (new_AGEMA_signal_12830), .Q (new_AGEMA_signal_12831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5010 ( .C (clk), .D (new_AGEMA_signal_12834), .Q (new_AGEMA_signal_12835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5014 ( .C (clk), .D (new_AGEMA_signal_12838), .Q (new_AGEMA_signal_12839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5018 ( .C (clk), .D (new_AGEMA_signal_12842), .Q (new_AGEMA_signal_12843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5022 ( .C (clk), .D (new_AGEMA_signal_12846), .Q (new_AGEMA_signal_12847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5026 ( .C (clk), .D (new_AGEMA_signal_12850), .Q (new_AGEMA_signal_12851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5030 ( .C (clk), .D (new_AGEMA_signal_12854), .Q (new_AGEMA_signal_12855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5034 ( .C (clk), .D (new_AGEMA_signal_12858), .Q (new_AGEMA_signal_12859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5038 ( .C (clk), .D (new_AGEMA_signal_12862), .Q (new_AGEMA_signal_12863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5042 ( .C (clk), .D (new_AGEMA_signal_12866), .Q (new_AGEMA_signal_12867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5046 ( .C (clk), .D (new_AGEMA_signal_12870), .Q (new_AGEMA_signal_12871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5050 ( .C (clk), .D (new_AGEMA_signal_12874), .Q (new_AGEMA_signal_12875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5054 ( .C (clk), .D (new_AGEMA_signal_12878), .Q (new_AGEMA_signal_12879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5058 ( .C (clk), .D (new_AGEMA_signal_12882), .Q (new_AGEMA_signal_12883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5062 ( .C (clk), .D (new_AGEMA_signal_12886), .Q (new_AGEMA_signal_12887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5066 ( .C (clk), .D (new_AGEMA_signal_12890), .Q (new_AGEMA_signal_12891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5070 ( .C (clk), .D (new_AGEMA_signal_12894), .Q (new_AGEMA_signal_12895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5074 ( .C (clk), .D (new_AGEMA_signal_12898), .Q (new_AGEMA_signal_12899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5078 ( .C (clk), .D (new_AGEMA_signal_12902), .Q (new_AGEMA_signal_12903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5082 ( .C (clk), .D (new_AGEMA_signal_12906), .Q (new_AGEMA_signal_12907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5086 ( .C (clk), .D (new_AGEMA_signal_12910), .Q (new_AGEMA_signal_12911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5090 ( .C (clk), .D (new_AGEMA_signal_12914), .Q (new_AGEMA_signal_12915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5094 ( .C (clk), .D (new_AGEMA_signal_12918), .Q (new_AGEMA_signal_12919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5098 ( .C (clk), .D (new_AGEMA_signal_12922), .Q (new_AGEMA_signal_12923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5102 ( .C (clk), .D (new_AGEMA_signal_12926), .Q (new_AGEMA_signal_12927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5106 ( .C (clk), .D (new_AGEMA_signal_12930), .Q (new_AGEMA_signal_12931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5110 ( .C (clk), .D (new_AGEMA_signal_12934), .Q (new_AGEMA_signal_12935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5114 ( .C (clk), .D (new_AGEMA_signal_12938), .Q (new_AGEMA_signal_12939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5118 ( .C (clk), .D (new_AGEMA_signal_12942), .Q (new_AGEMA_signal_12943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5122 ( .C (clk), .D (new_AGEMA_signal_12946), .Q (new_AGEMA_signal_12947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5126 ( .C (clk), .D (new_AGEMA_signal_12950), .Q (new_AGEMA_signal_12951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5130 ( .C (clk), .D (new_AGEMA_signal_12954), .Q (new_AGEMA_signal_12955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5134 ( .C (clk), .D (new_AGEMA_signal_12958), .Q (new_AGEMA_signal_12959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5138 ( .C (clk), .D (new_AGEMA_signal_12962), .Q (new_AGEMA_signal_12963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5142 ( .C (clk), .D (new_AGEMA_signal_12966), .Q (new_AGEMA_signal_12967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5146 ( .C (clk), .D (new_AGEMA_signal_12970), .Q (new_AGEMA_signal_12971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5150 ( .C (clk), .D (new_AGEMA_signal_12974), .Q (new_AGEMA_signal_12975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5154 ( .C (clk), .D (new_AGEMA_signal_12978), .Q (new_AGEMA_signal_12979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5158 ( .C (clk), .D (new_AGEMA_signal_12982), .Q (new_AGEMA_signal_12983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5162 ( .C (clk), .D (new_AGEMA_signal_12986), .Q (new_AGEMA_signal_12987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5166 ( .C (clk), .D (new_AGEMA_signal_12990), .Q (new_AGEMA_signal_12991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5170 ( .C (clk), .D (new_AGEMA_signal_12994), .Q (new_AGEMA_signal_12995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5174 ( .C (clk), .D (new_AGEMA_signal_12998), .Q (new_AGEMA_signal_12999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5178 ( .C (clk), .D (new_AGEMA_signal_13002), .Q (new_AGEMA_signal_13003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5182 ( .C (clk), .D (new_AGEMA_signal_13006), .Q (new_AGEMA_signal_13007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5186 ( .C (clk), .D (new_AGEMA_signal_13010), .Q (new_AGEMA_signal_13011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5190 ( .C (clk), .D (new_AGEMA_signal_13014), .Q (new_AGEMA_signal_13015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5194 ( .C (clk), .D (new_AGEMA_signal_13018), .Q (new_AGEMA_signal_13019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5198 ( .C (clk), .D (new_AGEMA_signal_13022), .Q (new_AGEMA_signal_13023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5202 ( .C (clk), .D (new_AGEMA_signal_13026), .Q (new_AGEMA_signal_13027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5206 ( .C (clk), .D (new_AGEMA_signal_13030), .Q (new_AGEMA_signal_13031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5210 ( .C (clk), .D (new_AGEMA_signal_13034), .Q (new_AGEMA_signal_13035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5214 ( .C (clk), .D (new_AGEMA_signal_13038), .Q (new_AGEMA_signal_13039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5218 ( .C (clk), .D (new_AGEMA_signal_13042), .Q (new_AGEMA_signal_13043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5222 ( .C (clk), .D (new_AGEMA_signal_13046), .Q (new_AGEMA_signal_13047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5226 ( .C (clk), .D (new_AGEMA_signal_13050), .Q (new_AGEMA_signal_13051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5230 ( .C (clk), .D (new_AGEMA_signal_13054), .Q (new_AGEMA_signal_13055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5234 ( .C (clk), .D (new_AGEMA_signal_13058), .Q (new_AGEMA_signal_13059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5238 ( .C (clk), .D (new_AGEMA_signal_13062), .Q (new_AGEMA_signal_13063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5242 ( .C (clk), .D (new_AGEMA_signal_13066), .Q (new_AGEMA_signal_13067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5246 ( .C (clk), .D (new_AGEMA_signal_13070), .Q (new_AGEMA_signal_13071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5250 ( .C (clk), .D (new_AGEMA_signal_13074), .Q (new_AGEMA_signal_13075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5254 ( .C (clk), .D (new_AGEMA_signal_13078), .Q (new_AGEMA_signal_13079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5258 ( .C (clk), .D (new_AGEMA_signal_13082), .Q (new_AGEMA_signal_13083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5262 ( .C (clk), .D (new_AGEMA_signal_13086), .Q (new_AGEMA_signal_13087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5266 ( .C (clk), .D (new_AGEMA_signal_13090), .Q (new_AGEMA_signal_13091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5270 ( .C (clk), .D (new_AGEMA_signal_13094), .Q (new_AGEMA_signal_13095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5274 ( .C (clk), .D (new_AGEMA_signal_13098), .Q (new_AGEMA_signal_13099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5278 ( .C (clk), .D (new_AGEMA_signal_13102), .Q (new_AGEMA_signal_13103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5282 ( .C (clk), .D (new_AGEMA_signal_13106), .Q (new_AGEMA_signal_13107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5286 ( .C (clk), .D (new_AGEMA_signal_13110), .Q (new_AGEMA_signal_13111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5290 ( .C (clk), .D (new_AGEMA_signal_13114), .Q (new_AGEMA_signal_13115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5294 ( .C (clk), .D (new_AGEMA_signal_13118), .Q (new_AGEMA_signal_13119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5298 ( .C (clk), .D (new_AGEMA_signal_13122), .Q (new_AGEMA_signal_13123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5302 ( .C (clk), .D (new_AGEMA_signal_13126), .Q (new_AGEMA_signal_13127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5306 ( .C (clk), .D (new_AGEMA_signal_13130), .Q (new_AGEMA_signal_13131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5310 ( .C (clk), .D (new_AGEMA_signal_13134), .Q (new_AGEMA_signal_13135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5314 ( .C (clk), .D (new_AGEMA_signal_13138), .Q (new_AGEMA_signal_13139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5318 ( .C (clk), .D (new_AGEMA_signal_13142), .Q (new_AGEMA_signal_13143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5322 ( .C (clk), .D (new_AGEMA_signal_13146), .Q (new_AGEMA_signal_13147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5326 ( .C (clk), .D (new_AGEMA_signal_13150), .Q (new_AGEMA_signal_13151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5330 ( .C (clk), .D (new_AGEMA_signal_13154), .Q (new_AGEMA_signal_13155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5334 ( .C (clk), .D (new_AGEMA_signal_13158), .Q (new_AGEMA_signal_13159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5338 ( .C (clk), .D (new_AGEMA_signal_13162), .Q (new_AGEMA_signal_13163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5342 ( .C (clk), .D (new_AGEMA_signal_13166), .Q (new_AGEMA_signal_13167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5346 ( .C (clk), .D (new_AGEMA_signal_13170), .Q (new_AGEMA_signal_13171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5350 ( .C (clk), .D (new_AGEMA_signal_13174), .Q (new_AGEMA_signal_13175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5354 ( .C (clk), .D (new_AGEMA_signal_13178), .Q (new_AGEMA_signal_13179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5358 ( .C (clk), .D (new_AGEMA_signal_13182), .Q (new_AGEMA_signal_13183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5362 ( .C (clk), .D (new_AGEMA_signal_13186), .Q (new_AGEMA_signal_13187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5366 ( .C (clk), .D (new_AGEMA_signal_13190), .Q (new_AGEMA_signal_13191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5370 ( .C (clk), .D (new_AGEMA_signal_13194), .Q (new_AGEMA_signal_13195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5374 ( .C (clk), .D (new_AGEMA_signal_13198), .Q (new_AGEMA_signal_13199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5378 ( .C (clk), .D (new_AGEMA_signal_13202), .Q (new_AGEMA_signal_13203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5382 ( .C (clk), .D (new_AGEMA_signal_13206), .Q (new_AGEMA_signal_13207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5386 ( .C (clk), .D (new_AGEMA_signal_13210), .Q (new_AGEMA_signal_13211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5390 ( .C (clk), .D (new_AGEMA_signal_13214), .Q (new_AGEMA_signal_13215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5394 ( .C (clk), .D (new_AGEMA_signal_13218), .Q (new_AGEMA_signal_13219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5398 ( .C (clk), .D (new_AGEMA_signal_13222), .Q (new_AGEMA_signal_13223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5402 ( .C (clk), .D (new_AGEMA_signal_13226), .Q (new_AGEMA_signal_13227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5406 ( .C (clk), .D (new_AGEMA_signal_13230), .Q (new_AGEMA_signal_13231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5410 ( .C (clk), .D (new_AGEMA_signal_13234), .Q (new_AGEMA_signal_13235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5414 ( .C (clk), .D (new_AGEMA_signal_13238), .Q (new_AGEMA_signal_13239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5418 ( .C (clk), .D (new_AGEMA_signal_13242), .Q (new_AGEMA_signal_13243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5422 ( .C (clk), .D (new_AGEMA_signal_13246), .Q (new_AGEMA_signal_13247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5426 ( .C (clk), .D (new_AGEMA_signal_13250), .Q (new_AGEMA_signal_13251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5430 ( .C (clk), .D (new_AGEMA_signal_13254), .Q (new_AGEMA_signal_13255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5434 ( .C (clk), .D (new_AGEMA_signal_13258), .Q (new_AGEMA_signal_13259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5438 ( .C (clk), .D (new_AGEMA_signal_13262), .Q (new_AGEMA_signal_13263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5442 ( .C (clk), .D (new_AGEMA_signal_13266), .Q (new_AGEMA_signal_13267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5446 ( .C (clk), .D (new_AGEMA_signal_13270), .Q (new_AGEMA_signal_13271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5450 ( .C (clk), .D (new_AGEMA_signal_13274), .Q (new_AGEMA_signal_13275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5454 ( .C (clk), .D (new_AGEMA_signal_13278), .Q (new_AGEMA_signal_13279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5458 ( .C (clk), .D (new_AGEMA_signal_13282), .Q (new_AGEMA_signal_13283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5462 ( .C (clk), .D (new_AGEMA_signal_13286), .Q (new_AGEMA_signal_13287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5466 ( .C (clk), .D (new_AGEMA_signal_13290), .Q (new_AGEMA_signal_13291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5470 ( .C (clk), .D (new_AGEMA_signal_13294), .Q (new_AGEMA_signal_13295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5474 ( .C (clk), .D (new_AGEMA_signal_13298), .Q (new_AGEMA_signal_13299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5478 ( .C (clk), .D (new_AGEMA_signal_13302), .Q (new_AGEMA_signal_13303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5482 ( .C (clk), .D (new_AGEMA_signal_13306), .Q (new_AGEMA_signal_13307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5486 ( .C (clk), .D (new_AGEMA_signal_13310), .Q (new_AGEMA_signal_13311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5490 ( .C (clk), .D (new_AGEMA_signal_13314), .Q (new_AGEMA_signal_13315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5494 ( .C (clk), .D (new_AGEMA_signal_13318), .Q (new_AGEMA_signal_13319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5498 ( .C (clk), .D (new_AGEMA_signal_13322), .Q (new_AGEMA_signal_13323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5502 ( .C (clk), .D (new_AGEMA_signal_13326), .Q (new_AGEMA_signal_13327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5506 ( .C (clk), .D (new_AGEMA_signal_13330), .Q (new_AGEMA_signal_13331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5510 ( .C (clk), .D (new_AGEMA_signal_13334), .Q (new_AGEMA_signal_13335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5514 ( .C (clk), .D (new_AGEMA_signal_13338), .Q (new_AGEMA_signal_13339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5518 ( .C (clk), .D (new_AGEMA_signal_13342), .Q (new_AGEMA_signal_13343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5522 ( .C (clk), .D (new_AGEMA_signal_13346), .Q (new_AGEMA_signal_13347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5526 ( .C (clk), .D (new_AGEMA_signal_13350), .Q (new_AGEMA_signal_13351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5530 ( .C (clk), .D (new_AGEMA_signal_13354), .Q (new_AGEMA_signal_13355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5534 ( .C (clk), .D (new_AGEMA_signal_13358), .Q (new_AGEMA_signal_13359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5538 ( .C (clk), .D (new_AGEMA_signal_13362), .Q (new_AGEMA_signal_13363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5542 ( .C (clk), .D (new_AGEMA_signal_13366), .Q (new_AGEMA_signal_13367) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5546 ( .C (clk), .D (new_AGEMA_signal_13370), .Q (new_AGEMA_signal_13371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5550 ( .C (clk), .D (new_AGEMA_signal_13374), .Q (new_AGEMA_signal_13375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5554 ( .C (clk), .D (new_AGEMA_signal_13378), .Q (new_AGEMA_signal_13379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5558 ( .C (clk), .D (new_AGEMA_signal_13382), .Q (new_AGEMA_signal_13383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5562 ( .C (clk), .D (new_AGEMA_signal_13386), .Q (new_AGEMA_signal_13387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5566 ( .C (clk), .D (new_AGEMA_signal_13390), .Q (new_AGEMA_signal_13391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5570 ( .C (clk), .D (new_AGEMA_signal_13394), .Q (new_AGEMA_signal_13395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5574 ( .C (clk), .D (new_AGEMA_signal_13398), .Q (new_AGEMA_signal_13399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5578 ( .C (clk), .D (new_AGEMA_signal_13402), .Q (new_AGEMA_signal_13403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5582 ( .C (clk), .D (new_AGEMA_signal_13406), .Q (new_AGEMA_signal_13407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5586 ( .C (clk), .D (new_AGEMA_signal_13410), .Q (new_AGEMA_signal_13411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5590 ( .C (clk), .D (new_AGEMA_signal_13414), .Q (new_AGEMA_signal_13415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5594 ( .C (clk), .D (new_AGEMA_signal_13418), .Q (new_AGEMA_signal_13419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5598 ( .C (clk), .D (new_AGEMA_signal_13422), .Q (new_AGEMA_signal_13423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5602 ( .C (clk), .D (new_AGEMA_signal_13426), .Q (new_AGEMA_signal_13427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5606 ( .C (clk), .D (new_AGEMA_signal_13430), .Q (new_AGEMA_signal_13431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5610 ( .C (clk), .D (new_AGEMA_signal_13434), .Q (new_AGEMA_signal_13435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5614 ( .C (clk), .D (new_AGEMA_signal_13438), .Q (new_AGEMA_signal_13439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5618 ( .C (clk), .D (new_AGEMA_signal_13442), .Q (new_AGEMA_signal_13443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5622 ( .C (clk), .D (new_AGEMA_signal_13446), .Q (new_AGEMA_signal_13447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5626 ( .C (clk), .D (new_AGEMA_signal_13450), .Q (new_AGEMA_signal_13451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5630 ( .C (clk), .D (new_AGEMA_signal_13454), .Q (new_AGEMA_signal_13455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5634 ( .C (clk), .D (new_AGEMA_signal_13458), .Q (new_AGEMA_signal_13459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5638 ( .C (clk), .D (new_AGEMA_signal_13462), .Q (new_AGEMA_signal_13463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5642 ( .C (clk), .D (new_AGEMA_signal_13466), .Q (new_AGEMA_signal_13467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5646 ( .C (clk), .D (new_AGEMA_signal_13470), .Q (new_AGEMA_signal_13471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5650 ( .C (clk), .D (new_AGEMA_signal_13474), .Q (new_AGEMA_signal_13475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5654 ( .C (clk), .D (new_AGEMA_signal_13478), .Q (new_AGEMA_signal_13479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5658 ( .C (clk), .D (new_AGEMA_signal_13482), .Q (new_AGEMA_signal_13483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5662 ( .C (clk), .D (new_AGEMA_signal_13486), .Q (new_AGEMA_signal_13487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5666 ( .C (clk), .D (new_AGEMA_signal_13490), .Q (new_AGEMA_signal_13491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5670 ( .C (clk), .D (new_AGEMA_signal_13494), .Q (new_AGEMA_signal_13495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5674 ( .C (clk), .D (new_AGEMA_signal_13498), .Q (new_AGEMA_signal_13499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5678 ( .C (clk), .D (new_AGEMA_signal_13502), .Q (new_AGEMA_signal_13503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5682 ( .C (clk), .D (new_AGEMA_signal_13506), .Q (new_AGEMA_signal_13507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5686 ( .C (clk), .D (new_AGEMA_signal_13510), .Q (new_AGEMA_signal_13511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5690 ( .C (clk), .D (new_AGEMA_signal_13514), .Q (new_AGEMA_signal_13515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5694 ( .C (clk), .D (new_AGEMA_signal_13518), .Q (new_AGEMA_signal_13519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5698 ( .C (clk), .D (new_AGEMA_signal_13522), .Q (new_AGEMA_signal_13523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5702 ( .C (clk), .D (new_AGEMA_signal_13526), .Q (new_AGEMA_signal_13527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5706 ( .C (clk), .D (new_AGEMA_signal_13530), .Q (new_AGEMA_signal_13531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5710 ( .C (clk), .D (new_AGEMA_signal_13534), .Q (new_AGEMA_signal_13535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5714 ( .C (clk), .D (new_AGEMA_signal_13538), .Q (new_AGEMA_signal_13539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5718 ( .C (clk), .D (new_AGEMA_signal_13542), .Q (new_AGEMA_signal_13543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5722 ( .C (clk), .D (new_AGEMA_signal_13546), .Q (new_AGEMA_signal_13547) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5726 ( .C (clk), .D (new_AGEMA_signal_13550), .Q (new_AGEMA_signal_13551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5730 ( .C (clk), .D (new_AGEMA_signal_13554), .Q (new_AGEMA_signal_13555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5734 ( .C (clk), .D (new_AGEMA_signal_13558), .Q (new_AGEMA_signal_13559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5738 ( .C (clk), .D (new_AGEMA_signal_13562), .Q (new_AGEMA_signal_13563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5742 ( .C (clk), .D (new_AGEMA_signal_13566), .Q (new_AGEMA_signal_13567) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5746 ( .C (clk), .D (new_AGEMA_signal_13570), .Q (new_AGEMA_signal_13571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5750 ( .C (clk), .D (new_AGEMA_signal_13574), .Q (new_AGEMA_signal_13575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5754 ( .C (clk), .D (new_AGEMA_signal_13578), .Q (new_AGEMA_signal_13579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5758 ( .C (clk), .D (new_AGEMA_signal_13582), .Q (new_AGEMA_signal_13583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5762 ( .C (clk), .D (new_AGEMA_signal_13586), .Q (new_AGEMA_signal_13587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5766 ( .C (clk), .D (new_AGEMA_signal_13590), .Q (new_AGEMA_signal_13591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5770 ( .C (clk), .D (new_AGEMA_signal_13594), .Q (new_AGEMA_signal_13595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5774 ( .C (clk), .D (new_AGEMA_signal_13598), .Q (new_AGEMA_signal_13599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5778 ( .C (clk), .D (new_AGEMA_signal_13602), .Q (new_AGEMA_signal_13603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5782 ( .C (clk), .D (new_AGEMA_signal_13606), .Q (new_AGEMA_signal_13607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5786 ( .C (clk), .D (new_AGEMA_signal_13610), .Q (new_AGEMA_signal_13611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5790 ( .C (clk), .D (new_AGEMA_signal_13614), .Q (new_AGEMA_signal_13615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5794 ( .C (clk), .D (new_AGEMA_signal_13618), .Q (new_AGEMA_signal_13619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5798 ( .C (clk), .D (new_AGEMA_signal_13622), .Q (new_AGEMA_signal_13623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5802 ( .C (clk), .D (new_AGEMA_signal_13626), .Q (new_AGEMA_signal_13627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5806 ( .C (clk), .D (new_AGEMA_signal_13630), .Q (new_AGEMA_signal_13631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5810 ( .C (clk), .D (new_AGEMA_signal_13634), .Q (new_AGEMA_signal_13635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5814 ( .C (clk), .D (new_AGEMA_signal_13638), .Q (new_AGEMA_signal_13639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5818 ( .C (clk), .D (new_AGEMA_signal_13642), .Q (new_AGEMA_signal_13643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5822 ( .C (clk), .D (new_AGEMA_signal_13646), .Q (new_AGEMA_signal_13647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5826 ( .C (clk), .D (new_AGEMA_signal_13650), .Q (new_AGEMA_signal_13651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5830 ( .C (clk), .D (new_AGEMA_signal_13654), .Q (new_AGEMA_signal_13655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5834 ( .C (clk), .D (new_AGEMA_signal_13658), .Q (new_AGEMA_signal_13659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5838 ( .C (clk), .D (new_AGEMA_signal_13662), .Q (new_AGEMA_signal_13663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5842 ( .C (clk), .D (new_AGEMA_signal_13666), .Q (new_AGEMA_signal_13667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5846 ( .C (clk), .D (new_AGEMA_signal_13670), .Q (new_AGEMA_signal_13671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5850 ( .C (clk), .D (new_AGEMA_signal_13674), .Q (new_AGEMA_signal_13675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5854 ( .C (clk), .D (new_AGEMA_signal_13678), .Q (new_AGEMA_signal_13679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5858 ( .C (clk), .D (new_AGEMA_signal_13682), .Q (new_AGEMA_signal_13683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5862 ( .C (clk), .D (new_AGEMA_signal_13686), .Q (new_AGEMA_signal_13687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5866 ( .C (clk), .D (new_AGEMA_signal_13690), .Q (new_AGEMA_signal_13691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5870 ( .C (clk), .D (new_AGEMA_signal_13694), .Q (new_AGEMA_signal_13695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5874 ( .C (clk), .D (new_AGEMA_signal_13698), .Q (new_AGEMA_signal_13699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5878 ( .C (clk), .D (new_AGEMA_signal_13702), .Q (new_AGEMA_signal_13703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5882 ( .C (clk), .D (new_AGEMA_signal_13706), .Q (new_AGEMA_signal_13707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5886 ( .C (clk), .D (new_AGEMA_signal_13710), .Q (new_AGEMA_signal_13711) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5890 ( .C (clk), .D (new_AGEMA_signal_13714), .Q (new_AGEMA_signal_13715) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5894 ( .C (clk), .D (new_AGEMA_signal_13718), .Q (new_AGEMA_signal_13719) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5898 ( .C (clk), .D (new_AGEMA_signal_13722), .Q (new_AGEMA_signal_13723) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5902 ( .C (clk), .D (new_AGEMA_signal_13726), .Q (new_AGEMA_signal_13727) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5906 ( .C (clk), .D (new_AGEMA_signal_13730), .Q (new_AGEMA_signal_13731) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5910 ( .C (clk), .D (new_AGEMA_signal_13734), .Q (new_AGEMA_signal_13735) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5914 ( .C (clk), .D (new_AGEMA_signal_13738), .Q (new_AGEMA_signal_13739) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5918 ( .C (clk), .D (new_AGEMA_signal_13742), .Q (new_AGEMA_signal_13743) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5922 ( .C (clk), .D (new_AGEMA_signal_13746), .Q (new_AGEMA_signal_13747) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5926 ( .C (clk), .D (new_AGEMA_signal_13750), .Q (new_AGEMA_signal_13751) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5930 ( .C (clk), .D (new_AGEMA_signal_13754), .Q (new_AGEMA_signal_13755) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5934 ( .C (clk), .D (new_AGEMA_signal_13758), .Q (new_AGEMA_signal_13759) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5938 ( .C (clk), .D (new_AGEMA_signal_13762), .Q (new_AGEMA_signal_13763) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5942 ( .C (clk), .D (new_AGEMA_signal_13766), .Q (new_AGEMA_signal_13767) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5946 ( .C (clk), .D (new_AGEMA_signal_13770), .Q (new_AGEMA_signal_13771) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5950 ( .C (clk), .D (new_AGEMA_signal_13774), .Q (new_AGEMA_signal_13775) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5954 ( .C (clk), .D (new_AGEMA_signal_13778), .Q (new_AGEMA_signal_13779) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5958 ( .C (clk), .D (new_AGEMA_signal_13782), .Q (new_AGEMA_signal_13783) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5962 ( .C (clk), .D (new_AGEMA_signal_13786), .Q (new_AGEMA_signal_13787) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5966 ( .C (clk), .D (new_AGEMA_signal_13790), .Q (new_AGEMA_signal_13791) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5970 ( .C (clk), .D (new_AGEMA_signal_13794), .Q (new_AGEMA_signal_13795) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5974 ( .C (clk), .D (new_AGEMA_signal_13798), .Q (new_AGEMA_signal_13799) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5978 ( .C (clk), .D (new_AGEMA_signal_13802), .Q (new_AGEMA_signal_13803) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5982 ( .C (clk), .D (new_AGEMA_signal_13806), .Q (new_AGEMA_signal_13807) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5986 ( .C (clk), .D (new_AGEMA_signal_13810), .Q (new_AGEMA_signal_13811) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5990 ( .C (clk), .D (new_AGEMA_signal_13814), .Q (new_AGEMA_signal_13815) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5994 ( .C (clk), .D (new_AGEMA_signal_13818), .Q (new_AGEMA_signal_13819) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5998 ( .C (clk), .D (new_AGEMA_signal_13822), .Q (new_AGEMA_signal_13823) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6002 ( .C (clk), .D (new_AGEMA_signal_13826), .Q (new_AGEMA_signal_13827) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6006 ( .C (clk), .D (new_AGEMA_signal_13830), .Q (new_AGEMA_signal_13831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6010 ( .C (clk), .D (new_AGEMA_signal_13834), .Q (new_AGEMA_signal_13835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6014 ( .C (clk), .D (new_AGEMA_signal_13838), .Q (new_AGEMA_signal_13839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6018 ( .C (clk), .D (new_AGEMA_signal_13842), .Q (new_AGEMA_signal_13843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6022 ( .C (clk), .D (new_AGEMA_signal_13846), .Q (new_AGEMA_signal_13847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6026 ( .C (clk), .D (new_AGEMA_signal_13850), .Q (new_AGEMA_signal_13851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6030 ( .C (clk), .D (new_AGEMA_signal_13854), .Q (new_AGEMA_signal_13855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6034 ( .C (clk), .D (new_AGEMA_signal_13858), .Q (new_AGEMA_signal_13859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6038 ( .C (clk), .D (new_AGEMA_signal_13862), .Q (new_AGEMA_signal_13863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6042 ( .C (clk), .D (new_AGEMA_signal_13866), .Q (new_AGEMA_signal_13867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6046 ( .C (clk), .D (new_AGEMA_signal_13870), .Q (new_AGEMA_signal_13871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6050 ( .C (clk), .D (new_AGEMA_signal_13874), .Q (new_AGEMA_signal_13875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6054 ( .C (clk), .D (new_AGEMA_signal_13878), .Q (new_AGEMA_signal_13879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6058 ( .C (clk), .D (new_AGEMA_signal_13882), .Q (new_AGEMA_signal_13883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6062 ( .C (clk), .D (new_AGEMA_signal_13886), .Q (new_AGEMA_signal_13887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6066 ( .C (clk), .D (new_AGEMA_signal_13890), .Q (new_AGEMA_signal_13891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6070 ( .C (clk), .D (new_AGEMA_signal_13894), .Q (new_AGEMA_signal_13895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6074 ( .C (clk), .D (new_AGEMA_signal_13898), .Q (new_AGEMA_signal_13899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6078 ( .C (clk), .D (new_AGEMA_signal_13902), .Q (new_AGEMA_signal_13903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6082 ( .C (clk), .D (new_AGEMA_signal_13906), .Q (new_AGEMA_signal_13907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6086 ( .C (clk), .D (new_AGEMA_signal_13910), .Q (new_AGEMA_signal_13911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6090 ( .C (clk), .D (new_AGEMA_signal_13914), .Q (new_AGEMA_signal_13915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6094 ( .C (clk), .D (new_AGEMA_signal_13918), .Q (new_AGEMA_signal_13919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6098 ( .C (clk), .D (new_AGEMA_signal_13922), .Q (new_AGEMA_signal_13923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6102 ( .C (clk), .D (new_AGEMA_signal_13926), .Q (new_AGEMA_signal_13927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6106 ( .C (clk), .D (new_AGEMA_signal_13930), .Q (new_AGEMA_signal_13931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6110 ( .C (clk), .D (new_AGEMA_signal_13934), .Q (new_AGEMA_signal_13935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6114 ( .C (clk), .D (new_AGEMA_signal_13938), .Q (new_AGEMA_signal_13939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6118 ( .C (clk), .D (new_AGEMA_signal_13942), .Q (new_AGEMA_signal_13943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6122 ( .C (clk), .D (new_AGEMA_signal_13946), .Q (new_AGEMA_signal_13947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6126 ( .C (clk), .D (new_AGEMA_signal_13950), .Q (new_AGEMA_signal_13951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6130 ( .C (clk), .D (new_AGEMA_signal_13954), .Q (new_AGEMA_signal_13955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6134 ( .C (clk), .D (new_AGEMA_signal_13958), .Q (new_AGEMA_signal_13959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6138 ( .C (clk), .D (new_AGEMA_signal_13962), .Q (new_AGEMA_signal_13963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6142 ( .C (clk), .D (new_AGEMA_signal_13966), .Q (new_AGEMA_signal_13967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6146 ( .C (clk), .D (new_AGEMA_signal_13970), .Q (new_AGEMA_signal_13971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6150 ( .C (clk), .D (new_AGEMA_signal_13974), .Q (new_AGEMA_signal_13975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6154 ( .C (clk), .D (new_AGEMA_signal_13978), .Q (new_AGEMA_signal_13979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6158 ( .C (clk), .D (new_AGEMA_signal_13982), .Q (new_AGEMA_signal_13983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6162 ( .C (clk), .D (new_AGEMA_signal_13986), .Q (new_AGEMA_signal_13987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6166 ( .C (clk), .D (new_AGEMA_signal_13990), .Q (new_AGEMA_signal_13991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6170 ( .C (clk), .D (new_AGEMA_signal_13994), .Q (new_AGEMA_signal_13995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6174 ( .C (clk), .D (new_AGEMA_signal_13998), .Q (new_AGEMA_signal_13999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6178 ( .C (clk), .D (new_AGEMA_signal_14002), .Q (new_AGEMA_signal_14003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6182 ( .C (clk), .D (new_AGEMA_signal_14006), .Q (new_AGEMA_signal_14007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6186 ( .C (clk), .D (new_AGEMA_signal_14010), .Q (new_AGEMA_signal_14011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6190 ( .C (clk), .D (new_AGEMA_signal_14014), .Q (new_AGEMA_signal_14015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6194 ( .C (clk), .D (new_AGEMA_signal_14018), .Q (new_AGEMA_signal_14019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6198 ( .C (clk), .D (new_AGEMA_signal_14022), .Q (new_AGEMA_signal_14023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6202 ( .C (clk), .D (new_AGEMA_signal_14026), .Q (new_AGEMA_signal_14027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6206 ( .C (clk), .D (new_AGEMA_signal_14030), .Q (new_AGEMA_signal_14031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6210 ( .C (clk), .D (new_AGEMA_signal_14034), .Q (new_AGEMA_signal_14035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6214 ( .C (clk), .D (new_AGEMA_signal_14038), .Q (new_AGEMA_signal_14039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6218 ( .C (clk), .D (new_AGEMA_signal_14042), .Q (new_AGEMA_signal_14043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6222 ( .C (clk), .D (new_AGEMA_signal_14046), .Q (new_AGEMA_signal_14047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6226 ( .C (clk), .D (new_AGEMA_signal_14050), .Q (new_AGEMA_signal_14051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6230 ( .C (clk), .D (new_AGEMA_signal_14054), .Q (new_AGEMA_signal_14055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6234 ( .C (clk), .D (new_AGEMA_signal_14058), .Q (new_AGEMA_signal_14059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6238 ( .C (clk), .D (new_AGEMA_signal_14062), .Q (new_AGEMA_signal_14063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6242 ( .C (clk), .D (new_AGEMA_signal_14066), .Q (new_AGEMA_signal_14067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6246 ( .C (clk), .D (new_AGEMA_signal_14070), .Q (new_AGEMA_signal_14071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6250 ( .C (clk), .D (new_AGEMA_signal_14074), .Q (new_AGEMA_signal_14075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6254 ( .C (clk), .D (new_AGEMA_signal_14078), .Q (new_AGEMA_signal_14079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6258 ( .C (clk), .D (new_AGEMA_signal_14082), .Q (new_AGEMA_signal_14083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6262 ( .C (clk), .D (new_AGEMA_signal_14086), .Q (new_AGEMA_signal_14087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6266 ( .C (clk), .D (new_AGEMA_signal_14090), .Q (new_AGEMA_signal_14091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6270 ( .C (clk), .D (new_AGEMA_signal_14094), .Q (new_AGEMA_signal_14095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6274 ( .C (clk), .D (new_AGEMA_signal_14098), .Q (new_AGEMA_signal_14099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6278 ( .C (clk), .D (new_AGEMA_signal_14102), .Q (new_AGEMA_signal_14103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6282 ( .C (clk), .D (new_AGEMA_signal_14106), .Q (new_AGEMA_signal_14107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6286 ( .C (clk), .D (new_AGEMA_signal_14110), .Q (new_AGEMA_signal_14111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6290 ( .C (clk), .D (new_AGEMA_signal_14114), .Q (new_AGEMA_signal_14115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6294 ( .C (clk), .D (new_AGEMA_signal_14118), .Q (new_AGEMA_signal_14119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6298 ( .C (clk), .D (new_AGEMA_signal_14122), .Q (new_AGEMA_signal_14123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6302 ( .C (clk), .D (new_AGEMA_signal_14126), .Q (new_AGEMA_signal_14127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6306 ( .C (clk), .D (new_AGEMA_signal_14130), .Q (new_AGEMA_signal_14131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6310 ( .C (clk), .D (new_AGEMA_signal_14134), .Q (new_AGEMA_signal_14135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6314 ( .C (clk), .D (new_AGEMA_signal_14138), .Q (new_AGEMA_signal_14139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6318 ( .C (clk), .D (new_AGEMA_signal_14142), .Q (new_AGEMA_signal_14143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6322 ( .C (clk), .D (new_AGEMA_signal_14146), .Q (new_AGEMA_signal_14147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6326 ( .C (clk), .D (new_AGEMA_signal_14150), .Q (new_AGEMA_signal_14151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6330 ( .C (clk), .D (new_AGEMA_signal_14154), .Q (new_AGEMA_signal_14155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6334 ( .C (clk), .D (new_AGEMA_signal_14158), .Q (new_AGEMA_signal_14159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6338 ( .C (clk), .D (new_AGEMA_signal_14162), .Q (new_AGEMA_signal_14163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6342 ( .C (clk), .D (new_AGEMA_signal_14166), .Q (new_AGEMA_signal_14167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6346 ( .C (clk), .D (new_AGEMA_signal_14170), .Q (new_AGEMA_signal_14171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6350 ( .C (clk), .D (new_AGEMA_signal_14174), .Q (new_AGEMA_signal_14175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6354 ( .C (clk), .D (new_AGEMA_signal_14178), .Q (new_AGEMA_signal_14179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6358 ( .C (clk), .D (new_AGEMA_signal_14182), .Q (new_AGEMA_signal_14183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6362 ( .C (clk), .D (new_AGEMA_signal_14186), .Q (new_AGEMA_signal_14187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6366 ( .C (clk), .D (new_AGEMA_signal_14190), .Q (new_AGEMA_signal_14191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6370 ( .C (clk), .D (new_AGEMA_signal_14194), .Q (new_AGEMA_signal_14195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6374 ( .C (clk), .D (new_AGEMA_signal_14198), .Q (new_AGEMA_signal_14199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6378 ( .C (clk), .D (new_AGEMA_signal_14202), .Q (new_AGEMA_signal_14203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6382 ( .C (clk), .D (new_AGEMA_signal_14206), .Q (new_AGEMA_signal_14207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6386 ( .C (clk), .D (new_AGEMA_signal_14210), .Q (new_AGEMA_signal_14211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6390 ( .C (clk), .D (new_AGEMA_signal_14214), .Q (new_AGEMA_signal_14215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6394 ( .C (clk), .D (new_AGEMA_signal_14218), .Q (new_AGEMA_signal_14219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6398 ( .C (clk), .D (new_AGEMA_signal_14222), .Q (new_AGEMA_signal_14223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6402 ( .C (clk), .D (new_AGEMA_signal_14226), .Q (new_AGEMA_signal_14227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6406 ( .C (clk), .D (new_AGEMA_signal_14230), .Q (new_AGEMA_signal_14231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6410 ( .C (clk), .D (new_AGEMA_signal_14234), .Q (new_AGEMA_signal_14235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6414 ( .C (clk), .D (new_AGEMA_signal_14238), .Q (new_AGEMA_signal_14239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6418 ( .C (clk), .D (new_AGEMA_signal_14242), .Q (new_AGEMA_signal_14243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6422 ( .C (clk), .D (new_AGEMA_signal_14246), .Q (new_AGEMA_signal_14247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6426 ( .C (clk), .D (new_AGEMA_signal_14250), .Q (new_AGEMA_signal_14251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6430 ( .C (clk), .D (new_AGEMA_signal_14254), .Q (new_AGEMA_signal_14255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6434 ( .C (clk), .D (new_AGEMA_signal_14258), .Q (new_AGEMA_signal_14259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6438 ( .C (clk), .D (new_AGEMA_signal_14262), .Q (new_AGEMA_signal_14263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6442 ( .C (clk), .D (new_AGEMA_signal_14266), .Q (new_AGEMA_signal_14267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6446 ( .C (clk), .D (new_AGEMA_signal_14270), .Q (new_AGEMA_signal_14271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6450 ( .C (clk), .D (new_AGEMA_signal_14274), .Q (new_AGEMA_signal_14275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6454 ( .C (clk), .D (new_AGEMA_signal_14278), .Q (new_AGEMA_signal_14279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6458 ( .C (clk), .D (new_AGEMA_signal_14282), .Q (new_AGEMA_signal_14283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6462 ( .C (clk), .D (new_AGEMA_signal_14286), .Q (new_AGEMA_signal_14287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6466 ( .C (clk), .D (new_AGEMA_signal_14290), .Q (new_AGEMA_signal_14291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6470 ( .C (clk), .D (new_AGEMA_signal_14294), .Q (new_AGEMA_signal_14295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6474 ( .C (clk), .D (new_AGEMA_signal_14298), .Q (new_AGEMA_signal_14299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6478 ( .C (clk), .D (new_AGEMA_signal_14302), .Q (new_AGEMA_signal_14303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6482 ( .C (clk), .D (new_AGEMA_signal_14306), .Q (new_AGEMA_signal_14307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6486 ( .C (clk), .D (new_AGEMA_signal_14310), .Q (new_AGEMA_signal_14311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6490 ( .C (clk), .D (new_AGEMA_signal_14314), .Q (new_AGEMA_signal_14315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6494 ( .C (clk), .D (new_AGEMA_signal_14318), .Q (new_AGEMA_signal_14319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6498 ( .C (clk), .D (new_AGEMA_signal_14322), .Q (new_AGEMA_signal_14323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6502 ( .C (clk), .D (new_AGEMA_signal_14326), .Q (new_AGEMA_signal_14327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6506 ( .C (clk), .D (new_AGEMA_signal_14330), .Q (new_AGEMA_signal_14331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6510 ( .C (clk), .D (new_AGEMA_signal_14334), .Q (new_AGEMA_signal_14335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6514 ( .C (clk), .D (new_AGEMA_signal_14338), .Q (new_AGEMA_signal_14339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6518 ( .C (clk), .D (new_AGEMA_signal_14342), .Q (new_AGEMA_signal_14343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6522 ( .C (clk), .D (new_AGEMA_signal_14346), .Q (new_AGEMA_signal_14347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6526 ( .C (clk), .D (new_AGEMA_signal_14350), .Q (new_AGEMA_signal_14351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6530 ( .C (clk), .D (new_AGEMA_signal_14354), .Q (new_AGEMA_signal_14355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6534 ( .C (clk), .D (new_AGEMA_signal_14358), .Q (new_AGEMA_signal_14359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6538 ( .C (clk), .D (new_AGEMA_signal_14362), .Q (new_AGEMA_signal_14363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6542 ( .C (clk), .D (new_AGEMA_signal_14366), .Q (new_AGEMA_signal_14367) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6546 ( .C (clk), .D (new_AGEMA_signal_14370), .Q (new_AGEMA_signal_14371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6550 ( .C (clk), .D (new_AGEMA_signal_14374), .Q (new_AGEMA_signal_14375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6554 ( .C (clk), .D (new_AGEMA_signal_14378), .Q (new_AGEMA_signal_14379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6558 ( .C (clk), .D (new_AGEMA_signal_14382), .Q (new_AGEMA_signal_14383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6562 ( .C (clk), .D (new_AGEMA_signal_14386), .Q (new_AGEMA_signal_14387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6566 ( .C (clk), .D (new_AGEMA_signal_14390), .Q (new_AGEMA_signal_14391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6570 ( .C (clk), .D (new_AGEMA_signal_14394), .Q (new_AGEMA_signal_14395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6574 ( .C (clk), .D (new_AGEMA_signal_14398), .Q (new_AGEMA_signal_14399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6578 ( .C (clk), .D (new_AGEMA_signal_14402), .Q (new_AGEMA_signal_14403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6582 ( .C (clk), .D (new_AGEMA_signal_14406), .Q (new_AGEMA_signal_14407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6586 ( .C (clk), .D (new_AGEMA_signal_14410), .Q (new_AGEMA_signal_14411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6590 ( .C (clk), .D (new_AGEMA_signal_14414), .Q (new_AGEMA_signal_14415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6594 ( .C (clk), .D (new_AGEMA_signal_14418), .Q (new_AGEMA_signal_14419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6598 ( .C (clk), .D (new_AGEMA_signal_14422), .Q (new_AGEMA_signal_14423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6602 ( .C (clk), .D (new_AGEMA_signal_14426), .Q (new_AGEMA_signal_14427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6606 ( .C (clk), .D (new_AGEMA_signal_14430), .Q (new_AGEMA_signal_14431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6610 ( .C (clk), .D (new_AGEMA_signal_14434), .Q (new_AGEMA_signal_14435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6614 ( .C (clk), .D (new_AGEMA_signal_14438), .Q (new_AGEMA_signal_14439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6618 ( .C (clk), .D (new_AGEMA_signal_14442), .Q (new_AGEMA_signal_14443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6622 ( .C (clk), .D (new_AGEMA_signal_14446), .Q (new_AGEMA_signal_14447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6626 ( .C (clk), .D (new_AGEMA_signal_14450), .Q (new_AGEMA_signal_14451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6630 ( .C (clk), .D (new_AGEMA_signal_14454), .Q (new_AGEMA_signal_14455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6634 ( .C (clk), .D (new_AGEMA_signal_14458), .Q (new_AGEMA_signal_14459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6638 ( .C (clk), .D (new_AGEMA_signal_14462), .Q (new_AGEMA_signal_14463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6642 ( .C (clk), .D (new_AGEMA_signal_14466), .Q (new_AGEMA_signal_14467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6646 ( .C (clk), .D (new_AGEMA_signal_14470), .Q (new_AGEMA_signal_14471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6650 ( .C (clk), .D (new_AGEMA_signal_14474), .Q (new_AGEMA_signal_14475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6654 ( .C (clk), .D (new_AGEMA_signal_14478), .Q (new_AGEMA_signal_14479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6658 ( .C (clk), .D (new_AGEMA_signal_14482), .Q (new_AGEMA_signal_14483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6662 ( .C (clk), .D (new_AGEMA_signal_14486), .Q (new_AGEMA_signal_14487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6666 ( .C (clk), .D (new_AGEMA_signal_14490), .Q (new_AGEMA_signal_14491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6670 ( .C (clk), .D (new_AGEMA_signal_14494), .Q (new_AGEMA_signal_14495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6674 ( .C (clk), .D (new_AGEMA_signal_14498), .Q (new_AGEMA_signal_14499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6678 ( .C (clk), .D (new_AGEMA_signal_14502), .Q (new_AGEMA_signal_14503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6682 ( .C (clk), .D (new_AGEMA_signal_14506), .Q (new_AGEMA_signal_14507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6686 ( .C (clk), .D (new_AGEMA_signal_14510), .Q (new_AGEMA_signal_14511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6690 ( .C (clk), .D (new_AGEMA_signal_14514), .Q (new_AGEMA_signal_14515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6694 ( .C (clk), .D (new_AGEMA_signal_14518), .Q (new_AGEMA_signal_14519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6698 ( .C (clk), .D (new_AGEMA_signal_14522), .Q (new_AGEMA_signal_14523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6702 ( .C (clk), .D (new_AGEMA_signal_14526), .Q (new_AGEMA_signal_14527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6706 ( .C (clk), .D (new_AGEMA_signal_14530), .Q (new_AGEMA_signal_14531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6710 ( .C (clk), .D (new_AGEMA_signal_14534), .Q (new_AGEMA_signal_14535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6714 ( .C (clk), .D (new_AGEMA_signal_14538), .Q (new_AGEMA_signal_14539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6718 ( .C (clk), .D (new_AGEMA_signal_14542), .Q (new_AGEMA_signal_14543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6722 ( .C (clk), .D (new_AGEMA_signal_14546), .Q (new_AGEMA_signal_14547) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6726 ( .C (clk), .D (new_AGEMA_signal_14550), .Q (new_AGEMA_signal_14551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6730 ( .C (clk), .D (new_AGEMA_signal_14554), .Q (new_AGEMA_signal_14555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6734 ( .C (clk), .D (new_AGEMA_signal_14558), .Q (new_AGEMA_signal_14559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6738 ( .C (clk), .D (new_AGEMA_signal_14562), .Q (new_AGEMA_signal_14563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6742 ( .C (clk), .D (new_AGEMA_signal_14566), .Q (new_AGEMA_signal_14567) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6746 ( .C (clk), .D (new_AGEMA_signal_14570), .Q (new_AGEMA_signal_14571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6750 ( .C (clk), .D (new_AGEMA_signal_14574), .Q (new_AGEMA_signal_14575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6754 ( .C (clk), .D (new_AGEMA_signal_14578), .Q (new_AGEMA_signal_14579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6758 ( .C (clk), .D (new_AGEMA_signal_14582), .Q (new_AGEMA_signal_14583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6762 ( .C (clk), .D (new_AGEMA_signal_14586), .Q (new_AGEMA_signal_14587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6766 ( .C (clk), .D (new_AGEMA_signal_14590), .Q (new_AGEMA_signal_14591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6770 ( .C (clk), .D (new_AGEMA_signal_14594), .Q (new_AGEMA_signal_14595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6774 ( .C (clk), .D (new_AGEMA_signal_14598), .Q (new_AGEMA_signal_14599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6778 ( .C (clk), .D (new_AGEMA_signal_14602), .Q (new_AGEMA_signal_14603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6782 ( .C (clk), .D (new_AGEMA_signal_14606), .Q (new_AGEMA_signal_14607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6786 ( .C (clk), .D (new_AGEMA_signal_14610), .Q (new_AGEMA_signal_14611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6790 ( .C (clk), .D (new_AGEMA_signal_14614), .Q (new_AGEMA_signal_14615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6794 ( .C (clk), .D (new_AGEMA_signal_14618), .Q (new_AGEMA_signal_14619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6798 ( .C (clk), .D (new_AGEMA_signal_14622), .Q (new_AGEMA_signal_14623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6802 ( .C (clk), .D (new_AGEMA_signal_14626), .Q (new_AGEMA_signal_14627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6806 ( .C (clk), .D (new_AGEMA_signal_14630), .Q (new_AGEMA_signal_14631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6810 ( .C (clk), .D (new_AGEMA_signal_14634), .Q (new_AGEMA_signal_14635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6814 ( .C (clk), .D (new_AGEMA_signal_14638), .Q (new_AGEMA_signal_14639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6818 ( .C (clk), .D (new_AGEMA_signal_14642), .Q (new_AGEMA_signal_14643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6822 ( .C (clk), .D (new_AGEMA_signal_14646), .Q (new_AGEMA_signal_14647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6826 ( .C (clk), .D (new_AGEMA_signal_14650), .Q (new_AGEMA_signal_14651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6830 ( .C (clk), .D (new_AGEMA_signal_14654), .Q (new_AGEMA_signal_14655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6834 ( .C (clk), .D (new_AGEMA_signal_14658), .Q (new_AGEMA_signal_14659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6838 ( .C (clk), .D (new_AGEMA_signal_14662), .Q (new_AGEMA_signal_14663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6842 ( .C (clk), .D (new_AGEMA_signal_14666), .Q (new_AGEMA_signal_14667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6846 ( .C (clk), .D (new_AGEMA_signal_14670), .Q (new_AGEMA_signal_14671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6850 ( .C (clk), .D (new_AGEMA_signal_14674), .Q (new_AGEMA_signal_14675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6854 ( .C (clk), .D (new_AGEMA_signal_14678), .Q (new_AGEMA_signal_14679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6858 ( .C (clk), .D (new_AGEMA_signal_14682), .Q (new_AGEMA_signal_14683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6862 ( .C (clk), .D (new_AGEMA_signal_14686), .Q (new_AGEMA_signal_14687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6866 ( .C (clk), .D (new_AGEMA_signal_14690), .Q (new_AGEMA_signal_14691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6870 ( .C (clk), .D (new_AGEMA_signal_14694), .Q (new_AGEMA_signal_14695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6874 ( .C (clk), .D (new_AGEMA_signal_14698), .Q (new_AGEMA_signal_14699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6878 ( .C (clk), .D (new_AGEMA_signal_14702), .Q (new_AGEMA_signal_14703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6882 ( .C (clk), .D (new_AGEMA_signal_14706), .Q (new_AGEMA_signal_14707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6886 ( .C (clk), .D (new_AGEMA_signal_14710), .Q (new_AGEMA_signal_14711) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6890 ( .C (clk), .D (new_AGEMA_signal_14714), .Q (new_AGEMA_signal_14715) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6894 ( .C (clk), .D (new_AGEMA_signal_14718), .Q (new_AGEMA_signal_14719) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6898 ( .C (clk), .D (new_AGEMA_signal_14722), .Q (new_AGEMA_signal_14723) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6902 ( .C (clk), .D (new_AGEMA_signal_14726), .Q (new_AGEMA_signal_14727) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6906 ( .C (clk), .D (new_AGEMA_signal_14730), .Q (new_AGEMA_signal_14731) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6910 ( .C (clk), .D (new_AGEMA_signal_14734), .Q (new_AGEMA_signal_14735) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6914 ( .C (clk), .D (new_AGEMA_signal_14738), .Q (new_AGEMA_signal_14739) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6918 ( .C (clk), .D (new_AGEMA_signal_14742), .Q (new_AGEMA_signal_14743) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6922 ( .C (clk), .D (new_AGEMA_signal_14746), .Q (new_AGEMA_signal_14747) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6926 ( .C (clk), .D (new_AGEMA_signal_14750), .Q (new_AGEMA_signal_14751) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6930 ( .C (clk), .D (new_AGEMA_signal_14754), .Q (new_AGEMA_signal_14755) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6934 ( .C (clk), .D (new_AGEMA_signal_14758), .Q (new_AGEMA_signal_14759) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6938 ( .C (clk), .D (new_AGEMA_signal_14762), .Q (new_AGEMA_signal_14763) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6942 ( .C (clk), .D (new_AGEMA_signal_14766), .Q (new_AGEMA_signal_14767) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6946 ( .C (clk), .D (new_AGEMA_signal_14770), .Q (new_AGEMA_signal_14771) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6950 ( .C (clk), .D (new_AGEMA_signal_14774), .Q (new_AGEMA_signal_14775) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6954 ( .C (clk), .D (new_AGEMA_signal_14778), .Q (new_AGEMA_signal_14779) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6958 ( .C (clk), .D (new_AGEMA_signal_14782), .Q (new_AGEMA_signal_14783) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6962 ( .C (clk), .D (new_AGEMA_signal_14786), .Q (new_AGEMA_signal_14787) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6966 ( .C (clk), .D (new_AGEMA_signal_14790), .Q (new_AGEMA_signal_14791) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6970 ( .C (clk), .D (new_AGEMA_signal_14794), .Q (new_AGEMA_signal_14795) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6974 ( .C (clk), .D (new_AGEMA_signal_14798), .Q (new_AGEMA_signal_14799) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6978 ( .C (clk), .D (new_AGEMA_signal_14802), .Q (new_AGEMA_signal_14803) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6982 ( .C (clk), .D (new_AGEMA_signal_14806), .Q (new_AGEMA_signal_14807) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6986 ( .C (clk), .D (new_AGEMA_signal_14810), .Q (new_AGEMA_signal_14811) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6990 ( .C (clk), .D (new_AGEMA_signal_14814), .Q (new_AGEMA_signal_14815) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6994 ( .C (clk), .D (new_AGEMA_signal_14818), .Q (new_AGEMA_signal_14819) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6998 ( .C (clk), .D (new_AGEMA_signal_14822), .Q (new_AGEMA_signal_14823) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7002 ( .C (clk), .D (new_AGEMA_signal_14826), .Q (new_AGEMA_signal_14827) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7006 ( .C (clk), .D (new_AGEMA_signal_14830), .Q (new_AGEMA_signal_14831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7010 ( .C (clk), .D (new_AGEMA_signal_14834), .Q (new_AGEMA_signal_14835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7014 ( .C (clk), .D (new_AGEMA_signal_14838), .Q (new_AGEMA_signal_14839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7018 ( .C (clk), .D (new_AGEMA_signal_14842), .Q (new_AGEMA_signal_14843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7022 ( .C (clk), .D (new_AGEMA_signal_14846), .Q (new_AGEMA_signal_14847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7026 ( .C (clk), .D (new_AGEMA_signal_14850), .Q (new_AGEMA_signal_14851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7030 ( .C (clk), .D (new_AGEMA_signal_14854), .Q (new_AGEMA_signal_14855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7034 ( .C (clk), .D (new_AGEMA_signal_14858), .Q (new_AGEMA_signal_14859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7038 ( .C (clk), .D (new_AGEMA_signal_14862), .Q (new_AGEMA_signal_14863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7042 ( .C (clk), .D (new_AGEMA_signal_14866), .Q (new_AGEMA_signal_14867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7046 ( .C (clk), .D (new_AGEMA_signal_14870), .Q (new_AGEMA_signal_14871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7050 ( .C (clk), .D (new_AGEMA_signal_14874), .Q (new_AGEMA_signal_14875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7054 ( .C (clk), .D (new_AGEMA_signal_14878), .Q (new_AGEMA_signal_14879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7058 ( .C (clk), .D (new_AGEMA_signal_14882), .Q (new_AGEMA_signal_14883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7062 ( .C (clk), .D (new_AGEMA_signal_14886), .Q (new_AGEMA_signal_14887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7066 ( .C (clk), .D (new_AGEMA_signal_14890), .Q (new_AGEMA_signal_14891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7070 ( .C (clk), .D (new_AGEMA_signal_14894), .Q (new_AGEMA_signal_14895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7074 ( .C (clk), .D (new_AGEMA_signal_14898), .Q (new_AGEMA_signal_14899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7078 ( .C (clk), .D (new_AGEMA_signal_14902), .Q (new_AGEMA_signal_14903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7082 ( .C (clk), .D (new_AGEMA_signal_14906), .Q (new_AGEMA_signal_14907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7086 ( .C (clk), .D (new_AGEMA_signal_14910), .Q (new_AGEMA_signal_14911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7090 ( .C (clk), .D (new_AGEMA_signal_14914), .Q (new_AGEMA_signal_14915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7094 ( .C (clk), .D (new_AGEMA_signal_14918), .Q (new_AGEMA_signal_14919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7098 ( .C (clk), .D (new_AGEMA_signal_14922), .Q (new_AGEMA_signal_14923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7102 ( .C (clk), .D (new_AGEMA_signal_14926), .Q (new_AGEMA_signal_14927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7106 ( .C (clk), .D (new_AGEMA_signal_14930), .Q (new_AGEMA_signal_14931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7110 ( .C (clk), .D (new_AGEMA_signal_14934), .Q (new_AGEMA_signal_14935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7114 ( .C (clk), .D (new_AGEMA_signal_14938), .Q (new_AGEMA_signal_14939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7118 ( .C (clk), .D (new_AGEMA_signal_14942), .Q (new_AGEMA_signal_14943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7122 ( .C (clk), .D (new_AGEMA_signal_14946), .Q (new_AGEMA_signal_14947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7126 ( .C (clk), .D (new_AGEMA_signal_14950), .Q (new_AGEMA_signal_14951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7130 ( .C (clk), .D (new_AGEMA_signal_14954), .Q (new_AGEMA_signal_14955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7134 ( .C (clk), .D (new_AGEMA_signal_14958), .Q (new_AGEMA_signal_14959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7138 ( .C (clk), .D (new_AGEMA_signal_14962), .Q (new_AGEMA_signal_14963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7142 ( .C (clk), .D (new_AGEMA_signal_14966), .Q (new_AGEMA_signal_14967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7146 ( .C (clk), .D (new_AGEMA_signal_14970), .Q (new_AGEMA_signal_14971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7150 ( .C (clk), .D (new_AGEMA_signal_14974), .Q (new_AGEMA_signal_14975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7154 ( .C (clk), .D (new_AGEMA_signal_14978), .Q (new_AGEMA_signal_14979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7158 ( .C (clk), .D (new_AGEMA_signal_14982), .Q (new_AGEMA_signal_14983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7162 ( .C (clk), .D (new_AGEMA_signal_14986), .Q (new_AGEMA_signal_14987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7166 ( .C (clk), .D (new_AGEMA_signal_14990), .Q (new_AGEMA_signal_14991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7170 ( .C (clk), .D (new_AGEMA_signal_14994), .Q (new_AGEMA_signal_14995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7174 ( .C (clk), .D (new_AGEMA_signal_14998), .Q (new_AGEMA_signal_14999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7178 ( .C (clk), .D (new_AGEMA_signal_15002), .Q (new_AGEMA_signal_15003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7182 ( .C (clk), .D (new_AGEMA_signal_15006), .Q (new_AGEMA_signal_15007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7186 ( .C (clk), .D (new_AGEMA_signal_15010), .Q (new_AGEMA_signal_15011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7190 ( .C (clk), .D (new_AGEMA_signal_15014), .Q (new_AGEMA_signal_15015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7194 ( .C (clk), .D (new_AGEMA_signal_15018), .Q (new_AGEMA_signal_15019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7198 ( .C (clk), .D (new_AGEMA_signal_15022), .Q (new_AGEMA_signal_15023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7202 ( .C (clk), .D (new_AGEMA_signal_15026), .Q (new_AGEMA_signal_15027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7206 ( .C (clk), .D (new_AGEMA_signal_15030), .Q (new_AGEMA_signal_15031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7210 ( .C (clk), .D (new_AGEMA_signal_15034), .Q (new_AGEMA_signal_15035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7214 ( .C (clk), .D (new_AGEMA_signal_15038), .Q (new_AGEMA_signal_15039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7218 ( .C (clk), .D (new_AGEMA_signal_15042), .Q (new_AGEMA_signal_15043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7222 ( .C (clk), .D (new_AGEMA_signal_15046), .Q (new_AGEMA_signal_15047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7226 ( .C (clk), .D (new_AGEMA_signal_15050), .Q (new_AGEMA_signal_15051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7230 ( .C (clk), .D (new_AGEMA_signal_15054), .Q (new_AGEMA_signal_15055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7234 ( .C (clk), .D (new_AGEMA_signal_15058), .Q (new_AGEMA_signal_15059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7238 ( .C (clk), .D (new_AGEMA_signal_15062), .Q (new_AGEMA_signal_15063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7242 ( .C (clk), .D (new_AGEMA_signal_15066), .Q (new_AGEMA_signal_15067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7246 ( .C (clk), .D (new_AGEMA_signal_15070), .Q (new_AGEMA_signal_15071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7250 ( .C (clk), .D (new_AGEMA_signal_15074), .Q (new_AGEMA_signal_15075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7254 ( .C (clk), .D (new_AGEMA_signal_15078), .Q (new_AGEMA_signal_15079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7258 ( .C (clk), .D (new_AGEMA_signal_15082), .Q (new_AGEMA_signal_15083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7262 ( .C (clk), .D (new_AGEMA_signal_15086), .Q (new_AGEMA_signal_15087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7266 ( .C (clk), .D (new_AGEMA_signal_15090), .Q (new_AGEMA_signal_15091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7270 ( .C (clk), .D (new_AGEMA_signal_15094), .Q (new_AGEMA_signal_15095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7274 ( .C (clk), .D (new_AGEMA_signal_15098), .Q (new_AGEMA_signal_15099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7278 ( .C (clk), .D (new_AGEMA_signal_15102), .Q (new_AGEMA_signal_15103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7282 ( .C (clk), .D (new_AGEMA_signal_15106), .Q (new_AGEMA_signal_15107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7286 ( .C (clk), .D (new_AGEMA_signal_15110), .Q (new_AGEMA_signal_15111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7290 ( .C (clk), .D (new_AGEMA_signal_15114), .Q (new_AGEMA_signal_15115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7294 ( .C (clk), .D (new_AGEMA_signal_15118), .Q (new_AGEMA_signal_15119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7298 ( .C (clk), .D (new_AGEMA_signal_15122), .Q (new_AGEMA_signal_15123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7302 ( .C (clk), .D (new_AGEMA_signal_15126), .Q (new_AGEMA_signal_15127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7306 ( .C (clk), .D (new_AGEMA_signal_15130), .Q (new_AGEMA_signal_15131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7310 ( .C (clk), .D (new_AGEMA_signal_15134), .Q (new_AGEMA_signal_15135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7314 ( .C (clk), .D (new_AGEMA_signal_15138), .Q (new_AGEMA_signal_15139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7318 ( .C (clk), .D (new_AGEMA_signal_15142), .Q (new_AGEMA_signal_15143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7322 ( .C (clk), .D (new_AGEMA_signal_15146), .Q (new_AGEMA_signal_15147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7326 ( .C (clk), .D (new_AGEMA_signal_15150), .Q (new_AGEMA_signal_15151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7330 ( .C (clk), .D (new_AGEMA_signal_15154), .Q (new_AGEMA_signal_15155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7334 ( .C (clk), .D (new_AGEMA_signal_15158), .Q (new_AGEMA_signal_15159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7338 ( .C (clk), .D (new_AGEMA_signal_15162), .Q (new_AGEMA_signal_15163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7342 ( .C (clk), .D (new_AGEMA_signal_15166), .Q (new_AGEMA_signal_15167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7346 ( .C (clk), .D (new_AGEMA_signal_15170), .Q (new_AGEMA_signal_15171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7350 ( .C (clk), .D (new_AGEMA_signal_15174), .Q (new_AGEMA_signal_15175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7354 ( .C (clk), .D (new_AGEMA_signal_15178), .Q (new_AGEMA_signal_15179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7358 ( .C (clk), .D (new_AGEMA_signal_15182), .Q (new_AGEMA_signal_15183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7362 ( .C (clk), .D (new_AGEMA_signal_15186), .Q (new_AGEMA_signal_15187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7366 ( .C (clk), .D (new_AGEMA_signal_15190), .Q (new_AGEMA_signal_15191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7370 ( .C (clk), .D (new_AGEMA_signal_15194), .Q (new_AGEMA_signal_15195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7374 ( .C (clk), .D (new_AGEMA_signal_15198), .Q (new_AGEMA_signal_15199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7378 ( .C (clk), .D (new_AGEMA_signal_15202), .Q (new_AGEMA_signal_15203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7382 ( .C (clk), .D (new_AGEMA_signal_15206), .Q (new_AGEMA_signal_15207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7386 ( .C (clk), .D (new_AGEMA_signal_15210), .Q (new_AGEMA_signal_15211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7390 ( .C (clk), .D (new_AGEMA_signal_15214), .Q (new_AGEMA_signal_15215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7394 ( .C (clk), .D (new_AGEMA_signal_15218), .Q (new_AGEMA_signal_15219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7398 ( .C (clk), .D (new_AGEMA_signal_15222), .Q (new_AGEMA_signal_15223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7402 ( .C (clk), .D (new_AGEMA_signal_15226), .Q (new_AGEMA_signal_15227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7406 ( .C (clk), .D (new_AGEMA_signal_15230), .Q (new_AGEMA_signal_15231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7410 ( .C (clk), .D (new_AGEMA_signal_15234), .Q (new_AGEMA_signal_15235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7414 ( .C (clk), .D (new_AGEMA_signal_15238), .Q (new_AGEMA_signal_15239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7418 ( .C (clk), .D (new_AGEMA_signal_15242), .Q (new_AGEMA_signal_15243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7422 ( .C (clk), .D (new_AGEMA_signal_15246), .Q (new_AGEMA_signal_15247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7426 ( .C (clk), .D (new_AGEMA_signal_15250), .Q (new_AGEMA_signal_15251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7430 ( .C (clk), .D (new_AGEMA_signal_15254), .Q (new_AGEMA_signal_15255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7434 ( .C (clk), .D (new_AGEMA_signal_15258), .Q (new_AGEMA_signal_15259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7438 ( .C (clk), .D (new_AGEMA_signal_15262), .Q (new_AGEMA_signal_15263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7442 ( .C (clk), .D (new_AGEMA_signal_15266), .Q (new_AGEMA_signal_15267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7446 ( .C (clk), .D (new_AGEMA_signal_15270), .Q (new_AGEMA_signal_15271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7450 ( .C (clk), .D (new_AGEMA_signal_15274), .Q (new_AGEMA_signal_15275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7454 ( .C (clk), .D (new_AGEMA_signal_15278), .Q (new_AGEMA_signal_15279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7458 ( .C (clk), .D (new_AGEMA_signal_15282), .Q (new_AGEMA_signal_15283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7462 ( .C (clk), .D (new_AGEMA_signal_15286), .Q (new_AGEMA_signal_15287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7466 ( .C (clk), .D (new_AGEMA_signal_15290), .Q (new_AGEMA_signal_15291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7470 ( .C (clk), .D (new_AGEMA_signal_15294), .Q (new_AGEMA_signal_15295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7474 ( .C (clk), .D (new_AGEMA_signal_15298), .Q (new_AGEMA_signal_15299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7478 ( .C (clk), .D (new_AGEMA_signal_15302), .Q (new_AGEMA_signal_15303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7482 ( .C (clk), .D (new_AGEMA_signal_15306), .Q (new_AGEMA_signal_15307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7486 ( .C (clk), .D (new_AGEMA_signal_15310), .Q (new_AGEMA_signal_15311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7490 ( .C (clk), .D (new_AGEMA_signal_15314), .Q (new_AGEMA_signal_15315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7494 ( .C (clk), .D (new_AGEMA_signal_15318), .Q (new_AGEMA_signal_15319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7498 ( .C (clk), .D (new_AGEMA_signal_15322), .Q (new_AGEMA_signal_15323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7502 ( .C (clk), .D (new_AGEMA_signal_15326), .Q (new_AGEMA_signal_15327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7506 ( .C (clk), .D (new_AGEMA_signal_15330), .Q (new_AGEMA_signal_15331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7510 ( .C (clk), .D (new_AGEMA_signal_15334), .Q (new_AGEMA_signal_15335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7514 ( .C (clk), .D (new_AGEMA_signal_15338), .Q (new_AGEMA_signal_15339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7518 ( .C (clk), .D (new_AGEMA_signal_15342), .Q (new_AGEMA_signal_15343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7522 ( .C (clk), .D (new_AGEMA_signal_15346), .Q (new_AGEMA_signal_15347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7526 ( .C (clk), .D (new_AGEMA_signal_15350), .Q (new_AGEMA_signal_15351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7530 ( .C (clk), .D (new_AGEMA_signal_15354), .Q (new_AGEMA_signal_15355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7534 ( .C (clk), .D (new_AGEMA_signal_15358), .Q (new_AGEMA_signal_15359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7538 ( .C (clk), .D (new_AGEMA_signal_15362), .Q (new_AGEMA_signal_15363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7542 ( .C (clk), .D (new_AGEMA_signal_15366), .Q (new_AGEMA_signal_15367) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7546 ( .C (clk), .D (new_AGEMA_signal_15370), .Q (new_AGEMA_signal_15371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7550 ( .C (clk), .D (new_AGEMA_signal_15374), .Q (new_AGEMA_signal_15375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7554 ( .C (clk), .D (new_AGEMA_signal_15378), .Q (new_AGEMA_signal_15379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7558 ( .C (clk), .D (new_AGEMA_signal_15382), .Q (new_AGEMA_signal_15383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7562 ( .C (clk), .D (new_AGEMA_signal_15386), .Q (new_AGEMA_signal_15387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7566 ( .C (clk), .D (new_AGEMA_signal_15390), .Q (new_AGEMA_signal_15391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7570 ( .C (clk), .D (new_AGEMA_signal_15394), .Q (new_AGEMA_signal_15395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7574 ( .C (clk), .D (new_AGEMA_signal_15398), .Q (new_AGEMA_signal_15399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7578 ( .C (clk), .D (new_AGEMA_signal_15402), .Q (new_AGEMA_signal_15403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7582 ( .C (clk), .D (new_AGEMA_signal_15406), .Q (new_AGEMA_signal_15407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7586 ( .C (clk), .D (new_AGEMA_signal_15410), .Q (new_AGEMA_signal_15411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7590 ( .C (clk), .D (new_AGEMA_signal_15414), .Q (new_AGEMA_signal_15415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7594 ( .C (clk), .D (new_AGEMA_signal_15418), .Q (new_AGEMA_signal_15419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7598 ( .C (clk), .D (new_AGEMA_signal_15422), .Q (new_AGEMA_signal_15423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7602 ( .C (clk), .D (new_AGEMA_signal_15426), .Q (new_AGEMA_signal_15427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7606 ( .C (clk), .D (new_AGEMA_signal_15430), .Q (new_AGEMA_signal_15431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7610 ( .C (clk), .D (new_AGEMA_signal_15434), .Q (new_AGEMA_signal_15435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7614 ( .C (clk), .D (new_AGEMA_signal_15438), .Q (new_AGEMA_signal_15439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7618 ( .C (clk), .D (new_AGEMA_signal_15442), .Q (new_AGEMA_signal_15443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7622 ( .C (clk), .D (new_AGEMA_signal_15446), .Q (new_AGEMA_signal_15447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7626 ( .C (clk), .D (new_AGEMA_signal_15450), .Q (new_AGEMA_signal_15451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7630 ( .C (clk), .D (new_AGEMA_signal_15454), .Q (new_AGEMA_signal_15455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7634 ( .C (clk), .D (new_AGEMA_signal_15458), .Q (new_AGEMA_signal_15459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7638 ( .C (clk), .D (new_AGEMA_signal_15462), .Q (new_AGEMA_signal_15463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7642 ( .C (clk), .D (new_AGEMA_signal_15466), .Q (new_AGEMA_signal_15467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7646 ( .C (clk), .D (new_AGEMA_signal_15470), .Q (new_AGEMA_signal_15471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7650 ( .C (clk), .D (new_AGEMA_signal_15474), .Q (new_AGEMA_signal_15475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7654 ( .C (clk), .D (new_AGEMA_signal_15478), .Q (new_AGEMA_signal_15479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7658 ( .C (clk), .D (new_AGEMA_signal_15482), .Q (new_AGEMA_signal_15483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7662 ( .C (clk), .D (new_AGEMA_signal_15486), .Q (new_AGEMA_signal_15487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7666 ( .C (clk), .D (new_AGEMA_signal_15490), .Q (new_AGEMA_signal_15491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7670 ( .C (clk), .D (new_AGEMA_signal_15494), .Q (new_AGEMA_signal_15495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7674 ( .C (clk), .D (new_AGEMA_signal_15498), .Q (new_AGEMA_signal_15499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7678 ( .C (clk), .D (new_AGEMA_signal_15502), .Q (new_AGEMA_signal_15503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7682 ( .C (clk), .D (new_AGEMA_signal_15506), .Q (new_AGEMA_signal_15507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7686 ( .C (clk), .D (new_AGEMA_signal_15510), .Q (new_AGEMA_signal_15511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7690 ( .C (clk), .D (new_AGEMA_signal_15514), .Q (new_AGEMA_signal_15515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7694 ( .C (clk), .D (new_AGEMA_signal_15518), .Q (new_AGEMA_signal_15519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7698 ( .C (clk), .D (new_AGEMA_signal_15522), .Q (new_AGEMA_signal_15523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7702 ( .C (clk), .D (new_AGEMA_signal_15526), .Q (new_AGEMA_signal_15527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7706 ( .C (clk), .D (new_AGEMA_signal_15530), .Q (new_AGEMA_signal_15531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7710 ( .C (clk), .D (new_AGEMA_signal_15534), .Q (new_AGEMA_signal_15535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7714 ( .C (clk), .D (new_AGEMA_signal_15538), .Q (new_AGEMA_signal_15539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7718 ( .C (clk), .D (new_AGEMA_signal_15542), .Q (new_AGEMA_signal_15543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7722 ( .C (clk), .D (new_AGEMA_signal_15546), .Q (new_AGEMA_signal_15547) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7726 ( .C (clk), .D (new_AGEMA_signal_15550), .Q (new_AGEMA_signal_15551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7730 ( .C (clk), .D (new_AGEMA_signal_15554), .Q (new_AGEMA_signal_15555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7734 ( .C (clk), .D (new_AGEMA_signal_15558), .Q (new_AGEMA_signal_15559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7738 ( .C (clk), .D (new_AGEMA_signal_15562), .Q (new_AGEMA_signal_15563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7742 ( .C (clk), .D (new_AGEMA_signal_15566), .Q (new_AGEMA_signal_15567) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7746 ( .C (clk), .D (new_AGEMA_signal_15570), .Q (new_AGEMA_signal_15571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7750 ( .C (clk), .D (new_AGEMA_signal_15574), .Q (new_AGEMA_signal_15575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7754 ( .C (clk), .D (new_AGEMA_signal_15578), .Q (new_AGEMA_signal_15579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7758 ( .C (clk), .D (new_AGEMA_signal_15582), .Q (new_AGEMA_signal_15583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7762 ( .C (clk), .D (new_AGEMA_signal_15586), .Q (new_AGEMA_signal_15587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7766 ( .C (clk), .D (new_AGEMA_signal_15590), .Q (new_AGEMA_signal_15591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7770 ( .C (clk), .D (new_AGEMA_signal_15594), .Q (new_AGEMA_signal_15595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7774 ( .C (clk), .D (new_AGEMA_signal_15598), .Q (new_AGEMA_signal_15599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7778 ( .C (clk), .D (new_AGEMA_signal_15602), .Q (new_AGEMA_signal_15603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7782 ( .C (clk), .D (new_AGEMA_signal_15606), .Q (new_AGEMA_signal_15607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7786 ( .C (clk), .D (new_AGEMA_signal_15610), .Q (new_AGEMA_signal_15611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7790 ( .C (clk), .D (new_AGEMA_signal_15614), .Q (new_AGEMA_signal_15615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7794 ( .C (clk), .D (new_AGEMA_signal_15618), .Q (new_AGEMA_signal_15619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7798 ( .C (clk), .D (new_AGEMA_signal_15622), .Q (new_AGEMA_signal_15623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7802 ( .C (clk), .D (new_AGEMA_signal_15626), .Q (new_AGEMA_signal_15627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7806 ( .C (clk), .D (new_AGEMA_signal_15630), .Q (new_AGEMA_signal_15631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7810 ( .C (clk), .D (new_AGEMA_signal_15634), .Q (new_AGEMA_signal_15635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7814 ( .C (clk), .D (new_AGEMA_signal_15638), .Q (new_AGEMA_signal_15639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7818 ( .C (clk), .D (new_AGEMA_signal_15642), .Q (new_AGEMA_signal_15643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7822 ( .C (clk), .D (new_AGEMA_signal_15646), .Q (new_AGEMA_signal_15647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7826 ( .C (clk), .D (new_AGEMA_signal_15650), .Q (new_AGEMA_signal_15651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7830 ( .C (clk), .D (new_AGEMA_signal_15654), .Q (new_AGEMA_signal_15655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7834 ( .C (clk), .D (new_AGEMA_signal_15658), .Q (new_AGEMA_signal_15659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7838 ( .C (clk), .D (new_AGEMA_signal_15662), .Q (new_AGEMA_signal_15663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7842 ( .C (clk), .D (new_AGEMA_signal_15666), .Q (new_AGEMA_signal_15667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7846 ( .C (clk), .D (new_AGEMA_signal_15670), .Q (new_AGEMA_signal_15671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7850 ( .C (clk), .D (new_AGEMA_signal_15674), .Q (new_AGEMA_signal_15675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7854 ( .C (clk), .D (new_AGEMA_signal_15678), .Q (new_AGEMA_signal_15679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7858 ( .C (clk), .D (new_AGEMA_signal_15682), .Q (new_AGEMA_signal_15683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7862 ( .C (clk), .D (new_AGEMA_signal_15686), .Q (new_AGEMA_signal_15687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7866 ( .C (clk), .D (new_AGEMA_signal_15690), .Q (new_AGEMA_signal_15691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7870 ( .C (clk), .D (new_AGEMA_signal_15694), .Q (new_AGEMA_signal_15695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7874 ( .C (clk), .D (new_AGEMA_signal_15698), .Q (new_AGEMA_signal_15699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7878 ( .C (clk), .D (new_AGEMA_signal_15702), .Q (new_AGEMA_signal_15703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7882 ( .C (clk), .D (new_AGEMA_signal_15706), .Q (new_AGEMA_signal_15707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7886 ( .C (clk), .D (new_AGEMA_signal_15710), .Q (new_AGEMA_signal_15711) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7890 ( .C (clk), .D (new_AGEMA_signal_15714), .Q (new_AGEMA_signal_15715) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7894 ( .C (clk), .D (new_AGEMA_signal_15718), .Q (new_AGEMA_signal_15719) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7898 ( .C (clk), .D (new_AGEMA_signal_15722), .Q (new_AGEMA_signal_15723) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7902 ( .C (clk), .D (new_AGEMA_signal_15726), .Q (new_AGEMA_signal_15727) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7906 ( .C (clk), .D (new_AGEMA_signal_15730), .Q (new_AGEMA_signal_15731) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7910 ( .C (clk), .D (new_AGEMA_signal_15734), .Q (new_AGEMA_signal_15735) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7914 ( .C (clk), .D (new_AGEMA_signal_15738), .Q (new_AGEMA_signal_15739) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7918 ( .C (clk), .D (new_AGEMA_signal_15742), .Q (new_AGEMA_signal_15743) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7922 ( .C (clk), .D (new_AGEMA_signal_15746), .Q (new_AGEMA_signal_15747) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7926 ( .C (clk), .D (new_AGEMA_signal_15750), .Q (new_AGEMA_signal_15751) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7930 ( .C (clk), .D (new_AGEMA_signal_15754), .Q (new_AGEMA_signal_15755) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7934 ( .C (clk), .D (new_AGEMA_signal_15758), .Q (new_AGEMA_signal_15759) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7938 ( .C (clk), .D (new_AGEMA_signal_15762), .Q (new_AGEMA_signal_15763) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7942 ( .C (clk), .D (new_AGEMA_signal_15766), .Q (new_AGEMA_signal_15767) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7946 ( .C (clk), .D (new_AGEMA_signal_15770), .Q (new_AGEMA_signal_15771) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7950 ( .C (clk), .D (new_AGEMA_signal_15774), .Q (new_AGEMA_signal_15775) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7954 ( .C (clk), .D (new_AGEMA_signal_15778), .Q (new_AGEMA_signal_15779) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7958 ( .C (clk), .D (new_AGEMA_signal_15782), .Q (new_AGEMA_signal_15783) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7962 ( .C (clk), .D (new_AGEMA_signal_15786), .Q (new_AGEMA_signal_15787) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7966 ( .C (clk), .D (new_AGEMA_signal_15790), .Q (new_AGEMA_signal_15791) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7970 ( .C (clk), .D (new_AGEMA_signal_15794), .Q (new_AGEMA_signal_15795) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7974 ( .C (clk), .D (new_AGEMA_signal_15798), .Q (new_AGEMA_signal_15799) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7978 ( .C (clk), .D (new_AGEMA_signal_15802), .Q (new_AGEMA_signal_15803) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7982 ( .C (clk), .D (new_AGEMA_signal_15806), .Q (new_AGEMA_signal_15807) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7986 ( .C (clk), .D (new_AGEMA_signal_15810), .Q (new_AGEMA_signal_15811) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7990 ( .C (clk), .D (new_AGEMA_signal_15814), .Q (new_AGEMA_signal_15815) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7994 ( .C (clk), .D (new_AGEMA_signal_15818), .Q (new_AGEMA_signal_15819) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7998 ( .C (clk), .D (new_AGEMA_signal_15822), .Q (new_AGEMA_signal_15823) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8002 ( .C (clk), .D (new_AGEMA_signal_15826), .Q (new_AGEMA_signal_15827) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8006 ( .C (clk), .D (new_AGEMA_signal_15830), .Q (new_AGEMA_signal_15831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8010 ( .C (clk), .D (new_AGEMA_signal_15834), .Q (new_AGEMA_signal_15835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8014 ( .C (clk), .D (new_AGEMA_signal_15838), .Q (new_AGEMA_signal_15839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8018 ( .C (clk), .D (new_AGEMA_signal_15842), .Q (new_AGEMA_signal_15843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8022 ( .C (clk), .D (new_AGEMA_signal_15846), .Q (new_AGEMA_signal_15847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8026 ( .C (clk), .D (new_AGEMA_signal_15850), .Q (new_AGEMA_signal_15851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8030 ( .C (clk), .D (new_AGEMA_signal_15854), .Q (new_AGEMA_signal_15855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8034 ( .C (clk), .D (new_AGEMA_signal_15858), .Q (new_AGEMA_signal_15859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8038 ( .C (clk), .D (new_AGEMA_signal_15862), .Q (new_AGEMA_signal_15863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8042 ( .C (clk), .D (new_AGEMA_signal_15866), .Q (new_AGEMA_signal_15867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8046 ( .C (clk), .D (new_AGEMA_signal_15870), .Q (new_AGEMA_signal_15871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8050 ( .C (clk), .D (new_AGEMA_signal_15874), .Q (new_AGEMA_signal_15875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8054 ( .C (clk), .D (new_AGEMA_signal_15878), .Q (new_AGEMA_signal_15879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8058 ( .C (clk), .D (new_AGEMA_signal_15882), .Q (new_AGEMA_signal_15883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8062 ( .C (clk), .D (new_AGEMA_signal_15886), .Q (new_AGEMA_signal_15887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8066 ( .C (clk), .D (new_AGEMA_signal_15890), .Q (new_AGEMA_signal_15891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8070 ( .C (clk), .D (new_AGEMA_signal_15894), .Q (new_AGEMA_signal_15895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8074 ( .C (clk), .D (new_AGEMA_signal_15898), .Q (new_AGEMA_signal_15899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8078 ( .C (clk), .D (new_AGEMA_signal_15902), .Q (new_AGEMA_signal_15903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8082 ( .C (clk), .D (new_AGEMA_signal_15906), .Q (new_AGEMA_signal_15907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8086 ( .C (clk), .D (new_AGEMA_signal_15910), .Q (new_AGEMA_signal_15911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8090 ( .C (clk), .D (new_AGEMA_signal_15914), .Q (new_AGEMA_signal_15915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8094 ( .C (clk), .D (new_AGEMA_signal_15918), .Q (new_AGEMA_signal_15919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8098 ( .C (clk), .D (new_AGEMA_signal_15922), .Q (new_AGEMA_signal_15923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8102 ( .C (clk), .D (new_AGEMA_signal_15926), .Q (new_AGEMA_signal_15927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8106 ( .C (clk), .D (new_AGEMA_signal_15930), .Q (new_AGEMA_signal_15931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8110 ( .C (clk), .D (new_AGEMA_signal_15934), .Q (new_AGEMA_signal_15935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8114 ( .C (clk), .D (new_AGEMA_signal_15938), .Q (new_AGEMA_signal_15939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8118 ( .C (clk), .D (new_AGEMA_signal_15942), .Q (new_AGEMA_signal_15943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8122 ( .C (clk), .D (new_AGEMA_signal_15946), .Q (new_AGEMA_signal_15947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8126 ( .C (clk), .D (new_AGEMA_signal_15950), .Q (new_AGEMA_signal_15951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8130 ( .C (clk), .D (new_AGEMA_signal_15954), .Q (new_AGEMA_signal_15955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8134 ( .C (clk), .D (new_AGEMA_signal_15958), .Q (new_AGEMA_signal_15959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8138 ( .C (clk), .D (new_AGEMA_signal_15962), .Q (new_AGEMA_signal_15963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8142 ( .C (clk), .D (new_AGEMA_signal_15966), .Q (new_AGEMA_signal_15967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8146 ( .C (clk), .D (new_AGEMA_signal_15970), .Q (new_AGEMA_signal_15971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8150 ( .C (clk), .D (new_AGEMA_signal_15974), .Q (new_AGEMA_signal_15975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8154 ( .C (clk), .D (new_AGEMA_signal_15978), .Q (new_AGEMA_signal_15979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8158 ( .C (clk), .D (new_AGEMA_signal_15982), .Q (new_AGEMA_signal_15983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8162 ( .C (clk), .D (new_AGEMA_signal_15986), .Q (new_AGEMA_signal_15987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8166 ( .C (clk), .D (new_AGEMA_signal_15990), .Q (new_AGEMA_signal_15991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8170 ( .C (clk), .D (new_AGEMA_signal_15994), .Q (new_AGEMA_signal_15995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8174 ( .C (clk), .D (new_AGEMA_signal_15998), .Q (new_AGEMA_signal_15999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8178 ( .C (clk), .D (new_AGEMA_signal_16002), .Q (new_AGEMA_signal_16003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8182 ( .C (clk), .D (new_AGEMA_signal_16006), .Q (new_AGEMA_signal_16007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8186 ( .C (clk), .D (new_AGEMA_signal_16010), .Q (new_AGEMA_signal_16011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8190 ( .C (clk), .D (new_AGEMA_signal_16014), .Q (new_AGEMA_signal_16015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8194 ( .C (clk), .D (new_AGEMA_signal_16018), .Q (new_AGEMA_signal_16019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8198 ( .C (clk), .D (new_AGEMA_signal_16022), .Q (new_AGEMA_signal_16023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8202 ( .C (clk), .D (new_AGEMA_signal_16026), .Q (new_AGEMA_signal_16027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8206 ( .C (clk), .D (new_AGEMA_signal_16030), .Q (new_AGEMA_signal_16031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8210 ( .C (clk), .D (new_AGEMA_signal_16034), .Q (new_AGEMA_signal_16035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8214 ( .C (clk), .D (new_AGEMA_signal_16038), .Q (new_AGEMA_signal_16039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8218 ( .C (clk), .D (new_AGEMA_signal_16042), .Q (new_AGEMA_signal_16043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8222 ( .C (clk), .D (new_AGEMA_signal_16046), .Q (new_AGEMA_signal_16047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8226 ( .C (clk), .D (new_AGEMA_signal_16050), .Q (new_AGEMA_signal_16051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8230 ( .C (clk), .D (new_AGEMA_signal_16054), .Q (new_AGEMA_signal_16055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8234 ( .C (clk), .D (new_AGEMA_signal_16058), .Q (new_AGEMA_signal_16059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8238 ( .C (clk), .D (new_AGEMA_signal_16062), .Q (new_AGEMA_signal_16063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8242 ( .C (clk), .D (new_AGEMA_signal_16066), .Q (new_AGEMA_signal_16067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8246 ( .C (clk), .D (new_AGEMA_signal_16070), .Q (new_AGEMA_signal_16071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8250 ( .C (clk), .D (new_AGEMA_signal_16074), .Q (new_AGEMA_signal_16075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8254 ( .C (clk), .D (new_AGEMA_signal_16078), .Q (new_AGEMA_signal_16079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8258 ( .C (clk), .D (new_AGEMA_signal_16082), .Q (new_AGEMA_signal_16083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8262 ( .C (clk), .D (new_AGEMA_signal_16086), .Q (new_AGEMA_signal_16087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8266 ( .C (clk), .D (new_AGEMA_signal_16090), .Q (new_AGEMA_signal_16091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8270 ( .C (clk), .D (new_AGEMA_signal_16094), .Q (new_AGEMA_signal_16095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8274 ( .C (clk), .D (new_AGEMA_signal_16098), .Q (new_AGEMA_signal_16099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8278 ( .C (clk), .D (new_AGEMA_signal_16102), .Q (new_AGEMA_signal_16103) ) ;
    buf_clk new_AGEMA_reg_buffer_8282 ( .C (clk), .D (new_AGEMA_signal_16106), .Q (new_AGEMA_signal_16107) ) ;
    buf_clk new_AGEMA_reg_buffer_8286 ( .C (clk), .D (new_AGEMA_signal_16110), .Q (new_AGEMA_signal_16111) ) ;
    buf_clk new_AGEMA_reg_buffer_8290 ( .C (clk), .D (new_AGEMA_signal_16114), .Q (new_AGEMA_signal_16115) ) ;
    buf_clk new_AGEMA_reg_buffer_8294 ( .C (clk), .D (new_AGEMA_signal_16118), .Q (new_AGEMA_signal_16119) ) ;
    buf_clk new_AGEMA_reg_buffer_8298 ( .C (clk), .D (new_AGEMA_signal_16122), .Q (new_AGEMA_signal_16123) ) ;
    buf_clk new_AGEMA_reg_buffer_8302 ( .C (clk), .D (new_AGEMA_signal_16126), .Q (new_AGEMA_signal_16127) ) ;
    buf_clk new_AGEMA_reg_buffer_8306 ( .C (clk), .D (new_AGEMA_signal_16130), .Q (new_AGEMA_signal_16131) ) ;
    buf_clk new_AGEMA_reg_buffer_8310 ( .C (clk), .D (new_AGEMA_signal_16134), .Q (new_AGEMA_signal_16135) ) ;
    buf_clk new_AGEMA_reg_buffer_8314 ( .C (clk), .D (new_AGEMA_signal_16138), .Q (new_AGEMA_signal_16139) ) ;
    buf_clk new_AGEMA_reg_buffer_8318 ( .C (clk), .D (new_AGEMA_signal_16142), .Q (new_AGEMA_signal_16143) ) ;
    buf_clk new_AGEMA_reg_buffer_8322 ( .C (clk), .D (new_AGEMA_signal_16146), .Q (new_AGEMA_signal_16147) ) ;
    buf_clk new_AGEMA_reg_buffer_8326 ( .C (clk), .D (new_AGEMA_signal_16150), .Q (new_AGEMA_signal_16151) ) ;
    buf_clk new_AGEMA_reg_buffer_8330 ( .C (clk), .D (new_AGEMA_signal_16154), .Q (new_AGEMA_signal_16155) ) ;
    buf_clk new_AGEMA_reg_buffer_8334 ( .C (clk), .D (new_AGEMA_signal_16158), .Q (new_AGEMA_signal_16159) ) ;
    buf_clk new_AGEMA_reg_buffer_8338 ( .C (clk), .D (new_AGEMA_signal_16162), .Q (new_AGEMA_signal_16163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8342 ( .C (clk), .D (new_AGEMA_signal_16166), .Q (new_AGEMA_signal_16167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8346 ( .C (clk), .D (new_AGEMA_signal_16170), .Q (new_AGEMA_signal_16171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8350 ( .C (clk), .D (new_AGEMA_signal_16174), .Q (new_AGEMA_signal_16175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8354 ( .C (clk), .D (new_AGEMA_signal_16178), .Q (new_AGEMA_signal_16179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8358 ( .C (clk), .D (new_AGEMA_signal_16182), .Q (new_AGEMA_signal_16183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8362 ( .C (clk), .D (new_AGEMA_signal_16186), .Q (new_AGEMA_signal_16187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8366 ( .C (clk), .D (new_AGEMA_signal_16190), .Q (new_AGEMA_signal_16191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8370 ( .C (clk), .D (new_AGEMA_signal_16194), .Q (new_AGEMA_signal_16195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8374 ( .C (clk), .D (new_AGEMA_signal_16198), .Q (new_AGEMA_signal_16199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8378 ( .C (clk), .D (new_AGEMA_signal_16202), .Q (new_AGEMA_signal_16203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8382 ( .C (clk), .D (new_AGEMA_signal_16206), .Q (new_AGEMA_signal_16207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8386 ( .C (clk), .D (new_AGEMA_signal_16210), .Q (new_AGEMA_signal_16211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8390 ( .C (clk), .D (new_AGEMA_signal_16214), .Q (new_AGEMA_signal_16215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8394 ( .C (clk), .D (new_AGEMA_signal_16218), .Q (new_AGEMA_signal_16219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8398 ( .C (clk), .D (new_AGEMA_signal_16222), .Q (new_AGEMA_signal_16223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8402 ( .C (clk), .D (new_AGEMA_signal_16226), .Q (new_AGEMA_signal_16227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8406 ( .C (clk), .D (new_AGEMA_signal_16230), .Q (new_AGEMA_signal_16231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8410 ( .C (clk), .D (new_AGEMA_signal_16234), .Q (new_AGEMA_signal_16235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8414 ( .C (clk), .D (new_AGEMA_signal_16238), .Q (new_AGEMA_signal_16239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8418 ( .C (clk), .D (new_AGEMA_signal_16242), .Q (new_AGEMA_signal_16243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8422 ( .C (clk), .D (new_AGEMA_signal_16246), .Q (new_AGEMA_signal_16247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8426 ( .C (clk), .D (new_AGEMA_signal_16250), .Q (new_AGEMA_signal_16251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8430 ( .C (clk), .D (new_AGEMA_signal_16254), .Q (new_AGEMA_signal_16255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8434 ( .C (clk), .D (new_AGEMA_signal_16258), .Q (new_AGEMA_signal_16259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8438 ( .C (clk), .D (new_AGEMA_signal_16262), .Q (new_AGEMA_signal_16263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8442 ( .C (clk), .D (new_AGEMA_signal_16266), .Q (new_AGEMA_signal_16267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8446 ( .C (clk), .D (new_AGEMA_signal_16270), .Q (new_AGEMA_signal_16271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8450 ( .C (clk), .D (new_AGEMA_signal_16274), .Q (new_AGEMA_signal_16275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8454 ( .C (clk), .D (new_AGEMA_signal_16278), .Q (new_AGEMA_signal_16279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8458 ( .C (clk), .D (new_AGEMA_signal_16282), .Q (new_AGEMA_signal_16283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8462 ( .C (clk), .D (new_AGEMA_signal_16286), .Q (new_AGEMA_signal_16287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8466 ( .C (clk), .D (new_AGEMA_signal_16290), .Q (new_AGEMA_signal_16291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8470 ( .C (clk), .D (new_AGEMA_signal_16294), .Q (new_AGEMA_signal_16295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8474 ( .C (clk), .D (new_AGEMA_signal_16298), .Q (new_AGEMA_signal_16299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8478 ( .C (clk), .D (new_AGEMA_signal_16302), .Q (new_AGEMA_signal_16303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8482 ( .C (clk), .D (new_AGEMA_signal_16306), .Q (new_AGEMA_signal_16307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8486 ( .C (clk), .D (new_AGEMA_signal_16310), .Q (new_AGEMA_signal_16311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8490 ( .C (clk), .D (new_AGEMA_signal_16314), .Q (new_AGEMA_signal_16315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8494 ( .C (clk), .D (new_AGEMA_signal_16318), .Q (new_AGEMA_signal_16319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8498 ( .C (clk), .D (new_AGEMA_signal_16322), .Q (new_AGEMA_signal_16323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8502 ( .C (clk), .D (new_AGEMA_signal_16326), .Q (new_AGEMA_signal_16327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8506 ( .C (clk), .D (new_AGEMA_signal_16330), .Q (new_AGEMA_signal_16331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8510 ( .C (clk), .D (new_AGEMA_signal_16334), .Q (new_AGEMA_signal_16335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8514 ( .C (clk), .D (new_AGEMA_signal_16338), .Q (new_AGEMA_signal_16339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8518 ( .C (clk), .D (new_AGEMA_signal_16342), .Q (new_AGEMA_signal_16343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8522 ( .C (clk), .D (new_AGEMA_signal_16346), .Q (new_AGEMA_signal_16347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8526 ( .C (clk), .D (new_AGEMA_signal_16350), .Q (new_AGEMA_signal_16351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8530 ( .C (clk), .D (new_AGEMA_signal_16354), .Q (new_AGEMA_signal_16355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8534 ( .C (clk), .D (new_AGEMA_signal_16358), .Q (new_AGEMA_signal_16359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8538 ( .C (clk), .D (new_AGEMA_signal_16362), .Q (new_AGEMA_signal_16363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8542 ( .C (clk), .D (new_AGEMA_signal_16366), .Q (new_AGEMA_signal_16367) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8546 ( .C (clk), .D (new_AGEMA_signal_16370), .Q (new_AGEMA_signal_16371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8550 ( .C (clk), .D (new_AGEMA_signal_16374), .Q (new_AGEMA_signal_16375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8554 ( .C (clk), .D (new_AGEMA_signal_16378), .Q (new_AGEMA_signal_16379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8558 ( .C (clk), .D (new_AGEMA_signal_16382), .Q (new_AGEMA_signal_16383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8562 ( .C (clk), .D (new_AGEMA_signal_16386), .Q (new_AGEMA_signal_16387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8566 ( .C (clk), .D (new_AGEMA_signal_16390), .Q (new_AGEMA_signal_16391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8570 ( .C (clk), .D (new_AGEMA_signal_16394), .Q (new_AGEMA_signal_16395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8574 ( .C (clk), .D (new_AGEMA_signal_16398), .Q (new_AGEMA_signal_16399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8578 ( .C (clk), .D (new_AGEMA_signal_16402), .Q (new_AGEMA_signal_16403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8582 ( .C (clk), .D (new_AGEMA_signal_16406), .Q (new_AGEMA_signal_16407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8586 ( .C (clk), .D (new_AGEMA_signal_16410), .Q (new_AGEMA_signal_16411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8590 ( .C (clk), .D (new_AGEMA_signal_16414), .Q (new_AGEMA_signal_16415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8594 ( .C (clk), .D (new_AGEMA_signal_16418), .Q (new_AGEMA_signal_16419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8598 ( .C (clk), .D (new_AGEMA_signal_16422), .Q (new_AGEMA_signal_16423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8602 ( .C (clk), .D (new_AGEMA_signal_16426), .Q (new_AGEMA_signal_16427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8606 ( .C (clk), .D (new_AGEMA_signal_16430), .Q (new_AGEMA_signal_16431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8610 ( .C (clk), .D (new_AGEMA_signal_16434), .Q (new_AGEMA_signal_16435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8614 ( .C (clk), .D (new_AGEMA_signal_16438), .Q (new_AGEMA_signal_16439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8618 ( .C (clk), .D (new_AGEMA_signal_16442), .Q (new_AGEMA_signal_16443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8622 ( .C (clk), .D (new_AGEMA_signal_16446), .Q (new_AGEMA_signal_16447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8626 ( .C (clk), .D (new_AGEMA_signal_16450), .Q (new_AGEMA_signal_16451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8630 ( .C (clk), .D (new_AGEMA_signal_16454), .Q (new_AGEMA_signal_16455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8634 ( .C (clk), .D (new_AGEMA_signal_16458), .Q (new_AGEMA_signal_16459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8638 ( .C (clk), .D (new_AGEMA_signal_16462), .Q (new_AGEMA_signal_16463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8642 ( .C (clk), .D (new_AGEMA_signal_16466), .Q (new_AGEMA_signal_16467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8646 ( .C (clk), .D (new_AGEMA_signal_16470), .Q (new_AGEMA_signal_16471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8650 ( .C (clk), .D (new_AGEMA_signal_16474), .Q (new_AGEMA_signal_16475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8654 ( .C (clk), .D (new_AGEMA_signal_16478), .Q (new_AGEMA_signal_16479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8658 ( .C (clk), .D (new_AGEMA_signal_16482), .Q (new_AGEMA_signal_16483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8662 ( .C (clk), .D (new_AGEMA_signal_16486), .Q (new_AGEMA_signal_16487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8666 ( .C (clk), .D (new_AGEMA_signal_16490), .Q (new_AGEMA_signal_16491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8670 ( .C (clk), .D (new_AGEMA_signal_16494), .Q (new_AGEMA_signal_16495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8674 ( .C (clk), .D (new_AGEMA_signal_16498), .Q (new_AGEMA_signal_16499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8678 ( .C (clk), .D (new_AGEMA_signal_16502), .Q (new_AGEMA_signal_16503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8682 ( .C (clk), .D (new_AGEMA_signal_16506), .Q (new_AGEMA_signal_16507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8686 ( .C (clk), .D (new_AGEMA_signal_16510), .Q (new_AGEMA_signal_16511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8690 ( .C (clk), .D (new_AGEMA_signal_16514), .Q (new_AGEMA_signal_16515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8694 ( .C (clk), .D (new_AGEMA_signal_16518), .Q (new_AGEMA_signal_16519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8698 ( .C (clk), .D (new_AGEMA_signal_16522), .Q (new_AGEMA_signal_16523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8702 ( .C (clk), .D (new_AGEMA_signal_16526), .Q (new_AGEMA_signal_16527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8706 ( .C (clk), .D (new_AGEMA_signal_16530), .Q (new_AGEMA_signal_16531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8710 ( .C (clk), .D (new_AGEMA_signal_16534), .Q (new_AGEMA_signal_16535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8714 ( .C (clk), .D (new_AGEMA_signal_16538), .Q (new_AGEMA_signal_16539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8718 ( .C (clk), .D (new_AGEMA_signal_16542), .Q (new_AGEMA_signal_16543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8722 ( .C (clk), .D (new_AGEMA_signal_16546), .Q (new_AGEMA_signal_16547) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8726 ( .C (clk), .D (new_AGEMA_signal_16550), .Q (new_AGEMA_signal_16551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8730 ( .C (clk), .D (new_AGEMA_signal_16554), .Q (new_AGEMA_signal_16555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8734 ( .C (clk), .D (new_AGEMA_signal_16558), .Q (new_AGEMA_signal_16559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8738 ( .C (clk), .D (new_AGEMA_signal_16562), .Q (new_AGEMA_signal_16563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8742 ( .C (clk), .D (new_AGEMA_signal_16566), .Q (new_AGEMA_signal_16567) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8746 ( .C (clk), .D (new_AGEMA_signal_16570), .Q (new_AGEMA_signal_16571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8750 ( .C (clk), .D (new_AGEMA_signal_16574), .Q (new_AGEMA_signal_16575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8754 ( .C (clk), .D (new_AGEMA_signal_16578), .Q (new_AGEMA_signal_16579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8758 ( .C (clk), .D (new_AGEMA_signal_16582), .Q (new_AGEMA_signal_16583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8762 ( .C (clk), .D (new_AGEMA_signal_16586), .Q (new_AGEMA_signal_16587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8766 ( .C (clk), .D (new_AGEMA_signal_16590), .Q (new_AGEMA_signal_16591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8770 ( .C (clk), .D (new_AGEMA_signal_16594), .Q (new_AGEMA_signal_16595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8774 ( .C (clk), .D (new_AGEMA_signal_16598), .Q (new_AGEMA_signal_16599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8778 ( .C (clk), .D (new_AGEMA_signal_16602), .Q (new_AGEMA_signal_16603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8782 ( .C (clk), .D (new_AGEMA_signal_16606), .Q (new_AGEMA_signal_16607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8786 ( .C (clk), .D (new_AGEMA_signal_16610), .Q (new_AGEMA_signal_16611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8790 ( .C (clk), .D (new_AGEMA_signal_16614), .Q (new_AGEMA_signal_16615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8794 ( .C (clk), .D (new_AGEMA_signal_16618), .Q (new_AGEMA_signal_16619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8798 ( .C (clk), .D (new_AGEMA_signal_16622), .Q (new_AGEMA_signal_16623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8802 ( .C (clk), .D (new_AGEMA_signal_16626), .Q (new_AGEMA_signal_16627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8806 ( .C (clk), .D (new_AGEMA_signal_16630), .Q (new_AGEMA_signal_16631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8810 ( .C (clk), .D (new_AGEMA_signal_16634), .Q (new_AGEMA_signal_16635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8814 ( .C (clk), .D (new_AGEMA_signal_16638), .Q (new_AGEMA_signal_16639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8818 ( .C (clk), .D (new_AGEMA_signal_16642), .Q (new_AGEMA_signal_16643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8822 ( .C (clk), .D (new_AGEMA_signal_16646), .Q (new_AGEMA_signal_16647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8826 ( .C (clk), .D (new_AGEMA_signal_16650), .Q (new_AGEMA_signal_16651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8830 ( .C (clk), .D (new_AGEMA_signal_16654), .Q (new_AGEMA_signal_16655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8834 ( .C (clk), .D (new_AGEMA_signal_16658), .Q (new_AGEMA_signal_16659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8838 ( .C (clk), .D (new_AGEMA_signal_16662), .Q (new_AGEMA_signal_16663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8842 ( .C (clk), .D (new_AGEMA_signal_16666), .Q (new_AGEMA_signal_16667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8846 ( .C (clk), .D (new_AGEMA_signal_16670), .Q (new_AGEMA_signal_16671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8850 ( .C (clk), .D (new_AGEMA_signal_16674), .Q (new_AGEMA_signal_16675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8854 ( .C (clk), .D (new_AGEMA_signal_16678), .Q (new_AGEMA_signal_16679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8858 ( .C (clk), .D (new_AGEMA_signal_16682), .Q (new_AGEMA_signal_16683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8862 ( .C (clk), .D (new_AGEMA_signal_16686), .Q (new_AGEMA_signal_16687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8866 ( .C (clk), .D (new_AGEMA_signal_16690), .Q (new_AGEMA_signal_16691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8870 ( .C (clk), .D (new_AGEMA_signal_16694), .Q (new_AGEMA_signal_16695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8874 ( .C (clk), .D (new_AGEMA_signal_16698), .Q (new_AGEMA_signal_16699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8878 ( .C (clk), .D (new_AGEMA_signal_16702), .Q (new_AGEMA_signal_16703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8882 ( .C (clk), .D (new_AGEMA_signal_16706), .Q (new_AGEMA_signal_16707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8886 ( .C (clk), .D (new_AGEMA_signal_16710), .Q (new_AGEMA_signal_16711) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8890 ( .C (clk), .D (new_AGEMA_signal_16714), .Q (new_AGEMA_signal_16715) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8894 ( .C (clk), .D (new_AGEMA_signal_16718), .Q (new_AGEMA_signal_16719) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8898 ( .C (clk), .D (new_AGEMA_signal_16722), .Q (new_AGEMA_signal_16723) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8902 ( .C (clk), .D (new_AGEMA_signal_16726), .Q (new_AGEMA_signal_16727) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8906 ( .C (clk), .D (new_AGEMA_signal_16730), .Q (new_AGEMA_signal_16731) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8910 ( .C (clk), .D (new_AGEMA_signal_16734), .Q (new_AGEMA_signal_16735) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8914 ( .C (clk), .D (new_AGEMA_signal_16738), .Q (new_AGEMA_signal_16739) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8918 ( .C (clk), .D (new_AGEMA_signal_16742), .Q (new_AGEMA_signal_16743) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8922 ( .C (clk), .D (new_AGEMA_signal_16746), .Q (new_AGEMA_signal_16747) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8926 ( .C (clk), .D (new_AGEMA_signal_16750), .Q (new_AGEMA_signal_16751) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8930 ( .C (clk), .D (new_AGEMA_signal_16754), .Q (new_AGEMA_signal_16755) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8934 ( .C (clk), .D (new_AGEMA_signal_16758), .Q (new_AGEMA_signal_16759) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8938 ( .C (clk), .D (new_AGEMA_signal_16762), .Q (new_AGEMA_signal_16763) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8942 ( .C (clk), .D (new_AGEMA_signal_16766), .Q (new_AGEMA_signal_16767) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8946 ( .C (clk), .D (new_AGEMA_signal_16770), .Q (new_AGEMA_signal_16771) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8950 ( .C (clk), .D (new_AGEMA_signal_16774), .Q (new_AGEMA_signal_16775) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8954 ( .C (clk), .D (new_AGEMA_signal_16778), .Q (new_AGEMA_signal_16779) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8958 ( .C (clk), .D (new_AGEMA_signal_16782), .Q (new_AGEMA_signal_16783) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8962 ( .C (clk), .D (new_AGEMA_signal_16786), .Q (new_AGEMA_signal_16787) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8966 ( .C (clk), .D (new_AGEMA_signal_16790), .Q (new_AGEMA_signal_16791) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8970 ( .C (clk), .D (new_AGEMA_signal_16794), .Q (new_AGEMA_signal_16795) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8974 ( .C (clk), .D (new_AGEMA_signal_16798), .Q (new_AGEMA_signal_16799) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8978 ( .C (clk), .D (new_AGEMA_signal_16802), .Q (new_AGEMA_signal_16803) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8982 ( .C (clk), .D (new_AGEMA_signal_16806), .Q (new_AGEMA_signal_16807) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8986 ( .C (clk), .D (new_AGEMA_signal_16810), .Q (new_AGEMA_signal_16811) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8990 ( .C (clk), .D (new_AGEMA_signal_16814), .Q (new_AGEMA_signal_16815) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8994 ( .C (clk), .D (new_AGEMA_signal_16818), .Q (new_AGEMA_signal_16819) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8998 ( .C (clk), .D (new_AGEMA_signal_16822), .Q (new_AGEMA_signal_16823) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9002 ( .C (clk), .D (new_AGEMA_signal_16826), .Q (new_AGEMA_signal_16827) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9006 ( .C (clk), .D (new_AGEMA_signal_16830), .Q (new_AGEMA_signal_16831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9010 ( .C (clk), .D (new_AGEMA_signal_16834), .Q (new_AGEMA_signal_16835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9014 ( .C (clk), .D (new_AGEMA_signal_16838), .Q (new_AGEMA_signal_16839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9018 ( .C (clk), .D (new_AGEMA_signal_16842), .Q (new_AGEMA_signal_16843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9022 ( .C (clk), .D (new_AGEMA_signal_16846), .Q (new_AGEMA_signal_16847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9026 ( .C (clk), .D (new_AGEMA_signal_16850), .Q (new_AGEMA_signal_16851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9030 ( .C (clk), .D (new_AGEMA_signal_16854), .Q (new_AGEMA_signal_16855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9034 ( .C (clk), .D (new_AGEMA_signal_16858), .Q (new_AGEMA_signal_16859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9038 ( .C (clk), .D (new_AGEMA_signal_16862), .Q (new_AGEMA_signal_16863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9042 ( .C (clk), .D (new_AGEMA_signal_16866), .Q (new_AGEMA_signal_16867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9046 ( .C (clk), .D (new_AGEMA_signal_16870), .Q (new_AGEMA_signal_16871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9050 ( .C (clk), .D (new_AGEMA_signal_16874), .Q (new_AGEMA_signal_16875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9054 ( .C (clk), .D (new_AGEMA_signal_16878), .Q (new_AGEMA_signal_16879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9058 ( .C (clk), .D (new_AGEMA_signal_16882), .Q (new_AGEMA_signal_16883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9062 ( .C (clk), .D (new_AGEMA_signal_16886), .Q (new_AGEMA_signal_16887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9066 ( .C (clk), .D (new_AGEMA_signal_16890), .Q (new_AGEMA_signal_16891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9070 ( .C (clk), .D (new_AGEMA_signal_16894), .Q (new_AGEMA_signal_16895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9074 ( .C (clk), .D (new_AGEMA_signal_16898), .Q (new_AGEMA_signal_16899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9078 ( .C (clk), .D (new_AGEMA_signal_16902), .Q (new_AGEMA_signal_16903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9082 ( .C (clk), .D (new_AGEMA_signal_16906), .Q (new_AGEMA_signal_16907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9086 ( .C (clk), .D (new_AGEMA_signal_16910), .Q (new_AGEMA_signal_16911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9090 ( .C (clk), .D (new_AGEMA_signal_16914), .Q (new_AGEMA_signal_16915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9094 ( .C (clk), .D (new_AGEMA_signal_16918), .Q (new_AGEMA_signal_16919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9098 ( .C (clk), .D (new_AGEMA_signal_16922), .Q (new_AGEMA_signal_16923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9102 ( .C (clk), .D (new_AGEMA_signal_16926), .Q (new_AGEMA_signal_16927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9106 ( .C (clk), .D (new_AGEMA_signal_16930), .Q (new_AGEMA_signal_16931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9110 ( .C (clk), .D (new_AGEMA_signal_16934), .Q (new_AGEMA_signal_16935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9114 ( .C (clk), .D (new_AGEMA_signal_16938), .Q (new_AGEMA_signal_16939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9118 ( .C (clk), .D (new_AGEMA_signal_16942), .Q (new_AGEMA_signal_16943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9122 ( .C (clk), .D (new_AGEMA_signal_16946), .Q (new_AGEMA_signal_16947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9126 ( .C (clk), .D (new_AGEMA_signal_16950), .Q (new_AGEMA_signal_16951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9130 ( .C (clk), .D (new_AGEMA_signal_16954), .Q (new_AGEMA_signal_16955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9134 ( .C (clk), .D (new_AGEMA_signal_16958), .Q (new_AGEMA_signal_16959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9138 ( .C (clk), .D (new_AGEMA_signal_16962), .Q (new_AGEMA_signal_16963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9142 ( .C (clk), .D (new_AGEMA_signal_16966), .Q (new_AGEMA_signal_16967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9146 ( .C (clk), .D (new_AGEMA_signal_16970), .Q (new_AGEMA_signal_16971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9150 ( .C (clk), .D (new_AGEMA_signal_16974), .Q (new_AGEMA_signal_16975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9154 ( .C (clk), .D (new_AGEMA_signal_16978), .Q (new_AGEMA_signal_16979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9158 ( .C (clk), .D (new_AGEMA_signal_16982), .Q (new_AGEMA_signal_16983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9162 ( .C (clk), .D (new_AGEMA_signal_16986), .Q (new_AGEMA_signal_16987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9166 ( .C (clk), .D (new_AGEMA_signal_16990), .Q (new_AGEMA_signal_16991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9170 ( .C (clk), .D (new_AGEMA_signal_16994), .Q (new_AGEMA_signal_16995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9174 ( .C (clk), .D (new_AGEMA_signal_16998), .Q (new_AGEMA_signal_16999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9178 ( .C (clk), .D (new_AGEMA_signal_17002), .Q (new_AGEMA_signal_17003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9182 ( .C (clk), .D (new_AGEMA_signal_17006), .Q (new_AGEMA_signal_17007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9186 ( .C (clk), .D (new_AGEMA_signal_17010), .Q (new_AGEMA_signal_17011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9190 ( .C (clk), .D (new_AGEMA_signal_17014), .Q (new_AGEMA_signal_17015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9194 ( .C (clk), .D (new_AGEMA_signal_17018), .Q (new_AGEMA_signal_17019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9198 ( .C (clk), .D (new_AGEMA_signal_17022), .Q (new_AGEMA_signal_17023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9202 ( .C (clk), .D (new_AGEMA_signal_17026), .Q (new_AGEMA_signal_17027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9206 ( .C (clk), .D (new_AGEMA_signal_17030), .Q (new_AGEMA_signal_17031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9210 ( .C (clk), .D (new_AGEMA_signal_17034), .Q (new_AGEMA_signal_17035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9214 ( .C (clk), .D (new_AGEMA_signal_17038), .Q (new_AGEMA_signal_17039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9218 ( .C (clk), .D (new_AGEMA_signal_17042), .Q (new_AGEMA_signal_17043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9222 ( .C (clk), .D (new_AGEMA_signal_17046), .Q (new_AGEMA_signal_17047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9226 ( .C (clk), .D (new_AGEMA_signal_17050), .Q (new_AGEMA_signal_17051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9230 ( .C (clk), .D (new_AGEMA_signal_17054), .Q (new_AGEMA_signal_17055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9234 ( .C (clk), .D (new_AGEMA_signal_17058), .Q (new_AGEMA_signal_17059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9238 ( .C (clk), .D (new_AGEMA_signal_17062), .Q (new_AGEMA_signal_17063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9242 ( .C (clk), .D (new_AGEMA_signal_17066), .Q (new_AGEMA_signal_17067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9246 ( .C (clk), .D (new_AGEMA_signal_17070), .Q (new_AGEMA_signal_17071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9250 ( .C (clk), .D (new_AGEMA_signal_17074), .Q (new_AGEMA_signal_17075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9254 ( .C (clk), .D (new_AGEMA_signal_17078), .Q (new_AGEMA_signal_17079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9258 ( .C (clk), .D (new_AGEMA_signal_17082), .Q (new_AGEMA_signal_17083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9262 ( .C (clk), .D (new_AGEMA_signal_17086), .Q (new_AGEMA_signal_17087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9266 ( .C (clk), .D (new_AGEMA_signal_17090), .Q (new_AGEMA_signal_17091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9270 ( .C (clk), .D (new_AGEMA_signal_17094), .Q (new_AGEMA_signal_17095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9274 ( .C (clk), .D (new_AGEMA_signal_17098), .Q (new_AGEMA_signal_17099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9278 ( .C (clk), .D (new_AGEMA_signal_17102), .Q (new_AGEMA_signal_17103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9282 ( .C (clk), .D (new_AGEMA_signal_17106), .Q (new_AGEMA_signal_17107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9286 ( .C (clk), .D (new_AGEMA_signal_17110), .Q (new_AGEMA_signal_17111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9290 ( .C (clk), .D (new_AGEMA_signal_17114), .Q (new_AGEMA_signal_17115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9294 ( .C (clk), .D (new_AGEMA_signal_17118), .Q (new_AGEMA_signal_17119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9298 ( .C (clk), .D (new_AGEMA_signal_17122), .Q (new_AGEMA_signal_17123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9302 ( .C (clk), .D (new_AGEMA_signal_17126), .Q (new_AGEMA_signal_17127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9306 ( .C (clk), .D (new_AGEMA_signal_17130), .Q (new_AGEMA_signal_17131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9310 ( .C (clk), .D (new_AGEMA_signal_17134), .Q (new_AGEMA_signal_17135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9314 ( .C (clk), .D (new_AGEMA_signal_17138), .Q (new_AGEMA_signal_17139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9318 ( .C (clk), .D (new_AGEMA_signal_17142), .Q (new_AGEMA_signal_17143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9322 ( .C (clk), .D (new_AGEMA_signal_17146), .Q (new_AGEMA_signal_17147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9326 ( .C (clk), .D (new_AGEMA_signal_17150), .Q (new_AGEMA_signal_17151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9330 ( .C (clk), .D (new_AGEMA_signal_17154), .Q (new_AGEMA_signal_17155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9334 ( .C (clk), .D (new_AGEMA_signal_17158), .Q (new_AGEMA_signal_17159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9338 ( .C (clk), .D (new_AGEMA_signal_17162), .Q (new_AGEMA_signal_17163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9342 ( .C (clk), .D (new_AGEMA_signal_17166), .Q (new_AGEMA_signal_17167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9346 ( .C (clk), .D (new_AGEMA_signal_17170), .Q (new_AGEMA_signal_17171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9350 ( .C (clk), .D (new_AGEMA_signal_17174), .Q (new_AGEMA_signal_17175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9354 ( .C (clk), .D (new_AGEMA_signal_17178), .Q (new_AGEMA_signal_17179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9358 ( .C (clk), .D (new_AGEMA_signal_17182), .Q (new_AGEMA_signal_17183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9362 ( .C (clk), .D (new_AGEMA_signal_17186), .Q (new_AGEMA_signal_17187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9366 ( .C (clk), .D (new_AGEMA_signal_17190), .Q (new_AGEMA_signal_17191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9370 ( .C (clk), .D (new_AGEMA_signal_17194), .Q (new_AGEMA_signal_17195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9374 ( .C (clk), .D (new_AGEMA_signal_17198), .Q (new_AGEMA_signal_17199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9378 ( .C (clk), .D (new_AGEMA_signal_17202), .Q (new_AGEMA_signal_17203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9382 ( .C (clk), .D (new_AGEMA_signal_17206), .Q (new_AGEMA_signal_17207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9386 ( .C (clk), .D (new_AGEMA_signal_17210), .Q (new_AGEMA_signal_17211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9390 ( .C (clk), .D (new_AGEMA_signal_17214), .Q (new_AGEMA_signal_17215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9394 ( .C (clk), .D (new_AGEMA_signal_17218), .Q (new_AGEMA_signal_17219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9398 ( .C (clk), .D (new_AGEMA_signal_17222), .Q (new_AGEMA_signal_17223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9402 ( .C (clk), .D (new_AGEMA_signal_17226), .Q (new_AGEMA_signal_17227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9406 ( .C (clk), .D (new_AGEMA_signal_17230), .Q (new_AGEMA_signal_17231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9410 ( .C (clk), .D (new_AGEMA_signal_17234), .Q (new_AGEMA_signal_17235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9414 ( .C (clk), .D (new_AGEMA_signal_17238), .Q (new_AGEMA_signal_17239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9418 ( .C (clk), .D (new_AGEMA_signal_17242), .Q (new_AGEMA_signal_17243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9422 ( .C (clk), .D (new_AGEMA_signal_17246), .Q (new_AGEMA_signal_17247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9426 ( .C (clk), .D (new_AGEMA_signal_17250), .Q (new_AGEMA_signal_17251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9430 ( .C (clk), .D (new_AGEMA_signal_17254), .Q (new_AGEMA_signal_17255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9434 ( .C (clk), .D (new_AGEMA_signal_17258), .Q (new_AGEMA_signal_17259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9438 ( .C (clk), .D (new_AGEMA_signal_17262), .Q (new_AGEMA_signal_17263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9442 ( .C (clk), .D (new_AGEMA_signal_17266), .Q (new_AGEMA_signal_17267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9446 ( .C (clk), .D (new_AGEMA_signal_17270), .Q (new_AGEMA_signal_17271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9450 ( .C (clk), .D (new_AGEMA_signal_17274), .Q (new_AGEMA_signal_17275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9454 ( .C (clk), .D (new_AGEMA_signal_17278), .Q (new_AGEMA_signal_17279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9458 ( .C (clk), .D (new_AGEMA_signal_17282), .Q (new_AGEMA_signal_17283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9462 ( .C (clk), .D (new_AGEMA_signal_17286), .Q (new_AGEMA_signal_17287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9466 ( .C (clk), .D (new_AGEMA_signal_17290), .Q (new_AGEMA_signal_17291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9470 ( .C (clk), .D (new_AGEMA_signal_17294), .Q (new_AGEMA_signal_17295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9474 ( .C (clk), .D (new_AGEMA_signal_17298), .Q (new_AGEMA_signal_17299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9478 ( .C (clk), .D (new_AGEMA_signal_17302), .Q (new_AGEMA_signal_17303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9482 ( .C (clk), .D (new_AGEMA_signal_17306), .Q (new_AGEMA_signal_17307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9486 ( .C (clk), .D (new_AGEMA_signal_17310), .Q (new_AGEMA_signal_17311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9490 ( .C (clk), .D (new_AGEMA_signal_17314), .Q (new_AGEMA_signal_17315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9494 ( .C (clk), .D (new_AGEMA_signal_17318), .Q (new_AGEMA_signal_17319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9498 ( .C (clk), .D (new_AGEMA_signal_17322), .Q (new_AGEMA_signal_17323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9502 ( .C (clk), .D (new_AGEMA_signal_17326), .Q (new_AGEMA_signal_17327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9506 ( .C (clk), .D (new_AGEMA_signal_17330), .Q (new_AGEMA_signal_17331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9510 ( .C (clk), .D (new_AGEMA_signal_17334), .Q (new_AGEMA_signal_17335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9514 ( .C (clk), .D (new_AGEMA_signal_17338), .Q (new_AGEMA_signal_17339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9518 ( .C (clk), .D (new_AGEMA_signal_17342), .Q (new_AGEMA_signal_17343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9522 ( .C (clk), .D (new_AGEMA_signal_17346), .Q (new_AGEMA_signal_17347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9526 ( .C (clk), .D (new_AGEMA_signal_17350), .Q (new_AGEMA_signal_17351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9530 ( .C (clk), .D (new_AGEMA_signal_17354), .Q (new_AGEMA_signal_17355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9534 ( .C (clk), .D (new_AGEMA_signal_17358), .Q (new_AGEMA_signal_17359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9538 ( .C (clk), .D (new_AGEMA_signal_17362), .Q (new_AGEMA_signal_17363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9542 ( .C (clk), .D (new_AGEMA_signal_17366), .Q (new_AGEMA_signal_17367) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9546 ( .C (clk), .D (new_AGEMA_signal_17370), .Q (new_AGEMA_signal_17371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9550 ( .C (clk), .D (new_AGEMA_signal_17374), .Q (new_AGEMA_signal_17375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9554 ( .C (clk), .D (new_AGEMA_signal_17378), .Q (new_AGEMA_signal_17379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9558 ( .C (clk), .D (new_AGEMA_signal_17382), .Q (new_AGEMA_signal_17383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9562 ( .C (clk), .D (new_AGEMA_signal_17386), .Q (new_AGEMA_signal_17387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9566 ( .C (clk), .D (new_AGEMA_signal_17390), .Q (new_AGEMA_signal_17391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9570 ( .C (clk), .D (new_AGEMA_signal_17394), .Q (new_AGEMA_signal_17395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9574 ( .C (clk), .D (new_AGEMA_signal_17398), .Q (new_AGEMA_signal_17399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9578 ( .C (clk), .D (new_AGEMA_signal_17402), .Q (new_AGEMA_signal_17403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9582 ( .C (clk), .D (new_AGEMA_signal_17406), .Q (new_AGEMA_signal_17407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9586 ( .C (clk), .D (new_AGEMA_signal_17410), .Q (new_AGEMA_signal_17411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9590 ( .C (clk), .D (new_AGEMA_signal_17414), .Q (new_AGEMA_signal_17415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9594 ( .C (clk), .D (new_AGEMA_signal_17418), .Q (new_AGEMA_signal_17419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9598 ( .C (clk), .D (new_AGEMA_signal_17422), .Q (new_AGEMA_signal_17423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9602 ( .C (clk), .D (new_AGEMA_signal_17426), .Q (new_AGEMA_signal_17427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9606 ( .C (clk), .D (new_AGEMA_signal_17430), .Q (new_AGEMA_signal_17431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9610 ( .C (clk), .D (new_AGEMA_signal_17434), .Q (new_AGEMA_signal_17435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9614 ( .C (clk), .D (new_AGEMA_signal_17438), .Q (new_AGEMA_signal_17439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9618 ( .C (clk), .D (new_AGEMA_signal_17442), .Q (new_AGEMA_signal_17443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9622 ( .C (clk), .D (new_AGEMA_signal_17446), .Q (new_AGEMA_signal_17447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9626 ( .C (clk), .D (new_AGEMA_signal_17450), .Q (new_AGEMA_signal_17451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9630 ( .C (clk), .D (new_AGEMA_signal_17454), .Q (new_AGEMA_signal_17455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9634 ( .C (clk), .D (new_AGEMA_signal_17458), .Q (new_AGEMA_signal_17459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9638 ( .C (clk), .D (new_AGEMA_signal_17462), .Q (new_AGEMA_signal_17463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9642 ( .C (clk), .D (new_AGEMA_signal_17466), .Q (new_AGEMA_signal_17467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9646 ( .C (clk), .D (new_AGEMA_signal_17470), .Q (new_AGEMA_signal_17471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9650 ( .C (clk), .D (new_AGEMA_signal_17474), .Q (new_AGEMA_signal_17475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9654 ( .C (clk), .D (new_AGEMA_signal_17478), .Q (new_AGEMA_signal_17479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9658 ( .C (clk), .D (new_AGEMA_signal_17482), .Q (new_AGEMA_signal_17483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9662 ( .C (clk), .D (new_AGEMA_signal_17486), .Q (new_AGEMA_signal_17487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9666 ( .C (clk), .D (new_AGEMA_signal_17490), .Q (new_AGEMA_signal_17491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9670 ( .C (clk), .D (new_AGEMA_signal_17494), .Q (new_AGEMA_signal_17495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9674 ( .C (clk), .D (new_AGEMA_signal_17498), .Q (new_AGEMA_signal_17499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9678 ( .C (clk), .D (new_AGEMA_signal_17502), .Q (new_AGEMA_signal_17503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9682 ( .C (clk), .D (new_AGEMA_signal_17506), .Q (new_AGEMA_signal_17507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9686 ( .C (clk), .D (new_AGEMA_signal_17510), .Q (new_AGEMA_signal_17511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9690 ( .C (clk), .D (new_AGEMA_signal_17514), .Q (new_AGEMA_signal_17515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9694 ( .C (clk), .D (new_AGEMA_signal_17518), .Q (new_AGEMA_signal_17519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9698 ( .C (clk), .D (new_AGEMA_signal_17522), .Q (new_AGEMA_signal_17523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9702 ( .C (clk), .D (new_AGEMA_signal_17526), .Q (new_AGEMA_signal_17527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9706 ( .C (clk), .D (new_AGEMA_signal_17530), .Q (new_AGEMA_signal_17531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9710 ( .C (clk), .D (new_AGEMA_signal_17534), .Q (new_AGEMA_signal_17535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9714 ( .C (clk), .D (new_AGEMA_signal_17538), .Q (new_AGEMA_signal_17539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9718 ( .C (clk), .D (new_AGEMA_signal_17542), .Q (new_AGEMA_signal_17543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9722 ( .C (clk), .D (new_AGEMA_signal_17546), .Q (new_AGEMA_signal_17547) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9726 ( .C (clk), .D (new_AGEMA_signal_17550), .Q (new_AGEMA_signal_17551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9730 ( .C (clk), .D (new_AGEMA_signal_17554), .Q (new_AGEMA_signal_17555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9734 ( .C (clk), .D (new_AGEMA_signal_17558), .Q (new_AGEMA_signal_17559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9738 ( .C (clk), .D (new_AGEMA_signal_17562), .Q (new_AGEMA_signal_17563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9742 ( .C (clk), .D (new_AGEMA_signal_17566), .Q (new_AGEMA_signal_17567) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9746 ( .C (clk), .D (new_AGEMA_signal_17570), .Q (new_AGEMA_signal_17571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9750 ( .C (clk), .D (new_AGEMA_signal_17574), .Q (new_AGEMA_signal_17575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9754 ( .C (clk), .D (new_AGEMA_signal_17578), .Q (new_AGEMA_signal_17579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9758 ( .C (clk), .D (new_AGEMA_signal_17582), .Q (new_AGEMA_signal_17583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9762 ( .C (clk), .D (new_AGEMA_signal_17586), .Q (new_AGEMA_signal_17587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9766 ( .C (clk), .D (new_AGEMA_signal_17590), .Q (new_AGEMA_signal_17591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9770 ( .C (clk), .D (new_AGEMA_signal_17594), .Q (new_AGEMA_signal_17595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9774 ( .C (clk), .D (new_AGEMA_signal_17598), .Q (new_AGEMA_signal_17599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9778 ( .C (clk), .D (new_AGEMA_signal_17602), .Q (new_AGEMA_signal_17603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9782 ( .C (clk), .D (new_AGEMA_signal_17606), .Q (new_AGEMA_signal_17607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9786 ( .C (clk), .D (new_AGEMA_signal_17610), .Q (new_AGEMA_signal_17611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9790 ( .C (clk), .D (new_AGEMA_signal_17614), .Q (new_AGEMA_signal_17615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9794 ( .C (clk), .D (new_AGEMA_signal_17618), .Q (new_AGEMA_signal_17619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9798 ( .C (clk), .D (new_AGEMA_signal_17622), .Q (new_AGEMA_signal_17623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9802 ( .C (clk), .D (new_AGEMA_signal_17626), .Q (new_AGEMA_signal_17627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9806 ( .C (clk), .D (new_AGEMA_signal_17630), .Q (new_AGEMA_signal_17631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9810 ( .C (clk), .D (new_AGEMA_signal_17634), .Q (new_AGEMA_signal_17635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9814 ( .C (clk), .D (new_AGEMA_signal_17638), .Q (new_AGEMA_signal_17639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9818 ( .C (clk), .D (new_AGEMA_signal_17642), .Q (new_AGEMA_signal_17643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9822 ( .C (clk), .D (new_AGEMA_signal_17646), .Q (new_AGEMA_signal_17647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9826 ( .C (clk), .D (new_AGEMA_signal_17650), .Q (new_AGEMA_signal_17651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9830 ( .C (clk), .D (new_AGEMA_signal_17654), .Q (new_AGEMA_signal_17655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9834 ( .C (clk), .D (new_AGEMA_signal_17658), .Q (new_AGEMA_signal_17659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9838 ( .C (clk), .D (new_AGEMA_signal_17662), .Q (new_AGEMA_signal_17663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9842 ( .C (clk), .D (new_AGEMA_signal_17666), .Q (new_AGEMA_signal_17667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9846 ( .C (clk), .D (new_AGEMA_signal_17670), .Q (new_AGEMA_signal_17671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9850 ( .C (clk), .D (new_AGEMA_signal_17674), .Q (new_AGEMA_signal_17675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9854 ( .C (clk), .D (new_AGEMA_signal_17678), .Q (new_AGEMA_signal_17679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9858 ( .C (clk), .D (new_AGEMA_signal_17682), .Q (new_AGEMA_signal_17683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9862 ( .C (clk), .D (new_AGEMA_signal_17686), .Q (new_AGEMA_signal_17687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9866 ( .C (clk), .D (new_AGEMA_signal_17690), .Q (new_AGEMA_signal_17691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9870 ( .C (clk), .D (new_AGEMA_signal_17694), .Q (new_AGEMA_signal_17695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9874 ( .C (clk), .D (new_AGEMA_signal_17698), .Q (new_AGEMA_signal_17699) ) ;
    buf_clk new_AGEMA_reg_buffer_9878 ( .C (clk), .D (new_AGEMA_signal_17702), .Q (new_AGEMA_signal_17703) ) ;
    buf_clk new_AGEMA_reg_buffer_9882 ( .C (clk), .D (new_AGEMA_signal_17706), .Q (new_AGEMA_signal_17707) ) ;
    buf_clk new_AGEMA_reg_buffer_9886 ( .C (clk), .D (new_AGEMA_signal_17710), .Q (new_AGEMA_signal_17711) ) ;
    buf_clk new_AGEMA_reg_buffer_9890 ( .C (clk), .D (new_AGEMA_signal_17714), .Q (new_AGEMA_signal_17715) ) ;
    buf_clk new_AGEMA_reg_buffer_9894 ( .C (clk), .D (new_AGEMA_signal_17718), .Q (new_AGEMA_signal_17719) ) ;
    buf_clk new_AGEMA_reg_buffer_9898 ( .C (clk), .D (new_AGEMA_signal_17722), .Q (new_AGEMA_signal_17723) ) ;
    buf_clk new_AGEMA_reg_buffer_9902 ( .C (clk), .D (new_AGEMA_signal_17726), .Q (new_AGEMA_signal_17727) ) ;

    /* cells in depth 3 */
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_5094, new_AGEMA_signal_5093, new_AGEMA_signal_5092, SubBytesIns_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_9961, new_AGEMA_signal_9960, new_AGEMA_signal_9959, new_AGEMA_signal_9958}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_5148, new_AGEMA_signal_5147, new_AGEMA_signal_5146, SubBytesIns_Inst_Sbox_0_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_5091, new_AGEMA_signal_5090, new_AGEMA_signal_5089, SubBytesIns_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_9965, new_AGEMA_signal_9964, new_AGEMA_signal_9963, new_AGEMA_signal_9962}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_5151, new_AGEMA_signal_5150, new_AGEMA_signal_5149, SubBytesIns_Inst_Sbox_0_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_9961, new_AGEMA_signal_9960, new_AGEMA_signal_9959, new_AGEMA_signal_9958}), .b ({new_AGEMA_signal_5097, new_AGEMA_signal_5096, new_AGEMA_signal_5095, SubBytesIns_Inst_Sbox_0_M31}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_5154, new_AGEMA_signal_5153, new_AGEMA_signal_5152, SubBytesIns_Inst_Sbox_0_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_9965, new_AGEMA_signal_9964, new_AGEMA_signal_9963, new_AGEMA_signal_9962}), .b ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, new_AGEMA_signal_5047, SubBytesIns_Inst_Sbox_0_M34}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_5157, new_AGEMA_signal_5156, new_AGEMA_signal_5155, SubBytesIns_Inst_Sbox_0_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_10017, new_AGEMA_signal_10016, new_AGEMA_signal_10015, new_AGEMA_signal_10014}), .b ({new_AGEMA_signal_5148, new_AGEMA_signal_5147, new_AGEMA_signal_5146, SubBytesIns_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_5208, new_AGEMA_signal_5207, new_AGEMA_signal_5206, SubBytesIns_Inst_Sbox_0_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_5154, new_AGEMA_signal_5153, new_AGEMA_signal_5152, SubBytesIns_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_10021, new_AGEMA_signal_10020, new_AGEMA_signal_10019, new_AGEMA_signal_10018}), .c ({new_AGEMA_signal_5211, new_AGEMA_signal_5210, new_AGEMA_signal_5209, SubBytesIns_Inst_Sbox_0_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_10025, new_AGEMA_signal_10024, new_AGEMA_signal_10023, new_AGEMA_signal_10022}), .b ({new_AGEMA_signal_5151, new_AGEMA_signal_5150, new_AGEMA_signal_5149, SubBytesIns_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_5214, new_AGEMA_signal_5213, new_AGEMA_signal_5212, SubBytesIns_Inst_Sbox_0_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_5157, new_AGEMA_signal_5156, new_AGEMA_signal_5155, SubBytesIns_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_10029, new_AGEMA_signal_10028, new_AGEMA_signal_10027, new_AGEMA_signal_10026}), .c ({new_AGEMA_signal_5217, new_AGEMA_signal_5216, new_AGEMA_signal_5215, SubBytesIns_Inst_Sbox_0_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_5211, new_AGEMA_signal_5210, new_AGEMA_signal_5209, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_5217, new_AGEMA_signal_5216, new_AGEMA_signal_5215, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_5256, new_AGEMA_signal_5255, new_AGEMA_signal_5254, SubBytesIns_Inst_Sbox_0_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_5208, new_AGEMA_signal_5207, new_AGEMA_signal_5206, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_5214, new_AGEMA_signal_5213, new_AGEMA_signal_5212, SubBytesIns_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_5259, new_AGEMA_signal_5258, new_AGEMA_signal_5257, SubBytesIns_Inst_Sbox_0_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_5208, new_AGEMA_signal_5207, new_AGEMA_signal_5206, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_5211, new_AGEMA_signal_5210, new_AGEMA_signal_5209, SubBytesIns_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_5262, new_AGEMA_signal_5261, new_AGEMA_signal_5260, SubBytesIns_Inst_Sbox_0_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_5214, new_AGEMA_signal_5213, new_AGEMA_signal_5212, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_5217, new_AGEMA_signal_5216, new_AGEMA_signal_5215, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_5265, new_AGEMA_signal_5264, new_AGEMA_signal_5263, SubBytesIns_Inst_Sbox_0_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_5259, new_AGEMA_signal_5258, new_AGEMA_signal_5257, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_5256, new_AGEMA_signal_5255, new_AGEMA_signal_5254, SubBytesIns_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, new_AGEMA_signal_5398, SubBytesIns_Inst_Sbox_0_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_5109, new_AGEMA_signal_5108, new_AGEMA_signal_5107, SubBytesIns_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_9977, new_AGEMA_signal_9976, new_AGEMA_signal_9975, new_AGEMA_signal_9974}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630], Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_5163, new_AGEMA_signal_5162, new_AGEMA_signal_5161, SubBytesIns_Inst_Sbox_1_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_5106, new_AGEMA_signal_5105, new_AGEMA_signal_5104, SubBytesIns_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_9981, new_AGEMA_signal_9980, new_AGEMA_signal_9979, new_AGEMA_signal_9978}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_5166, new_AGEMA_signal_5165, new_AGEMA_signal_5164, SubBytesIns_Inst_Sbox_1_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_9977, new_AGEMA_signal_9976, new_AGEMA_signal_9975, new_AGEMA_signal_9974}), .b ({new_AGEMA_signal_5112, new_AGEMA_signal_5111, new_AGEMA_signal_5110, SubBytesIns_Inst_Sbox_1_M31}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_5169, new_AGEMA_signal_5168, new_AGEMA_signal_5167, SubBytesIns_Inst_Sbox_1_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_9981, new_AGEMA_signal_9980, new_AGEMA_signal_9979, new_AGEMA_signal_9978}), .b ({new_AGEMA_signal_5061, new_AGEMA_signal_5060, new_AGEMA_signal_5059, SubBytesIns_Inst_Sbox_1_M34}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_5172, new_AGEMA_signal_5171, new_AGEMA_signal_5170, SubBytesIns_Inst_Sbox_1_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_10033, new_AGEMA_signal_10032, new_AGEMA_signal_10031, new_AGEMA_signal_10030}), .b ({new_AGEMA_signal_5163, new_AGEMA_signal_5162, new_AGEMA_signal_5161, SubBytesIns_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_5220, new_AGEMA_signal_5219, new_AGEMA_signal_5218, SubBytesIns_Inst_Sbox_1_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_5169, new_AGEMA_signal_5168, new_AGEMA_signal_5167, SubBytesIns_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_10037, new_AGEMA_signal_10036, new_AGEMA_signal_10035, new_AGEMA_signal_10034}), .c ({new_AGEMA_signal_5223, new_AGEMA_signal_5222, new_AGEMA_signal_5221, SubBytesIns_Inst_Sbox_1_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_10041, new_AGEMA_signal_10040, new_AGEMA_signal_10039, new_AGEMA_signal_10038}), .b ({new_AGEMA_signal_5166, new_AGEMA_signal_5165, new_AGEMA_signal_5164, SubBytesIns_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_5226, new_AGEMA_signal_5225, new_AGEMA_signal_5224, SubBytesIns_Inst_Sbox_1_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_5172, new_AGEMA_signal_5171, new_AGEMA_signal_5170, SubBytesIns_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_10045, new_AGEMA_signal_10044, new_AGEMA_signal_10043, new_AGEMA_signal_10042}), .c ({new_AGEMA_signal_5229, new_AGEMA_signal_5228, new_AGEMA_signal_5227, SubBytesIns_Inst_Sbox_1_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_5223, new_AGEMA_signal_5222, new_AGEMA_signal_5221, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_5229, new_AGEMA_signal_5228, new_AGEMA_signal_5227, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_5292, new_AGEMA_signal_5291, new_AGEMA_signal_5290, SubBytesIns_Inst_Sbox_1_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_5220, new_AGEMA_signal_5219, new_AGEMA_signal_5218, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_5226, new_AGEMA_signal_5225, new_AGEMA_signal_5224, SubBytesIns_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_5295, new_AGEMA_signal_5294, new_AGEMA_signal_5293, SubBytesIns_Inst_Sbox_1_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_5220, new_AGEMA_signal_5219, new_AGEMA_signal_5218, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_5223, new_AGEMA_signal_5222, new_AGEMA_signal_5221, SubBytesIns_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_5298, new_AGEMA_signal_5297, new_AGEMA_signal_5296, SubBytesIns_Inst_Sbox_1_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_5226, new_AGEMA_signal_5225, new_AGEMA_signal_5224, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_5229, new_AGEMA_signal_5228, new_AGEMA_signal_5227, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, new_AGEMA_signal_5299, SubBytesIns_Inst_Sbox_1_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_5295, new_AGEMA_signal_5294, new_AGEMA_signal_5293, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_5292, new_AGEMA_signal_5291, new_AGEMA_signal_5290, SubBytesIns_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_5436, new_AGEMA_signal_5435, new_AGEMA_signal_5434, SubBytesIns_Inst_Sbox_1_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_5124, new_AGEMA_signal_5123, new_AGEMA_signal_5122, SubBytesIns_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_9993, new_AGEMA_signal_9992, new_AGEMA_signal_9991, new_AGEMA_signal_9990}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_5178, new_AGEMA_signal_5177, new_AGEMA_signal_5176, SubBytesIns_Inst_Sbox_2_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_5121, new_AGEMA_signal_5120, new_AGEMA_signal_5119, SubBytesIns_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_9997, new_AGEMA_signal_9996, new_AGEMA_signal_9995, new_AGEMA_signal_9994}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690], Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_5181, new_AGEMA_signal_5180, new_AGEMA_signal_5179, SubBytesIns_Inst_Sbox_2_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_9993, new_AGEMA_signal_9992, new_AGEMA_signal_9991, new_AGEMA_signal_9990}), .b ({new_AGEMA_signal_5127, new_AGEMA_signal_5126, new_AGEMA_signal_5125, SubBytesIns_Inst_Sbox_2_M31}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702], Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_5184, new_AGEMA_signal_5183, new_AGEMA_signal_5182, SubBytesIns_Inst_Sbox_2_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_9997, new_AGEMA_signal_9996, new_AGEMA_signal_9995, new_AGEMA_signal_9994}), .b ({new_AGEMA_signal_5073, new_AGEMA_signal_5072, new_AGEMA_signal_5071, SubBytesIns_Inst_Sbox_2_M34}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_5187, new_AGEMA_signal_5186, new_AGEMA_signal_5185, SubBytesIns_Inst_Sbox_2_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_10049, new_AGEMA_signal_10048, new_AGEMA_signal_10047, new_AGEMA_signal_10046}), .b ({new_AGEMA_signal_5178, new_AGEMA_signal_5177, new_AGEMA_signal_5176, SubBytesIns_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_5232, new_AGEMA_signal_5231, new_AGEMA_signal_5230, SubBytesIns_Inst_Sbox_2_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_5184, new_AGEMA_signal_5183, new_AGEMA_signal_5182, SubBytesIns_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_10053, new_AGEMA_signal_10052, new_AGEMA_signal_10051, new_AGEMA_signal_10050}), .c ({new_AGEMA_signal_5235, new_AGEMA_signal_5234, new_AGEMA_signal_5233, SubBytesIns_Inst_Sbox_2_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_10057, new_AGEMA_signal_10056, new_AGEMA_signal_10055, new_AGEMA_signal_10054}), .b ({new_AGEMA_signal_5181, new_AGEMA_signal_5180, new_AGEMA_signal_5179, SubBytesIns_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_5238, new_AGEMA_signal_5237, new_AGEMA_signal_5236, SubBytesIns_Inst_Sbox_2_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_5187, new_AGEMA_signal_5186, new_AGEMA_signal_5185, SubBytesIns_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_10061, new_AGEMA_signal_10060, new_AGEMA_signal_10059, new_AGEMA_signal_10058}), .c ({new_AGEMA_signal_5241, new_AGEMA_signal_5240, new_AGEMA_signal_5239, SubBytesIns_Inst_Sbox_2_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_5235, new_AGEMA_signal_5234, new_AGEMA_signal_5233, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_5241, new_AGEMA_signal_5240, new_AGEMA_signal_5239, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, new_AGEMA_signal_5326, SubBytesIns_Inst_Sbox_2_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_5232, new_AGEMA_signal_5231, new_AGEMA_signal_5230, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_5238, new_AGEMA_signal_5237, new_AGEMA_signal_5236, SubBytesIns_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_5331, new_AGEMA_signal_5330, new_AGEMA_signal_5329, SubBytesIns_Inst_Sbox_2_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_5232, new_AGEMA_signal_5231, new_AGEMA_signal_5230, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_5235, new_AGEMA_signal_5234, new_AGEMA_signal_5233, SubBytesIns_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_5334, new_AGEMA_signal_5333, new_AGEMA_signal_5332, SubBytesIns_Inst_Sbox_2_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_5238, new_AGEMA_signal_5237, new_AGEMA_signal_5236, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_5241, new_AGEMA_signal_5240, new_AGEMA_signal_5239, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_5337, new_AGEMA_signal_5336, new_AGEMA_signal_5335, SubBytesIns_Inst_Sbox_2_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_5331, new_AGEMA_signal_5330, new_AGEMA_signal_5329, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, new_AGEMA_signal_5326, SubBytesIns_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_5472, new_AGEMA_signal_5471, new_AGEMA_signal_5470, SubBytesIns_Inst_Sbox_2_M45}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_5139, new_AGEMA_signal_5138, new_AGEMA_signal_5137, SubBytesIns_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_10009, new_AGEMA_signal_10008, new_AGEMA_signal_10007, new_AGEMA_signal_10006}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_5193, new_AGEMA_signal_5192, new_AGEMA_signal_5191, SubBytesIns_Inst_Sbox_3_M29}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_5136, new_AGEMA_signal_5135, new_AGEMA_signal_5134, SubBytesIns_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_10013, new_AGEMA_signal_10012, new_AGEMA_signal_10011, new_AGEMA_signal_10010}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738], Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_5196, new_AGEMA_signal_5195, new_AGEMA_signal_5194, SubBytesIns_Inst_Sbox_3_M30}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_10009, new_AGEMA_signal_10008, new_AGEMA_signal_10007, new_AGEMA_signal_10006}), .b ({new_AGEMA_signal_5142, new_AGEMA_signal_5141, new_AGEMA_signal_5140, SubBytesIns_Inst_Sbox_3_M31}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750], Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_5199, new_AGEMA_signal_5198, new_AGEMA_signal_5197, SubBytesIns_Inst_Sbox_3_M32}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_10013, new_AGEMA_signal_10012, new_AGEMA_signal_10011, new_AGEMA_signal_10010}), .b ({new_AGEMA_signal_5085, new_AGEMA_signal_5084, new_AGEMA_signal_5083, SubBytesIns_Inst_Sbox_3_M34}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_5202, new_AGEMA_signal_5201, new_AGEMA_signal_5200, SubBytesIns_Inst_Sbox_3_M35}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_10065, new_AGEMA_signal_10064, new_AGEMA_signal_10063, new_AGEMA_signal_10062}), .b ({new_AGEMA_signal_5193, new_AGEMA_signal_5192, new_AGEMA_signal_5191, SubBytesIns_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_5244, new_AGEMA_signal_5243, new_AGEMA_signal_5242, SubBytesIns_Inst_Sbox_3_M37}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_5199, new_AGEMA_signal_5198, new_AGEMA_signal_5197, SubBytesIns_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_10069, new_AGEMA_signal_10068, new_AGEMA_signal_10067, new_AGEMA_signal_10066}), .c ({new_AGEMA_signal_5247, new_AGEMA_signal_5246, new_AGEMA_signal_5245, SubBytesIns_Inst_Sbox_3_M38}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_10073, new_AGEMA_signal_10072, new_AGEMA_signal_10071, new_AGEMA_signal_10070}), .b ({new_AGEMA_signal_5196, new_AGEMA_signal_5195, new_AGEMA_signal_5194, SubBytesIns_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_5250, new_AGEMA_signal_5249, new_AGEMA_signal_5248, SubBytesIns_Inst_Sbox_3_M39}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_5202, new_AGEMA_signal_5201, new_AGEMA_signal_5200, SubBytesIns_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_10077, new_AGEMA_signal_10076, new_AGEMA_signal_10075, new_AGEMA_signal_10074}), .c ({new_AGEMA_signal_5253, new_AGEMA_signal_5252, new_AGEMA_signal_5251, SubBytesIns_Inst_Sbox_3_M40}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_5247, new_AGEMA_signal_5246, new_AGEMA_signal_5245, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_5253, new_AGEMA_signal_5252, new_AGEMA_signal_5251, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, new_AGEMA_signal_5362, SubBytesIns_Inst_Sbox_3_M41}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_5244, new_AGEMA_signal_5243, new_AGEMA_signal_5242, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_5250, new_AGEMA_signal_5249, new_AGEMA_signal_5248, SubBytesIns_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_5367, new_AGEMA_signal_5366, new_AGEMA_signal_5365, SubBytesIns_Inst_Sbox_3_M42}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_5244, new_AGEMA_signal_5243, new_AGEMA_signal_5242, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_5247, new_AGEMA_signal_5246, new_AGEMA_signal_5245, SubBytesIns_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_5370, new_AGEMA_signal_5369, new_AGEMA_signal_5368, SubBytesIns_Inst_Sbox_3_M43}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_5250, new_AGEMA_signal_5249, new_AGEMA_signal_5248, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_5253, new_AGEMA_signal_5252, new_AGEMA_signal_5251, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_5373, new_AGEMA_signal_5372, new_AGEMA_signal_5371, SubBytesIns_Inst_Sbox_3_M44}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_5367, new_AGEMA_signal_5366, new_AGEMA_signal_5365, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, new_AGEMA_signal_5362, SubBytesIns_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, new_AGEMA_signal_5506, SubBytesIns_Inst_Sbox_3_M45}) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2189 ( .C (clk), .D (new_AGEMA_signal_9950), .Q (new_AGEMA_signal_10014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2190 ( .C (clk), .D (new_AGEMA_signal_9951), .Q (new_AGEMA_signal_10015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2191 ( .C (clk), .D (new_AGEMA_signal_9952), .Q (new_AGEMA_signal_10016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2192 ( .C (clk), .D (new_AGEMA_signal_9953), .Q (new_AGEMA_signal_10017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2193 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M33), .Q (new_AGEMA_signal_10018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2194 ( .C (clk), .D (new_AGEMA_signal_5098), .Q (new_AGEMA_signal_10019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2195 ( .C (clk), .D (new_AGEMA_signal_5099), .Q (new_AGEMA_signal_10020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2196 ( .C (clk), .D (new_AGEMA_signal_5100), .Q (new_AGEMA_signal_10021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2197 ( .C (clk), .D (new_AGEMA_signal_9954), .Q (new_AGEMA_signal_10022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2198 ( .C (clk), .D (new_AGEMA_signal_9955), .Q (new_AGEMA_signal_10023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2199 ( .C (clk), .D (new_AGEMA_signal_9956), .Q (new_AGEMA_signal_10024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2200 ( .C (clk), .D (new_AGEMA_signal_9957), .Q (new_AGEMA_signal_10025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2201 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M36), .Q (new_AGEMA_signal_10026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2202 ( .C (clk), .D (new_AGEMA_signal_5158), .Q (new_AGEMA_signal_10027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2203 ( .C (clk), .D (new_AGEMA_signal_5159), .Q (new_AGEMA_signal_10028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2204 ( .C (clk), .D (new_AGEMA_signal_5160), .Q (new_AGEMA_signal_10029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2205 ( .C (clk), .D (new_AGEMA_signal_9966), .Q (new_AGEMA_signal_10030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2206 ( .C (clk), .D (new_AGEMA_signal_9967), .Q (new_AGEMA_signal_10031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2207 ( .C (clk), .D (new_AGEMA_signal_9968), .Q (new_AGEMA_signal_10032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2208 ( .C (clk), .D (new_AGEMA_signal_9969), .Q (new_AGEMA_signal_10033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2209 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M33), .Q (new_AGEMA_signal_10034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2210 ( .C (clk), .D (new_AGEMA_signal_5113), .Q (new_AGEMA_signal_10035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2211 ( .C (clk), .D (new_AGEMA_signal_5114), .Q (new_AGEMA_signal_10036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2212 ( .C (clk), .D (new_AGEMA_signal_5115), .Q (new_AGEMA_signal_10037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2213 ( .C (clk), .D (new_AGEMA_signal_9970), .Q (new_AGEMA_signal_10038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2214 ( .C (clk), .D (new_AGEMA_signal_9971), .Q (new_AGEMA_signal_10039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2215 ( .C (clk), .D (new_AGEMA_signal_9972), .Q (new_AGEMA_signal_10040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2216 ( .C (clk), .D (new_AGEMA_signal_9973), .Q (new_AGEMA_signal_10041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2217 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M36), .Q (new_AGEMA_signal_10042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2218 ( .C (clk), .D (new_AGEMA_signal_5173), .Q (new_AGEMA_signal_10043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2219 ( .C (clk), .D (new_AGEMA_signal_5174), .Q (new_AGEMA_signal_10044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2220 ( .C (clk), .D (new_AGEMA_signal_5175), .Q (new_AGEMA_signal_10045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2221 ( .C (clk), .D (new_AGEMA_signal_9982), .Q (new_AGEMA_signal_10046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2222 ( .C (clk), .D (new_AGEMA_signal_9983), .Q (new_AGEMA_signal_10047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2223 ( .C (clk), .D (new_AGEMA_signal_9984), .Q (new_AGEMA_signal_10048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2224 ( .C (clk), .D (new_AGEMA_signal_9985), .Q (new_AGEMA_signal_10049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2225 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M33), .Q (new_AGEMA_signal_10050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2226 ( .C (clk), .D (new_AGEMA_signal_5128), .Q (new_AGEMA_signal_10051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2227 ( .C (clk), .D (new_AGEMA_signal_5129), .Q (new_AGEMA_signal_10052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2228 ( .C (clk), .D (new_AGEMA_signal_5130), .Q (new_AGEMA_signal_10053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2229 ( .C (clk), .D (new_AGEMA_signal_9986), .Q (new_AGEMA_signal_10054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2230 ( .C (clk), .D (new_AGEMA_signal_9987), .Q (new_AGEMA_signal_10055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2231 ( .C (clk), .D (new_AGEMA_signal_9988), .Q (new_AGEMA_signal_10056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2232 ( .C (clk), .D (new_AGEMA_signal_9989), .Q (new_AGEMA_signal_10057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2233 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M36), .Q (new_AGEMA_signal_10058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2234 ( .C (clk), .D (new_AGEMA_signal_5188), .Q (new_AGEMA_signal_10059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2235 ( .C (clk), .D (new_AGEMA_signal_5189), .Q (new_AGEMA_signal_10060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2236 ( .C (clk), .D (new_AGEMA_signal_5190), .Q (new_AGEMA_signal_10061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2237 ( .C (clk), .D (new_AGEMA_signal_9998), .Q (new_AGEMA_signal_10062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2238 ( .C (clk), .D (new_AGEMA_signal_9999), .Q (new_AGEMA_signal_10063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2239 ( .C (clk), .D (new_AGEMA_signal_10000), .Q (new_AGEMA_signal_10064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2240 ( .C (clk), .D (new_AGEMA_signal_10001), .Q (new_AGEMA_signal_10065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2241 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M33), .Q (new_AGEMA_signal_10066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2242 ( .C (clk), .D (new_AGEMA_signal_5143), .Q (new_AGEMA_signal_10067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2243 ( .C (clk), .D (new_AGEMA_signal_5144), .Q (new_AGEMA_signal_10068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2244 ( .C (clk), .D (new_AGEMA_signal_5145), .Q (new_AGEMA_signal_10069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2245 ( .C (clk), .D (new_AGEMA_signal_10002), .Q (new_AGEMA_signal_10070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2246 ( .C (clk), .D (new_AGEMA_signal_10003), .Q (new_AGEMA_signal_10071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2247 ( .C (clk), .D (new_AGEMA_signal_10004), .Q (new_AGEMA_signal_10072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2248 ( .C (clk), .D (new_AGEMA_signal_10005), .Q (new_AGEMA_signal_10073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2249 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M36), .Q (new_AGEMA_signal_10074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2250 ( .C (clk), .D (new_AGEMA_signal_5203), .Q (new_AGEMA_signal_10075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2251 ( .C (clk), .D (new_AGEMA_signal_5204), .Q (new_AGEMA_signal_10076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2252 ( .C (clk), .D (new_AGEMA_signal_5205), .Q (new_AGEMA_signal_10077) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C (clk), .D (new_AGEMA_signal_10079), .Q (new_AGEMA_signal_10080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2259 ( .C (clk), .D (new_AGEMA_signal_10083), .Q (new_AGEMA_signal_10084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2263 ( .C (clk), .D (new_AGEMA_signal_10087), .Q (new_AGEMA_signal_10088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2267 ( .C (clk), .D (new_AGEMA_signal_10091), .Q (new_AGEMA_signal_10092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2271 ( .C (clk), .D (new_AGEMA_signal_10095), .Q (new_AGEMA_signal_10096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2275 ( .C (clk), .D (new_AGEMA_signal_10099), .Q (new_AGEMA_signal_10100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2279 ( .C (clk), .D (new_AGEMA_signal_10103), .Q (new_AGEMA_signal_10104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2283 ( .C (clk), .D (new_AGEMA_signal_10107), .Q (new_AGEMA_signal_10108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2287 ( .C (clk), .D (new_AGEMA_signal_10111), .Q (new_AGEMA_signal_10112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2291 ( .C (clk), .D (new_AGEMA_signal_10115), .Q (new_AGEMA_signal_10116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2295 ( .C (clk), .D (new_AGEMA_signal_10119), .Q (new_AGEMA_signal_10120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2299 ( .C (clk), .D (new_AGEMA_signal_10123), .Q (new_AGEMA_signal_10124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2303 ( .C (clk), .D (new_AGEMA_signal_10127), .Q (new_AGEMA_signal_10128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2307 ( .C (clk), .D (new_AGEMA_signal_10131), .Q (new_AGEMA_signal_10132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2311 ( .C (clk), .D (new_AGEMA_signal_10135), .Q (new_AGEMA_signal_10136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2315 ( .C (clk), .D (new_AGEMA_signal_10139), .Q (new_AGEMA_signal_10140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2319 ( .C (clk), .D (new_AGEMA_signal_10143), .Q (new_AGEMA_signal_10144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2323 ( .C (clk), .D (new_AGEMA_signal_10147), .Q (new_AGEMA_signal_10148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2327 ( .C (clk), .D (new_AGEMA_signal_10151), .Q (new_AGEMA_signal_10152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2331 ( .C (clk), .D (new_AGEMA_signal_10155), .Q (new_AGEMA_signal_10156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2335 ( .C (clk), .D (new_AGEMA_signal_10159), .Q (new_AGEMA_signal_10160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2339 ( .C (clk), .D (new_AGEMA_signal_10163), .Q (new_AGEMA_signal_10164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2343 ( .C (clk), .D (new_AGEMA_signal_10167), .Q (new_AGEMA_signal_10168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2347 ( .C (clk), .D (new_AGEMA_signal_10171), .Q (new_AGEMA_signal_10172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2351 ( .C (clk), .D (new_AGEMA_signal_10175), .Q (new_AGEMA_signal_10176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2355 ( .C (clk), .D (new_AGEMA_signal_10179), .Q (new_AGEMA_signal_10180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2359 ( .C (clk), .D (new_AGEMA_signal_10183), .Q (new_AGEMA_signal_10184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2363 ( .C (clk), .D (new_AGEMA_signal_10187), .Q (new_AGEMA_signal_10188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2367 ( .C (clk), .D (new_AGEMA_signal_10191), .Q (new_AGEMA_signal_10192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2371 ( .C (clk), .D (new_AGEMA_signal_10195), .Q (new_AGEMA_signal_10196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2375 ( .C (clk), .D (new_AGEMA_signal_10199), .Q (new_AGEMA_signal_10200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2379 ( .C (clk), .D (new_AGEMA_signal_10203), .Q (new_AGEMA_signal_10204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2383 ( .C (clk), .D (new_AGEMA_signal_10207), .Q (new_AGEMA_signal_10208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2387 ( .C (clk), .D (new_AGEMA_signal_10211), .Q (new_AGEMA_signal_10212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2391 ( .C (clk), .D (new_AGEMA_signal_10215), .Q (new_AGEMA_signal_10216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2395 ( .C (clk), .D (new_AGEMA_signal_10219), .Q (new_AGEMA_signal_10220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2399 ( .C (clk), .D (new_AGEMA_signal_10223), .Q (new_AGEMA_signal_10224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2403 ( .C (clk), .D (new_AGEMA_signal_10227), .Q (new_AGEMA_signal_10228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2407 ( .C (clk), .D (new_AGEMA_signal_10231), .Q (new_AGEMA_signal_10232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2411 ( .C (clk), .D (new_AGEMA_signal_10235), .Q (new_AGEMA_signal_10236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2415 ( .C (clk), .D (new_AGEMA_signal_10239), .Q (new_AGEMA_signal_10240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2419 ( .C (clk), .D (new_AGEMA_signal_10243), .Q (new_AGEMA_signal_10244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2423 ( .C (clk), .D (new_AGEMA_signal_10247), .Q (new_AGEMA_signal_10248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2427 ( .C (clk), .D (new_AGEMA_signal_10251), .Q (new_AGEMA_signal_10252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2431 ( .C (clk), .D (new_AGEMA_signal_10255), .Q (new_AGEMA_signal_10256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2435 ( .C (clk), .D (new_AGEMA_signal_10259), .Q (new_AGEMA_signal_10260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2439 ( .C (clk), .D (new_AGEMA_signal_10263), .Q (new_AGEMA_signal_10264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2443 ( .C (clk), .D (new_AGEMA_signal_10267), .Q (new_AGEMA_signal_10268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2447 ( .C (clk), .D (new_AGEMA_signal_10271), .Q (new_AGEMA_signal_10272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2451 ( .C (clk), .D (new_AGEMA_signal_10275), .Q (new_AGEMA_signal_10276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2455 ( .C (clk), .D (new_AGEMA_signal_10279), .Q (new_AGEMA_signal_10280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2459 ( .C (clk), .D (new_AGEMA_signal_10283), .Q (new_AGEMA_signal_10284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2463 ( .C (clk), .D (new_AGEMA_signal_10287), .Q (new_AGEMA_signal_10288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2467 ( .C (clk), .D (new_AGEMA_signal_10291), .Q (new_AGEMA_signal_10292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2471 ( .C (clk), .D (new_AGEMA_signal_10295), .Q (new_AGEMA_signal_10296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2475 ( .C (clk), .D (new_AGEMA_signal_10299), .Q (new_AGEMA_signal_10300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2479 ( .C (clk), .D (new_AGEMA_signal_10303), .Q (new_AGEMA_signal_10304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2483 ( .C (clk), .D (new_AGEMA_signal_10307), .Q (new_AGEMA_signal_10308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2487 ( .C (clk), .D (new_AGEMA_signal_10311), .Q (new_AGEMA_signal_10312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2491 ( .C (clk), .D (new_AGEMA_signal_10315), .Q (new_AGEMA_signal_10316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2495 ( .C (clk), .D (new_AGEMA_signal_10319), .Q (new_AGEMA_signal_10320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2499 ( .C (clk), .D (new_AGEMA_signal_10323), .Q (new_AGEMA_signal_10324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2503 ( .C (clk), .D (new_AGEMA_signal_10327), .Q (new_AGEMA_signal_10328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2507 ( .C (clk), .D (new_AGEMA_signal_10331), .Q (new_AGEMA_signal_10332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2511 ( .C (clk), .D (new_AGEMA_signal_10335), .Q (new_AGEMA_signal_10336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2515 ( .C (clk), .D (new_AGEMA_signal_10339), .Q (new_AGEMA_signal_10340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2519 ( .C (clk), .D (new_AGEMA_signal_10343), .Q (new_AGEMA_signal_10344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2523 ( .C (clk), .D (new_AGEMA_signal_10347), .Q (new_AGEMA_signal_10348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2527 ( .C (clk), .D (new_AGEMA_signal_10351), .Q (new_AGEMA_signal_10352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2531 ( .C (clk), .D (new_AGEMA_signal_10355), .Q (new_AGEMA_signal_10356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2535 ( .C (clk), .D (new_AGEMA_signal_10359), .Q (new_AGEMA_signal_10360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2539 ( .C (clk), .D (new_AGEMA_signal_10363), .Q (new_AGEMA_signal_10364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2543 ( .C (clk), .D (new_AGEMA_signal_10367), .Q (new_AGEMA_signal_10368) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2547 ( .C (clk), .D (new_AGEMA_signal_10371), .Q (new_AGEMA_signal_10372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2551 ( .C (clk), .D (new_AGEMA_signal_10375), .Q (new_AGEMA_signal_10376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2555 ( .C (clk), .D (new_AGEMA_signal_10379), .Q (new_AGEMA_signal_10380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2559 ( .C (clk), .D (new_AGEMA_signal_10383), .Q (new_AGEMA_signal_10384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2563 ( .C (clk), .D (new_AGEMA_signal_10387), .Q (new_AGEMA_signal_10388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2567 ( .C (clk), .D (new_AGEMA_signal_10391), .Q (new_AGEMA_signal_10392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2571 ( .C (clk), .D (new_AGEMA_signal_10395), .Q (new_AGEMA_signal_10396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2575 ( .C (clk), .D (new_AGEMA_signal_10399), .Q (new_AGEMA_signal_10400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2579 ( .C (clk), .D (new_AGEMA_signal_10403), .Q (new_AGEMA_signal_10404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2583 ( .C (clk), .D (new_AGEMA_signal_10407), .Q (new_AGEMA_signal_10408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2587 ( .C (clk), .D (new_AGEMA_signal_10411), .Q (new_AGEMA_signal_10412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2591 ( .C (clk), .D (new_AGEMA_signal_10415), .Q (new_AGEMA_signal_10416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2595 ( .C (clk), .D (new_AGEMA_signal_10419), .Q (new_AGEMA_signal_10420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2599 ( .C (clk), .D (new_AGEMA_signal_10423), .Q (new_AGEMA_signal_10424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2603 ( .C (clk), .D (new_AGEMA_signal_10427), .Q (new_AGEMA_signal_10428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2607 ( .C (clk), .D (new_AGEMA_signal_10431), .Q (new_AGEMA_signal_10432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2611 ( .C (clk), .D (new_AGEMA_signal_10435), .Q (new_AGEMA_signal_10436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2615 ( .C (clk), .D (new_AGEMA_signal_10439), .Q (new_AGEMA_signal_10440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2619 ( .C (clk), .D (new_AGEMA_signal_10443), .Q (new_AGEMA_signal_10444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2623 ( .C (clk), .D (new_AGEMA_signal_10447), .Q (new_AGEMA_signal_10448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2627 ( .C (clk), .D (new_AGEMA_signal_10451), .Q (new_AGEMA_signal_10452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2631 ( .C (clk), .D (new_AGEMA_signal_10455), .Q (new_AGEMA_signal_10456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2635 ( .C (clk), .D (new_AGEMA_signal_10459), .Q (new_AGEMA_signal_10460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2639 ( .C (clk), .D (new_AGEMA_signal_10463), .Q (new_AGEMA_signal_10464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2643 ( .C (clk), .D (new_AGEMA_signal_10467), .Q (new_AGEMA_signal_10468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2647 ( .C (clk), .D (new_AGEMA_signal_10471), .Q (new_AGEMA_signal_10472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2651 ( .C (clk), .D (new_AGEMA_signal_10475), .Q (new_AGEMA_signal_10476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2655 ( .C (clk), .D (new_AGEMA_signal_10479), .Q (new_AGEMA_signal_10480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2659 ( .C (clk), .D (new_AGEMA_signal_10483), .Q (new_AGEMA_signal_10484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2663 ( .C (clk), .D (new_AGEMA_signal_10487), .Q (new_AGEMA_signal_10488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2667 ( .C (clk), .D (new_AGEMA_signal_10491), .Q (new_AGEMA_signal_10492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2671 ( .C (clk), .D (new_AGEMA_signal_10495), .Q (new_AGEMA_signal_10496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2675 ( .C (clk), .D (new_AGEMA_signal_10499), .Q (new_AGEMA_signal_10500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2679 ( .C (clk), .D (new_AGEMA_signal_10503), .Q (new_AGEMA_signal_10504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2683 ( .C (clk), .D (new_AGEMA_signal_10507), .Q (new_AGEMA_signal_10508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2687 ( .C (clk), .D (new_AGEMA_signal_10511), .Q (new_AGEMA_signal_10512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2691 ( .C (clk), .D (new_AGEMA_signal_10515), .Q (new_AGEMA_signal_10516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2695 ( .C (clk), .D (new_AGEMA_signal_10519), .Q (new_AGEMA_signal_10520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2699 ( .C (clk), .D (new_AGEMA_signal_10523), .Q (new_AGEMA_signal_10524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2703 ( .C (clk), .D (new_AGEMA_signal_10527), .Q (new_AGEMA_signal_10528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2707 ( .C (clk), .D (new_AGEMA_signal_10531), .Q (new_AGEMA_signal_10532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2711 ( .C (clk), .D (new_AGEMA_signal_10535), .Q (new_AGEMA_signal_10536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2715 ( .C (clk), .D (new_AGEMA_signal_10539), .Q (new_AGEMA_signal_10540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2719 ( .C (clk), .D (new_AGEMA_signal_10543), .Q (new_AGEMA_signal_10544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2723 ( .C (clk), .D (new_AGEMA_signal_10547), .Q (new_AGEMA_signal_10548) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2727 ( .C (clk), .D (new_AGEMA_signal_10551), .Q (new_AGEMA_signal_10552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2731 ( .C (clk), .D (new_AGEMA_signal_10555), .Q (new_AGEMA_signal_10556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2735 ( .C (clk), .D (new_AGEMA_signal_10559), .Q (new_AGEMA_signal_10560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2739 ( .C (clk), .D (new_AGEMA_signal_10563), .Q (new_AGEMA_signal_10564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2743 ( .C (clk), .D (new_AGEMA_signal_10567), .Q (new_AGEMA_signal_10568) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2747 ( .C (clk), .D (new_AGEMA_signal_10571), .Q (new_AGEMA_signal_10572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2751 ( .C (clk), .D (new_AGEMA_signal_10575), .Q (new_AGEMA_signal_10576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2755 ( .C (clk), .D (new_AGEMA_signal_10579), .Q (new_AGEMA_signal_10580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2759 ( .C (clk), .D (new_AGEMA_signal_10583), .Q (new_AGEMA_signal_10584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2763 ( .C (clk), .D (new_AGEMA_signal_10587), .Q (new_AGEMA_signal_10588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2767 ( .C (clk), .D (new_AGEMA_signal_10591), .Q (new_AGEMA_signal_10592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2771 ( .C (clk), .D (new_AGEMA_signal_10595), .Q (new_AGEMA_signal_10596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2774 ( .C (clk), .D (new_AGEMA_signal_10598), .Q (new_AGEMA_signal_10599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2777 ( .C (clk), .D (new_AGEMA_signal_10601), .Q (new_AGEMA_signal_10602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2780 ( .C (clk), .D (new_AGEMA_signal_10604), .Q (new_AGEMA_signal_10605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2783 ( .C (clk), .D (new_AGEMA_signal_10607), .Q (new_AGEMA_signal_10608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2786 ( .C (clk), .D (new_AGEMA_signal_10610), .Q (new_AGEMA_signal_10611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2789 ( .C (clk), .D (new_AGEMA_signal_10613), .Q (new_AGEMA_signal_10614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2792 ( .C (clk), .D (new_AGEMA_signal_10616), .Q (new_AGEMA_signal_10617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2795 ( .C (clk), .D (new_AGEMA_signal_10619), .Q (new_AGEMA_signal_10620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2798 ( .C (clk), .D (new_AGEMA_signal_10622), .Q (new_AGEMA_signal_10623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2801 ( .C (clk), .D (new_AGEMA_signal_10625), .Q (new_AGEMA_signal_10626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2804 ( .C (clk), .D (new_AGEMA_signal_10628), .Q (new_AGEMA_signal_10629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2807 ( .C (clk), .D (new_AGEMA_signal_10631), .Q (new_AGEMA_signal_10632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2810 ( .C (clk), .D (new_AGEMA_signal_10634), .Q (new_AGEMA_signal_10635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2813 ( .C (clk), .D (new_AGEMA_signal_10637), .Q (new_AGEMA_signal_10638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2816 ( .C (clk), .D (new_AGEMA_signal_10640), .Q (new_AGEMA_signal_10641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2819 ( .C (clk), .D (new_AGEMA_signal_10643), .Q (new_AGEMA_signal_10644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2822 ( .C (clk), .D (new_AGEMA_signal_10646), .Q (new_AGEMA_signal_10647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2825 ( .C (clk), .D (new_AGEMA_signal_10649), .Q (new_AGEMA_signal_10650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2828 ( .C (clk), .D (new_AGEMA_signal_10652), .Q (new_AGEMA_signal_10653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2831 ( .C (clk), .D (new_AGEMA_signal_10655), .Q (new_AGEMA_signal_10656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2834 ( .C (clk), .D (new_AGEMA_signal_10658), .Q (new_AGEMA_signal_10659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2837 ( .C (clk), .D (new_AGEMA_signal_10661), .Q (new_AGEMA_signal_10662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2840 ( .C (clk), .D (new_AGEMA_signal_10664), .Q (new_AGEMA_signal_10665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2843 ( .C (clk), .D (new_AGEMA_signal_10667), .Q (new_AGEMA_signal_10668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2846 ( .C (clk), .D (new_AGEMA_signal_10670), .Q (new_AGEMA_signal_10671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2849 ( .C (clk), .D (new_AGEMA_signal_10673), .Q (new_AGEMA_signal_10674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2852 ( .C (clk), .D (new_AGEMA_signal_10676), .Q (new_AGEMA_signal_10677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2855 ( .C (clk), .D (new_AGEMA_signal_10679), .Q (new_AGEMA_signal_10680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2858 ( .C (clk), .D (new_AGEMA_signal_10682), .Q (new_AGEMA_signal_10683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2861 ( .C (clk), .D (new_AGEMA_signal_10685), .Q (new_AGEMA_signal_10686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2864 ( .C (clk), .D (new_AGEMA_signal_10688), .Q (new_AGEMA_signal_10689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2867 ( .C (clk), .D (new_AGEMA_signal_10691), .Q (new_AGEMA_signal_10692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2870 ( .C (clk), .D (new_AGEMA_signal_10694), .Q (new_AGEMA_signal_10695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2873 ( .C (clk), .D (new_AGEMA_signal_10697), .Q (new_AGEMA_signal_10698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2876 ( .C (clk), .D (new_AGEMA_signal_10700), .Q (new_AGEMA_signal_10701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2879 ( .C (clk), .D (new_AGEMA_signal_10703), .Q (new_AGEMA_signal_10704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2882 ( .C (clk), .D (new_AGEMA_signal_10706), .Q (new_AGEMA_signal_10707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2885 ( .C (clk), .D (new_AGEMA_signal_10709), .Q (new_AGEMA_signal_10710) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2888 ( .C (clk), .D (new_AGEMA_signal_10712), .Q (new_AGEMA_signal_10713) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2891 ( .C (clk), .D (new_AGEMA_signal_10715), .Q (new_AGEMA_signal_10716) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2894 ( .C (clk), .D (new_AGEMA_signal_10718), .Q (new_AGEMA_signal_10719) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2897 ( .C (clk), .D (new_AGEMA_signal_10721), .Q (new_AGEMA_signal_10722) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2900 ( .C (clk), .D (new_AGEMA_signal_10724), .Q (new_AGEMA_signal_10725) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2903 ( .C (clk), .D (new_AGEMA_signal_10727), .Q (new_AGEMA_signal_10728) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2906 ( .C (clk), .D (new_AGEMA_signal_10730), .Q (new_AGEMA_signal_10731) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2909 ( .C (clk), .D (new_AGEMA_signal_10733), .Q (new_AGEMA_signal_10734) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2912 ( .C (clk), .D (new_AGEMA_signal_10736), .Q (new_AGEMA_signal_10737) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2915 ( .C (clk), .D (new_AGEMA_signal_10739), .Q (new_AGEMA_signal_10740) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2918 ( .C (clk), .D (new_AGEMA_signal_10742), .Q (new_AGEMA_signal_10743) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2921 ( .C (clk), .D (new_AGEMA_signal_10745), .Q (new_AGEMA_signal_10746) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2924 ( .C (clk), .D (new_AGEMA_signal_10748), .Q (new_AGEMA_signal_10749) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2927 ( .C (clk), .D (new_AGEMA_signal_10751), .Q (new_AGEMA_signal_10752) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2930 ( .C (clk), .D (new_AGEMA_signal_10754), .Q (new_AGEMA_signal_10755) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2933 ( .C (clk), .D (new_AGEMA_signal_10757), .Q (new_AGEMA_signal_10758) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2936 ( .C (clk), .D (new_AGEMA_signal_10760), .Q (new_AGEMA_signal_10761) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2939 ( .C (clk), .D (new_AGEMA_signal_10763), .Q (new_AGEMA_signal_10764) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2942 ( .C (clk), .D (new_AGEMA_signal_10766), .Q (new_AGEMA_signal_10767) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2945 ( .C (clk), .D (new_AGEMA_signal_10769), .Q (new_AGEMA_signal_10770) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2948 ( .C (clk), .D (new_AGEMA_signal_10772), .Q (new_AGEMA_signal_10773) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2951 ( .C (clk), .D (new_AGEMA_signal_10775), .Q (new_AGEMA_signal_10776) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2954 ( .C (clk), .D (new_AGEMA_signal_10778), .Q (new_AGEMA_signal_10779) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2957 ( .C (clk), .D (new_AGEMA_signal_10781), .Q (new_AGEMA_signal_10782) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2960 ( .C (clk), .D (new_AGEMA_signal_10784), .Q (new_AGEMA_signal_10785) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2963 ( .C (clk), .D (new_AGEMA_signal_10787), .Q (new_AGEMA_signal_10788) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2966 ( .C (clk), .D (new_AGEMA_signal_10790), .Q (new_AGEMA_signal_10791) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2969 ( .C (clk), .D (new_AGEMA_signal_10793), .Q (new_AGEMA_signal_10794) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2972 ( .C (clk), .D (new_AGEMA_signal_10796), .Q (new_AGEMA_signal_10797) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2975 ( .C (clk), .D (new_AGEMA_signal_10799), .Q (new_AGEMA_signal_10800) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2978 ( .C (clk), .D (new_AGEMA_signal_10802), .Q (new_AGEMA_signal_10803) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2981 ( .C (clk), .D (new_AGEMA_signal_10805), .Q (new_AGEMA_signal_10806) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2984 ( .C (clk), .D (new_AGEMA_signal_10808), .Q (new_AGEMA_signal_10809) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2987 ( .C (clk), .D (new_AGEMA_signal_10811), .Q (new_AGEMA_signal_10812) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2990 ( .C (clk), .D (new_AGEMA_signal_10814), .Q (new_AGEMA_signal_10815) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2993 ( .C (clk), .D (new_AGEMA_signal_10817), .Q (new_AGEMA_signal_10818) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2996 ( .C (clk), .D (new_AGEMA_signal_10820), .Q (new_AGEMA_signal_10821) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2999 ( .C (clk), .D (new_AGEMA_signal_10823), .Q (new_AGEMA_signal_10824) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3002 ( .C (clk), .D (new_AGEMA_signal_10826), .Q (new_AGEMA_signal_10827) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3005 ( .C (clk), .D (new_AGEMA_signal_10829), .Q (new_AGEMA_signal_10830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3008 ( .C (clk), .D (new_AGEMA_signal_10832), .Q (new_AGEMA_signal_10833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3011 ( .C (clk), .D (new_AGEMA_signal_10835), .Q (new_AGEMA_signal_10836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3014 ( .C (clk), .D (new_AGEMA_signal_10838), .Q (new_AGEMA_signal_10839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3017 ( .C (clk), .D (new_AGEMA_signal_10841), .Q (new_AGEMA_signal_10842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3020 ( .C (clk), .D (new_AGEMA_signal_10844), .Q (new_AGEMA_signal_10845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3023 ( .C (clk), .D (new_AGEMA_signal_10847), .Q (new_AGEMA_signal_10848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3026 ( .C (clk), .D (new_AGEMA_signal_10850), .Q (new_AGEMA_signal_10851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3029 ( .C (clk), .D (new_AGEMA_signal_10853), .Q (new_AGEMA_signal_10854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3032 ( .C (clk), .D (new_AGEMA_signal_10856), .Q (new_AGEMA_signal_10857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3035 ( .C (clk), .D (new_AGEMA_signal_10859), .Q (new_AGEMA_signal_10860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3038 ( .C (clk), .D (new_AGEMA_signal_10862), .Q (new_AGEMA_signal_10863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3041 ( .C (clk), .D (new_AGEMA_signal_10865), .Q (new_AGEMA_signal_10866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3044 ( .C (clk), .D (new_AGEMA_signal_10868), .Q (new_AGEMA_signal_10869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3047 ( .C (clk), .D (new_AGEMA_signal_10871), .Q (new_AGEMA_signal_10872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3050 ( .C (clk), .D (new_AGEMA_signal_10874), .Q (new_AGEMA_signal_10875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3053 ( .C (clk), .D (new_AGEMA_signal_10877), .Q (new_AGEMA_signal_10878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3056 ( .C (clk), .D (new_AGEMA_signal_10880), .Q (new_AGEMA_signal_10881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3059 ( .C (clk), .D (new_AGEMA_signal_10883), .Q (new_AGEMA_signal_10884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3062 ( .C (clk), .D (new_AGEMA_signal_10886), .Q (new_AGEMA_signal_10887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3065 ( .C (clk), .D (new_AGEMA_signal_10889), .Q (new_AGEMA_signal_10890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3068 ( .C (clk), .D (new_AGEMA_signal_10892), .Q (new_AGEMA_signal_10893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3071 ( .C (clk), .D (new_AGEMA_signal_10895), .Q (new_AGEMA_signal_10896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3074 ( .C (clk), .D (new_AGEMA_signal_10898), .Q (new_AGEMA_signal_10899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3077 ( .C (clk), .D (new_AGEMA_signal_10901), .Q (new_AGEMA_signal_10902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3080 ( .C (clk), .D (new_AGEMA_signal_10904), .Q (new_AGEMA_signal_10905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3083 ( .C (clk), .D (new_AGEMA_signal_10907), .Q (new_AGEMA_signal_10908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3086 ( .C (clk), .D (new_AGEMA_signal_10910), .Q (new_AGEMA_signal_10911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3089 ( .C (clk), .D (new_AGEMA_signal_10913), .Q (new_AGEMA_signal_10914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3092 ( .C (clk), .D (new_AGEMA_signal_10916), .Q (new_AGEMA_signal_10917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3095 ( .C (clk), .D (new_AGEMA_signal_10919), .Q (new_AGEMA_signal_10920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3098 ( .C (clk), .D (new_AGEMA_signal_10922), .Q (new_AGEMA_signal_10923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3101 ( .C (clk), .D (new_AGEMA_signal_10925), .Q (new_AGEMA_signal_10926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3104 ( .C (clk), .D (new_AGEMA_signal_10928), .Q (new_AGEMA_signal_10929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3107 ( .C (clk), .D (new_AGEMA_signal_10931), .Q (new_AGEMA_signal_10932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3110 ( .C (clk), .D (new_AGEMA_signal_10934), .Q (new_AGEMA_signal_10935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3113 ( .C (clk), .D (new_AGEMA_signal_10937), .Q (new_AGEMA_signal_10938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3116 ( .C (clk), .D (new_AGEMA_signal_10940), .Q (new_AGEMA_signal_10941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3119 ( .C (clk), .D (new_AGEMA_signal_10943), .Q (new_AGEMA_signal_10944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3122 ( .C (clk), .D (new_AGEMA_signal_10946), .Q (new_AGEMA_signal_10947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3125 ( .C (clk), .D (new_AGEMA_signal_10949), .Q (new_AGEMA_signal_10950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3128 ( .C (clk), .D (new_AGEMA_signal_10952), .Q (new_AGEMA_signal_10953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3131 ( .C (clk), .D (new_AGEMA_signal_10955), .Q (new_AGEMA_signal_10956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3134 ( .C (clk), .D (new_AGEMA_signal_10958), .Q (new_AGEMA_signal_10959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3137 ( .C (clk), .D (new_AGEMA_signal_10961), .Q (new_AGEMA_signal_10962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3140 ( .C (clk), .D (new_AGEMA_signal_10964), .Q (new_AGEMA_signal_10965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3143 ( .C (clk), .D (new_AGEMA_signal_10967), .Q (new_AGEMA_signal_10968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3146 ( .C (clk), .D (new_AGEMA_signal_10970), .Q (new_AGEMA_signal_10971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3149 ( .C (clk), .D (new_AGEMA_signal_10973), .Q (new_AGEMA_signal_10974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3152 ( .C (clk), .D (new_AGEMA_signal_10976), .Q (new_AGEMA_signal_10977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3155 ( .C (clk), .D (new_AGEMA_signal_10979), .Q (new_AGEMA_signal_10980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3158 ( .C (clk), .D (new_AGEMA_signal_10982), .Q (new_AGEMA_signal_10983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3161 ( .C (clk), .D (new_AGEMA_signal_10985), .Q (new_AGEMA_signal_10986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3164 ( .C (clk), .D (new_AGEMA_signal_10988), .Q (new_AGEMA_signal_10989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3167 ( .C (clk), .D (new_AGEMA_signal_10991), .Q (new_AGEMA_signal_10992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3170 ( .C (clk), .D (new_AGEMA_signal_10994), .Q (new_AGEMA_signal_10995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3173 ( .C (clk), .D (new_AGEMA_signal_10997), .Q (new_AGEMA_signal_10998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3176 ( .C (clk), .D (new_AGEMA_signal_11000), .Q (new_AGEMA_signal_11001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3179 ( .C (clk), .D (new_AGEMA_signal_11003), .Q (new_AGEMA_signal_11004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3182 ( .C (clk), .D (new_AGEMA_signal_11006), .Q (new_AGEMA_signal_11007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3185 ( .C (clk), .D (new_AGEMA_signal_11009), .Q (new_AGEMA_signal_11010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3188 ( .C (clk), .D (new_AGEMA_signal_11012), .Q (new_AGEMA_signal_11013) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3191 ( .C (clk), .D (new_AGEMA_signal_11015), .Q (new_AGEMA_signal_11016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3194 ( .C (clk), .D (new_AGEMA_signal_11018), .Q (new_AGEMA_signal_11019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3197 ( .C (clk), .D (new_AGEMA_signal_11021), .Q (new_AGEMA_signal_11022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3200 ( .C (clk), .D (new_AGEMA_signal_11024), .Q (new_AGEMA_signal_11025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3203 ( .C (clk), .D (new_AGEMA_signal_11027), .Q (new_AGEMA_signal_11028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3206 ( .C (clk), .D (new_AGEMA_signal_11030), .Q (new_AGEMA_signal_11031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3209 ( .C (clk), .D (new_AGEMA_signal_11033), .Q (new_AGEMA_signal_11034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3212 ( .C (clk), .D (new_AGEMA_signal_11036), .Q (new_AGEMA_signal_11037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3215 ( .C (clk), .D (new_AGEMA_signal_11039), .Q (new_AGEMA_signal_11040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3218 ( .C (clk), .D (new_AGEMA_signal_11042), .Q (new_AGEMA_signal_11043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3221 ( .C (clk), .D (new_AGEMA_signal_11045), .Q (new_AGEMA_signal_11046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3224 ( .C (clk), .D (new_AGEMA_signal_11048), .Q (new_AGEMA_signal_11049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3227 ( .C (clk), .D (new_AGEMA_signal_11051), .Q (new_AGEMA_signal_11052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3230 ( .C (clk), .D (new_AGEMA_signal_11054), .Q (new_AGEMA_signal_11055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3233 ( .C (clk), .D (new_AGEMA_signal_11057), .Q (new_AGEMA_signal_11058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3236 ( .C (clk), .D (new_AGEMA_signal_11060), .Q (new_AGEMA_signal_11061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3239 ( .C (clk), .D (new_AGEMA_signal_11063), .Q (new_AGEMA_signal_11064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3242 ( .C (clk), .D (new_AGEMA_signal_11066), .Q (new_AGEMA_signal_11067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3245 ( .C (clk), .D (new_AGEMA_signal_11069), .Q (new_AGEMA_signal_11070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3248 ( .C (clk), .D (new_AGEMA_signal_11072), .Q (new_AGEMA_signal_11073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3251 ( .C (clk), .D (new_AGEMA_signal_11075), .Q (new_AGEMA_signal_11076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3254 ( .C (clk), .D (new_AGEMA_signal_11078), .Q (new_AGEMA_signal_11079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3257 ( .C (clk), .D (new_AGEMA_signal_11081), .Q (new_AGEMA_signal_11082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3260 ( .C (clk), .D (new_AGEMA_signal_11084), .Q (new_AGEMA_signal_11085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3263 ( .C (clk), .D (new_AGEMA_signal_11087), .Q (new_AGEMA_signal_11088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3266 ( .C (clk), .D (new_AGEMA_signal_11090), .Q (new_AGEMA_signal_11091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3269 ( .C (clk), .D (new_AGEMA_signal_11093), .Q (new_AGEMA_signal_11094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3272 ( .C (clk), .D (new_AGEMA_signal_11096), .Q (new_AGEMA_signal_11097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3275 ( .C (clk), .D (new_AGEMA_signal_11099), .Q (new_AGEMA_signal_11100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3278 ( .C (clk), .D (new_AGEMA_signal_11102), .Q (new_AGEMA_signal_11103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3281 ( .C (clk), .D (new_AGEMA_signal_11105), .Q (new_AGEMA_signal_11106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3284 ( .C (clk), .D (new_AGEMA_signal_11108), .Q (new_AGEMA_signal_11109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3287 ( .C (clk), .D (new_AGEMA_signal_11111), .Q (new_AGEMA_signal_11112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3290 ( .C (clk), .D (new_AGEMA_signal_11114), .Q (new_AGEMA_signal_11115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3293 ( .C (clk), .D (new_AGEMA_signal_11117), .Q (new_AGEMA_signal_11118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3296 ( .C (clk), .D (new_AGEMA_signal_11120), .Q (new_AGEMA_signal_11121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3299 ( .C (clk), .D (new_AGEMA_signal_11123), .Q (new_AGEMA_signal_11124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3302 ( .C (clk), .D (new_AGEMA_signal_11126), .Q (new_AGEMA_signal_11127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3305 ( .C (clk), .D (new_AGEMA_signal_11129), .Q (new_AGEMA_signal_11130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3308 ( .C (clk), .D (new_AGEMA_signal_11132), .Q (new_AGEMA_signal_11133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3311 ( .C (clk), .D (new_AGEMA_signal_11135), .Q (new_AGEMA_signal_11136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3314 ( .C (clk), .D (new_AGEMA_signal_11138), .Q (new_AGEMA_signal_11139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3317 ( .C (clk), .D (new_AGEMA_signal_11141), .Q (new_AGEMA_signal_11142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3320 ( .C (clk), .D (new_AGEMA_signal_11144), .Q (new_AGEMA_signal_11145) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3323 ( .C (clk), .D (new_AGEMA_signal_11147), .Q (new_AGEMA_signal_11148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3326 ( .C (clk), .D (new_AGEMA_signal_11150), .Q (new_AGEMA_signal_11151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3329 ( .C (clk), .D (new_AGEMA_signal_11153), .Q (new_AGEMA_signal_11154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3332 ( .C (clk), .D (new_AGEMA_signal_11156), .Q (new_AGEMA_signal_11157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3335 ( .C (clk), .D (new_AGEMA_signal_11159), .Q (new_AGEMA_signal_11160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3338 ( .C (clk), .D (new_AGEMA_signal_11162), .Q (new_AGEMA_signal_11163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3341 ( .C (clk), .D (new_AGEMA_signal_11165), .Q (new_AGEMA_signal_11166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3344 ( .C (clk), .D (new_AGEMA_signal_11168), .Q (new_AGEMA_signal_11169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3347 ( .C (clk), .D (new_AGEMA_signal_11171), .Q (new_AGEMA_signal_11172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3350 ( .C (clk), .D (new_AGEMA_signal_11174), .Q (new_AGEMA_signal_11175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3353 ( .C (clk), .D (new_AGEMA_signal_11177), .Q (new_AGEMA_signal_11178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3356 ( .C (clk), .D (new_AGEMA_signal_11180), .Q (new_AGEMA_signal_11181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3359 ( .C (clk), .D (new_AGEMA_signal_11183), .Q (new_AGEMA_signal_11184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3362 ( .C (clk), .D (new_AGEMA_signal_11186), .Q (new_AGEMA_signal_11187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3365 ( .C (clk), .D (new_AGEMA_signal_11189), .Q (new_AGEMA_signal_11190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3368 ( .C (clk), .D (new_AGEMA_signal_11192), .Q (new_AGEMA_signal_11193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3371 ( .C (clk), .D (new_AGEMA_signal_11195), .Q (new_AGEMA_signal_11196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3374 ( .C (clk), .D (new_AGEMA_signal_11198), .Q (new_AGEMA_signal_11199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3377 ( .C (clk), .D (new_AGEMA_signal_11201), .Q (new_AGEMA_signal_11202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3380 ( .C (clk), .D (new_AGEMA_signal_11204), .Q (new_AGEMA_signal_11205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3383 ( .C (clk), .D (new_AGEMA_signal_11207), .Q (new_AGEMA_signal_11208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3386 ( .C (clk), .D (new_AGEMA_signal_11210), .Q (new_AGEMA_signal_11211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3389 ( .C (clk), .D (new_AGEMA_signal_11213), .Q (new_AGEMA_signal_11214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3392 ( .C (clk), .D (new_AGEMA_signal_11216), .Q (new_AGEMA_signal_11217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3395 ( .C (clk), .D (new_AGEMA_signal_11219), .Q (new_AGEMA_signal_11220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3398 ( .C (clk), .D (new_AGEMA_signal_11222), .Q (new_AGEMA_signal_11223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3401 ( .C (clk), .D (new_AGEMA_signal_11225), .Q (new_AGEMA_signal_11226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3404 ( .C (clk), .D (new_AGEMA_signal_11228), .Q (new_AGEMA_signal_11229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3407 ( .C (clk), .D (new_AGEMA_signal_11231), .Q (new_AGEMA_signal_11232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3410 ( .C (clk), .D (new_AGEMA_signal_11234), .Q (new_AGEMA_signal_11235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3413 ( .C (clk), .D (new_AGEMA_signal_11237), .Q (new_AGEMA_signal_11238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3416 ( .C (clk), .D (new_AGEMA_signal_11240), .Q (new_AGEMA_signal_11241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3419 ( .C (clk), .D (new_AGEMA_signal_11243), .Q (new_AGEMA_signal_11244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3422 ( .C (clk), .D (new_AGEMA_signal_11246), .Q (new_AGEMA_signal_11247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3425 ( .C (clk), .D (new_AGEMA_signal_11249), .Q (new_AGEMA_signal_11250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3428 ( .C (clk), .D (new_AGEMA_signal_11252), .Q (new_AGEMA_signal_11253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3431 ( .C (clk), .D (new_AGEMA_signal_11255), .Q (new_AGEMA_signal_11256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3434 ( .C (clk), .D (new_AGEMA_signal_11258), .Q (new_AGEMA_signal_11259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3437 ( .C (clk), .D (new_AGEMA_signal_11261), .Q (new_AGEMA_signal_11262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3440 ( .C (clk), .D (new_AGEMA_signal_11264), .Q (new_AGEMA_signal_11265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3443 ( .C (clk), .D (new_AGEMA_signal_11267), .Q (new_AGEMA_signal_11268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3446 ( .C (clk), .D (new_AGEMA_signal_11270), .Q (new_AGEMA_signal_11271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3449 ( .C (clk), .D (new_AGEMA_signal_11273), .Q (new_AGEMA_signal_11274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3452 ( .C (clk), .D (new_AGEMA_signal_11276), .Q (new_AGEMA_signal_11277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3455 ( .C (clk), .D (new_AGEMA_signal_11279), .Q (new_AGEMA_signal_11280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3458 ( .C (clk), .D (new_AGEMA_signal_11282), .Q (new_AGEMA_signal_11283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3461 ( .C (clk), .D (new_AGEMA_signal_11285), .Q (new_AGEMA_signal_11286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3464 ( .C (clk), .D (new_AGEMA_signal_11288), .Q (new_AGEMA_signal_11289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3467 ( .C (clk), .D (new_AGEMA_signal_11291), .Q (new_AGEMA_signal_11292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3470 ( .C (clk), .D (new_AGEMA_signal_11294), .Q (new_AGEMA_signal_11295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3473 ( .C (clk), .D (new_AGEMA_signal_11297), .Q (new_AGEMA_signal_11298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3476 ( .C (clk), .D (new_AGEMA_signal_11300), .Q (new_AGEMA_signal_11301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3479 ( .C (clk), .D (new_AGEMA_signal_11303), .Q (new_AGEMA_signal_11304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3482 ( .C (clk), .D (new_AGEMA_signal_11306), .Q (new_AGEMA_signal_11307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3485 ( .C (clk), .D (new_AGEMA_signal_11309), .Q (new_AGEMA_signal_11310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3488 ( .C (clk), .D (new_AGEMA_signal_11312), .Q (new_AGEMA_signal_11313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3491 ( .C (clk), .D (new_AGEMA_signal_11315), .Q (new_AGEMA_signal_11316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3494 ( .C (clk), .D (new_AGEMA_signal_11318), .Q (new_AGEMA_signal_11319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3497 ( .C (clk), .D (new_AGEMA_signal_11321), .Q (new_AGEMA_signal_11322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3500 ( .C (clk), .D (new_AGEMA_signal_11324), .Q (new_AGEMA_signal_11325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3503 ( .C (clk), .D (new_AGEMA_signal_11327), .Q (new_AGEMA_signal_11328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3506 ( .C (clk), .D (new_AGEMA_signal_11330), .Q (new_AGEMA_signal_11331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3509 ( .C (clk), .D (new_AGEMA_signal_11333), .Q (new_AGEMA_signal_11334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3512 ( .C (clk), .D (new_AGEMA_signal_11336), .Q (new_AGEMA_signal_11337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3515 ( .C (clk), .D (new_AGEMA_signal_11339), .Q (new_AGEMA_signal_11340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3518 ( .C (clk), .D (new_AGEMA_signal_11342), .Q (new_AGEMA_signal_11343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3521 ( .C (clk), .D (new_AGEMA_signal_11345), .Q (new_AGEMA_signal_11346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3524 ( .C (clk), .D (new_AGEMA_signal_11348), .Q (new_AGEMA_signal_11349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3527 ( .C (clk), .D (new_AGEMA_signal_11351), .Q (new_AGEMA_signal_11352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3530 ( .C (clk), .D (new_AGEMA_signal_11354), .Q (new_AGEMA_signal_11355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3533 ( .C (clk), .D (new_AGEMA_signal_11357), .Q (new_AGEMA_signal_11358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3536 ( .C (clk), .D (new_AGEMA_signal_11360), .Q (new_AGEMA_signal_11361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3539 ( .C (clk), .D (new_AGEMA_signal_11363), .Q (new_AGEMA_signal_11364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3542 ( .C (clk), .D (new_AGEMA_signal_11366), .Q (new_AGEMA_signal_11367) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3545 ( .C (clk), .D (new_AGEMA_signal_11369), .Q (new_AGEMA_signal_11370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3548 ( .C (clk), .D (new_AGEMA_signal_11372), .Q (new_AGEMA_signal_11373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3551 ( .C (clk), .D (new_AGEMA_signal_11375), .Q (new_AGEMA_signal_11376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3554 ( .C (clk), .D (new_AGEMA_signal_11378), .Q (new_AGEMA_signal_11379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3557 ( .C (clk), .D (new_AGEMA_signal_11381), .Q (new_AGEMA_signal_11382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3560 ( .C (clk), .D (new_AGEMA_signal_11384), .Q (new_AGEMA_signal_11385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3563 ( .C (clk), .D (new_AGEMA_signal_11387), .Q (new_AGEMA_signal_11388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3566 ( .C (clk), .D (new_AGEMA_signal_11390), .Q (new_AGEMA_signal_11391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3569 ( .C (clk), .D (new_AGEMA_signal_11393), .Q (new_AGEMA_signal_11394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3572 ( .C (clk), .D (new_AGEMA_signal_11396), .Q (new_AGEMA_signal_11397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3575 ( .C (clk), .D (new_AGEMA_signal_11399), .Q (new_AGEMA_signal_11400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3578 ( .C (clk), .D (new_AGEMA_signal_11402), .Q (new_AGEMA_signal_11403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3581 ( .C (clk), .D (new_AGEMA_signal_11405), .Q (new_AGEMA_signal_11406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3584 ( .C (clk), .D (new_AGEMA_signal_11408), .Q (new_AGEMA_signal_11409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3587 ( .C (clk), .D (new_AGEMA_signal_11411), .Q (new_AGEMA_signal_11412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3590 ( .C (clk), .D (new_AGEMA_signal_11414), .Q (new_AGEMA_signal_11415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3593 ( .C (clk), .D (new_AGEMA_signal_11417), .Q (new_AGEMA_signal_11418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3596 ( .C (clk), .D (new_AGEMA_signal_11420), .Q (new_AGEMA_signal_11421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3599 ( .C (clk), .D (new_AGEMA_signal_11423), .Q (new_AGEMA_signal_11424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3602 ( .C (clk), .D (new_AGEMA_signal_11426), .Q (new_AGEMA_signal_11427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3605 ( .C (clk), .D (new_AGEMA_signal_11429), .Q (new_AGEMA_signal_11430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3608 ( .C (clk), .D (new_AGEMA_signal_11432), .Q (new_AGEMA_signal_11433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3611 ( .C (clk), .D (new_AGEMA_signal_11435), .Q (new_AGEMA_signal_11436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3614 ( .C (clk), .D (new_AGEMA_signal_11438), .Q (new_AGEMA_signal_11439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3617 ( .C (clk), .D (new_AGEMA_signal_11441), .Q (new_AGEMA_signal_11442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3620 ( .C (clk), .D (new_AGEMA_signal_11444), .Q (new_AGEMA_signal_11445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3623 ( .C (clk), .D (new_AGEMA_signal_11447), .Q (new_AGEMA_signal_11448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3626 ( .C (clk), .D (new_AGEMA_signal_11450), .Q (new_AGEMA_signal_11451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3629 ( .C (clk), .D (new_AGEMA_signal_11453), .Q (new_AGEMA_signal_11454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3632 ( .C (clk), .D (new_AGEMA_signal_11456), .Q (new_AGEMA_signal_11457) ) ;
    buf_clk new_AGEMA_reg_buffer_3635 ( .C (clk), .D (new_AGEMA_signal_11459), .Q (new_AGEMA_signal_11460) ) ;
    buf_clk new_AGEMA_reg_buffer_3639 ( .C (clk), .D (new_AGEMA_signal_11463), .Q (new_AGEMA_signal_11464) ) ;
    buf_clk new_AGEMA_reg_buffer_3643 ( .C (clk), .D (new_AGEMA_signal_11467), .Q (new_AGEMA_signal_11468) ) ;
    buf_clk new_AGEMA_reg_buffer_3647 ( .C (clk), .D (new_AGEMA_signal_11471), .Q (new_AGEMA_signal_11472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3651 ( .C (clk), .D (new_AGEMA_signal_11475), .Q (new_AGEMA_signal_11476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3655 ( .C (clk), .D (new_AGEMA_signal_11479), .Q (new_AGEMA_signal_11480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3659 ( .C (clk), .D (new_AGEMA_signal_11483), .Q (new_AGEMA_signal_11484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3663 ( .C (clk), .D (new_AGEMA_signal_11487), .Q (new_AGEMA_signal_11488) ) ;
    buf_clk new_AGEMA_reg_buffer_3667 ( .C (clk), .D (new_AGEMA_signal_11491), .Q (new_AGEMA_signal_11492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3671 ( .C (clk), .D (new_AGEMA_signal_11495), .Q (new_AGEMA_signal_11496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3675 ( .C (clk), .D (new_AGEMA_signal_11499), .Q (new_AGEMA_signal_11500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3679 ( .C (clk), .D (new_AGEMA_signal_11503), .Q (new_AGEMA_signal_11504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3683 ( .C (clk), .D (new_AGEMA_signal_11507), .Q (new_AGEMA_signal_11508) ) ;
    buf_clk new_AGEMA_reg_buffer_3687 ( .C (clk), .D (new_AGEMA_signal_11511), .Q (new_AGEMA_signal_11512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3691 ( .C (clk), .D (new_AGEMA_signal_11515), .Q (new_AGEMA_signal_11516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3695 ( .C (clk), .D (new_AGEMA_signal_11519), .Q (new_AGEMA_signal_11520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3699 ( .C (clk), .D (new_AGEMA_signal_11523), .Q (new_AGEMA_signal_11524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3703 ( .C (clk), .D (new_AGEMA_signal_11527), .Q (new_AGEMA_signal_11528) ) ;
    buf_clk new_AGEMA_reg_buffer_3707 ( .C (clk), .D (new_AGEMA_signal_11531), .Q (new_AGEMA_signal_11532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3711 ( .C (clk), .D (new_AGEMA_signal_11535), .Q (new_AGEMA_signal_11536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3715 ( .C (clk), .D (new_AGEMA_signal_11539), .Q (new_AGEMA_signal_11540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3719 ( .C (clk), .D (new_AGEMA_signal_11543), .Q (new_AGEMA_signal_11544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3723 ( .C (clk), .D (new_AGEMA_signal_11547), .Q (new_AGEMA_signal_11548) ) ;
    buf_clk new_AGEMA_reg_buffer_3727 ( .C (clk), .D (new_AGEMA_signal_11551), .Q (new_AGEMA_signal_11552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3731 ( .C (clk), .D (new_AGEMA_signal_11555), .Q (new_AGEMA_signal_11556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3735 ( .C (clk), .D (new_AGEMA_signal_11559), .Q (new_AGEMA_signal_11560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3739 ( .C (clk), .D (new_AGEMA_signal_11563), .Q (new_AGEMA_signal_11564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3743 ( .C (clk), .D (new_AGEMA_signal_11567), .Q (new_AGEMA_signal_11568) ) ;
    buf_clk new_AGEMA_reg_buffer_3747 ( .C (clk), .D (new_AGEMA_signal_11571), .Q (new_AGEMA_signal_11572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3751 ( .C (clk), .D (new_AGEMA_signal_11575), .Q (new_AGEMA_signal_11576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3755 ( .C (clk), .D (new_AGEMA_signal_11579), .Q (new_AGEMA_signal_11580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3759 ( .C (clk), .D (new_AGEMA_signal_11583), .Q (new_AGEMA_signal_11584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3763 ( .C (clk), .D (new_AGEMA_signal_11587), .Q (new_AGEMA_signal_11588) ) ;
    buf_clk new_AGEMA_reg_buffer_3767 ( .C (clk), .D (new_AGEMA_signal_11591), .Q (new_AGEMA_signal_11592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3771 ( .C (clk), .D (new_AGEMA_signal_11595), .Q (new_AGEMA_signal_11596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3775 ( .C (clk), .D (new_AGEMA_signal_11599), .Q (new_AGEMA_signal_11600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3779 ( .C (clk), .D (new_AGEMA_signal_11603), .Q (new_AGEMA_signal_11604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3783 ( .C (clk), .D (new_AGEMA_signal_11607), .Q (new_AGEMA_signal_11608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3787 ( .C (clk), .D (new_AGEMA_signal_11611), .Q (new_AGEMA_signal_11612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3791 ( .C (clk), .D (new_AGEMA_signal_11615), .Q (new_AGEMA_signal_11616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3795 ( .C (clk), .D (new_AGEMA_signal_11619), .Q (new_AGEMA_signal_11620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3799 ( .C (clk), .D (new_AGEMA_signal_11623), .Q (new_AGEMA_signal_11624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3803 ( .C (clk), .D (new_AGEMA_signal_11627), .Q (new_AGEMA_signal_11628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3807 ( .C (clk), .D (new_AGEMA_signal_11631), .Q (new_AGEMA_signal_11632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3811 ( .C (clk), .D (new_AGEMA_signal_11635), .Q (new_AGEMA_signal_11636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3815 ( .C (clk), .D (new_AGEMA_signal_11639), .Q (new_AGEMA_signal_11640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3819 ( .C (clk), .D (new_AGEMA_signal_11643), .Q (new_AGEMA_signal_11644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3823 ( .C (clk), .D (new_AGEMA_signal_11647), .Q (new_AGEMA_signal_11648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3827 ( .C (clk), .D (new_AGEMA_signal_11651), .Q (new_AGEMA_signal_11652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3831 ( .C (clk), .D (new_AGEMA_signal_11655), .Q (new_AGEMA_signal_11656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3835 ( .C (clk), .D (new_AGEMA_signal_11659), .Q (new_AGEMA_signal_11660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3839 ( .C (clk), .D (new_AGEMA_signal_11663), .Q (new_AGEMA_signal_11664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3843 ( .C (clk), .D (new_AGEMA_signal_11667), .Q (new_AGEMA_signal_11668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3847 ( .C (clk), .D (new_AGEMA_signal_11671), .Q (new_AGEMA_signal_11672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3851 ( .C (clk), .D (new_AGEMA_signal_11675), .Q (new_AGEMA_signal_11676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3855 ( .C (clk), .D (new_AGEMA_signal_11679), .Q (new_AGEMA_signal_11680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3859 ( .C (clk), .D (new_AGEMA_signal_11683), .Q (new_AGEMA_signal_11684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3863 ( .C (clk), .D (new_AGEMA_signal_11687), .Q (new_AGEMA_signal_11688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3867 ( .C (clk), .D (new_AGEMA_signal_11691), .Q (new_AGEMA_signal_11692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3871 ( .C (clk), .D (new_AGEMA_signal_11695), .Q (new_AGEMA_signal_11696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3875 ( .C (clk), .D (new_AGEMA_signal_11699), .Q (new_AGEMA_signal_11700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3879 ( .C (clk), .D (new_AGEMA_signal_11703), .Q (new_AGEMA_signal_11704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3883 ( .C (clk), .D (new_AGEMA_signal_11707), .Q (new_AGEMA_signal_11708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3887 ( .C (clk), .D (new_AGEMA_signal_11711), .Q (new_AGEMA_signal_11712) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3891 ( .C (clk), .D (new_AGEMA_signal_11715), .Q (new_AGEMA_signal_11716) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3895 ( .C (clk), .D (new_AGEMA_signal_11719), .Q (new_AGEMA_signal_11720) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3899 ( .C (clk), .D (new_AGEMA_signal_11723), .Q (new_AGEMA_signal_11724) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3903 ( .C (clk), .D (new_AGEMA_signal_11727), .Q (new_AGEMA_signal_11728) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3907 ( .C (clk), .D (new_AGEMA_signal_11731), .Q (new_AGEMA_signal_11732) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3911 ( .C (clk), .D (new_AGEMA_signal_11735), .Q (new_AGEMA_signal_11736) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3915 ( .C (clk), .D (new_AGEMA_signal_11739), .Q (new_AGEMA_signal_11740) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3919 ( .C (clk), .D (new_AGEMA_signal_11743), .Q (new_AGEMA_signal_11744) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3923 ( .C (clk), .D (new_AGEMA_signal_11747), .Q (new_AGEMA_signal_11748) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3927 ( .C (clk), .D (new_AGEMA_signal_11751), .Q (new_AGEMA_signal_11752) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3931 ( .C (clk), .D (new_AGEMA_signal_11755), .Q (new_AGEMA_signal_11756) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3935 ( .C (clk), .D (new_AGEMA_signal_11759), .Q (new_AGEMA_signal_11760) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3939 ( .C (clk), .D (new_AGEMA_signal_11763), .Q (new_AGEMA_signal_11764) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3943 ( .C (clk), .D (new_AGEMA_signal_11767), .Q (new_AGEMA_signal_11768) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3947 ( .C (clk), .D (new_AGEMA_signal_11771), .Q (new_AGEMA_signal_11772) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3951 ( .C (clk), .D (new_AGEMA_signal_11775), .Q (new_AGEMA_signal_11776) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3955 ( .C (clk), .D (new_AGEMA_signal_11779), .Q (new_AGEMA_signal_11780) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3959 ( .C (clk), .D (new_AGEMA_signal_11783), .Q (new_AGEMA_signal_11784) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3963 ( .C (clk), .D (new_AGEMA_signal_11787), .Q (new_AGEMA_signal_11788) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3967 ( .C (clk), .D (new_AGEMA_signal_11791), .Q (new_AGEMA_signal_11792) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3971 ( .C (clk), .D (new_AGEMA_signal_11795), .Q (new_AGEMA_signal_11796) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3975 ( .C (clk), .D (new_AGEMA_signal_11799), .Q (new_AGEMA_signal_11800) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3979 ( .C (clk), .D (new_AGEMA_signal_11803), .Q (new_AGEMA_signal_11804) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3983 ( .C (clk), .D (new_AGEMA_signal_11807), .Q (new_AGEMA_signal_11808) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3987 ( .C (clk), .D (new_AGEMA_signal_11811), .Q (new_AGEMA_signal_11812) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3991 ( .C (clk), .D (new_AGEMA_signal_11815), .Q (new_AGEMA_signal_11816) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3995 ( .C (clk), .D (new_AGEMA_signal_11819), .Q (new_AGEMA_signal_11820) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3999 ( .C (clk), .D (new_AGEMA_signal_11823), .Q (new_AGEMA_signal_11824) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4003 ( .C (clk), .D (new_AGEMA_signal_11827), .Q (new_AGEMA_signal_11828) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4007 ( .C (clk), .D (new_AGEMA_signal_11831), .Q (new_AGEMA_signal_11832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4011 ( .C (clk), .D (new_AGEMA_signal_11835), .Q (new_AGEMA_signal_11836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4015 ( .C (clk), .D (new_AGEMA_signal_11839), .Q (new_AGEMA_signal_11840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4019 ( .C (clk), .D (new_AGEMA_signal_11843), .Q (new_AGEMA_signal_11844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4023 ( .C (clk), .D (new_AGEMA_signal_11847), .Q (new_AGEMA_signal_11848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4027 ( .C (clk), .D (new_AGEMA_signal_11851), .Q (new_AGEMA_signal_11852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4031 ( .C (clk), .D (new_AGEMA_signal_11855), .Q (new_AGEMA_signal_11856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4035 ( .C (clk), .D (new_AGEMA_signal_11859), .Q (new_AGEMA_signal_11860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4039 ( .C (clk), .D (new_AGEMA_signal_11863), .Q (new_AGEMA_signal_11864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4043 ( .C (clk), .D (new_AGEMA_signal_11867), .Q (new_AGEMA_signal_11868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4047 ( .C (clk), .D (new_AGEMA_signal_11871), .Q (new_AGEMA_signal_11872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4051 ( .C (clk), .D (new_AGEMA_signal_11875), .Q (new_AGEMA_signal_11876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4055 ( .C (clk), .D (new_AGEMA_signal_11879), .Q (new_AGEMA_signal_11880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4059 ( .C (clk), .D (new_AGEMA_signal_11883), .Q (new_AGEMA_signal_11884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4063 ( .C (clk), .D (new_AGEMA_signal_11887), .Q (new_AGEMA_signal_11888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4067 ( .C (clk), .D (new_AGEMA_signal_11891), .Q (new_AGEMA_signal_11892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4071 ( .C (clk), .D (new_AGEMA_signal_11895), .Q (new_AGEMA_signal_11896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4075 ( .C (clk), .D (new_AGEMA_signal_11899), .Q (new_AGEMA_signal_11900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4079 ( .C (clk), .D (new_AGEMA_signal_11903), .Q (new_AGEMA_signal_11904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4083 ( .C (clk), .D (new_AGEMA_signal_11907), .Q (new_AGEMA_signal_11908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4087 ( .C (clk), .D (new_AGEMA_signal_11911), .Q (new_AGEMA_signal_11912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4091 ( .C (clk), .D (new_AGEMA_signal_11915), .Q (new_AGEMA_signal_11916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4095 ( .C (clk), .D (new_AGEMA_signal_11919), .Q (new_AGEMA_signal_11920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4099 ( .C (clk), .D (new_AGEMA_signal_11923), .Q (new_AGEMA_signal_11924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4103 ( .C (clk), .D (new_AGEMA_signal_11927), .Q (new_AGEMA_signal_11928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4107 ( .C (clk), .D (new_AGEMA_signal_11931), .Q (new_AGEMA_signal_11932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4111 ( .C (clk), .D (new_AGEMA_signal_11935), .Q (new_AGEMA_signal_11936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4115 ( .C (clk), .D (new_AGEMA_signal_11939), .Q (new_AGEMA_signal_11940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4119 ( .C (clk), .D (new_AGEMA_signal_11943), .Q (new_AGEMA_signal_11944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4123 ( .C (clk), .D (new_AGEMA_signal_11947), .Q (new_AGEMA_signal_11948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4127 ( .C (clk), .D (new_AGEMA_signal_11951), .Q (new_AGEMA_signal_11952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4131 ( .C (clk), .D (new_AGEMA_signal_11955), .Q (new_AGEMA_signal_11956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4135 ( .C (clk), .D (new_AGEMA_signal_11959), .Q (new_AGEMA_signal_11960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4139 ( .C (clk), .D (new_AGEMA_signal_11963), .Q (new_AGEMA_signal_11964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4143 ( .C (clk), .D (new_AGEMA_signal_11967), .Q (new_AGEMA_signal_11968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4147 ( .C (clk), .D (new_AGEMA_signal_11971), .Q (new_AGEMA_signal_11972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4151 ( .C (clk), .D (new_AGEMA_signal_11975), .Q (new_AGEMA_signal_11976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4155 ( .C (clk), .D (new_AGEMA_signal_11979), .Q (new_AGEMA_signal_11980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4159 ( .C (clk), .D (new_AGEMA_signal_11983), .Q (new_AGEMA_signal_11984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4163 ( .C (clk), .D (new_AGEMA_signal_11987), .Q (new_AGEMA_signal_11988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4167 ( .C (clk), .D (new_AGEMA_signal_11991), .Q (new_AGEMA_signal_11992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4171 ( .C (clk), .D (new_AGEMA_signal_11995), .Q (new_AGEMA_signal_11996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4175 ( .C (clk), .D (new_AGEMA_signal_11999), .Q (new_AGEMA_signal_12000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4179 ( .C (clk), .D (new_AGEMA_signal_12003), .Q (new_AGEMA_signal_12004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4183 ( .C (clk), .D (new_AGEMA_signal_12007), .Q (new_AGEMA_signal_12008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4187 ( .C (clk), .D (new_AGEMA_signal_12011), .Q (new_AGEMA_signal_12012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4191 ( .C (clk), .D (new_AGEMA_signal_12015), .Q (new_AGEMA_signal_12016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4195 ( .C (clk), .D (new_AGEMA_signal_12019), .Q (new_AGEMA_signal_12020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4199 ( .C (clk), .D (new_AGEMA_signal_12023), .Q (new_AGEMA_signal_12024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4203 ( .C (clk), .D (new_AGEMA_signal_12027), .Q (new_AGEMA_signal_12028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4207 ( .C (clk), .D (new_AGEMA_signal_12031), .Q (new_AGEMA_signal_12032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4211 ( .C (clk), .D (new_AGEMA_signal_12035), .Q (new_AGEMA_signal_12036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4215 ( .C (clk), .D (new_AGEMA_signal_12039), .Q (new_AGEMA_signal_12040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4219 ( .C (clk), .D (new_AGEMA_signal_12043), .Q (new_AGEMA_signal_12044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4223 ( .C (clk), .D (new_AGEMA_signal_12047), .Q (new_AGEMA_signal_12048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4227 ( .C (clk), .D (new_AGEMA_signal_12051), .Q (new_AGEMA_signal_12052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4231 ( .C (clk), .D (new_AGEMA_signal_12055), .Q (new_AGEMA_signal_12056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4235 ( .C (clk), .D (new_AGEMA_signal_12059), .Q (new_AGEMA_signal_12060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4239 ( .C (clk), .D (new_AGEMA_signal_12063), .Q (new_AGEMA_signal_12064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4243 ( .C (clk), .D (new_AGEMA_signal_12067), .Q (new_AGEMA_signal_12068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4247 ( .C (clk), .D (new_AGEMA_signal_12071), .Q (new_AGEMA_signal_12072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4251 ( .C (clk), .D (new_AGEMA_signal_12075), .Q (new_AGEMA_signal_12076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4255 ( .C (clk), .D (new_AGEMA_signal_12079), .Q (new_AGEMA_signal_12080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4259 ( .C (clk), .D (new_AGEMA_signal_12083), .Q (new_AGEMA_signal_12084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4263 ( .C (clk), .D (new_AGEMA_signal_12087), .Q (new_AGEMA_signal_12088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4267 ( .C (clk), .D (new_AGEMA_signal_12091), .Q (new_AGEMA_signal_12092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4271 ( .C (clk), .D (new_AGEMA_signal_12095), .Q (new_AGEMA_signal_12096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4275 ( .C (clk), .D (new_AGEMA_signal_12099), .Q (new_AGEMA_signal_12100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4279 ( .C (clk), .D (new_AGEMA_signal_12103), .Q (new_AGEMA_signal_12104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4283 ( .C (clk), .D (new_AGEMA_signal_12107), .Q (new_AGEMA_signal_12108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4287 ( .C (clk), .D (new_AGEMA_signal_12111), .Q (new_AGEMA_signal_12112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4291 ( .C (clk), .D (new_AGEMA_signal_12115), .Q (new_AGEMA_signal_12116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4295 ( .C (clk), .D (new_AGEMA_signal_12119), .Q (new_AGEMA_signal_12120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4299 ( .C (clk), .D (new_AGEMA_signal_12123), .Q (new_AGEMA_signal_12124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4303 ( .C (clk), .D (new_AGEMA_signal_12127), .Q (new_AGEMA_signal_12128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4307 ( .C (clk), .D (new_AGEMA_signal_12131), .Q (new_AGEMA_signal_12132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4311 ( .C (clk), .D (new_AGEMA_signal_12135), .Q (new_AGEMA_signal_12136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4315 ( .C (clk), .D (new_AGEMA_signal_12139), .Q (new_AGEMA_signal_12140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4319 ( .C (clk), .D (new_AGEMA_signal_12143), .Q (new_AGEMA_signal_12144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4323 ( .C (clk), .D (new_AGEMA_signal_12147), .Q (new_AGEMA_signal_12148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4327 ( .C (clk), .D (new_AGEMA_signal_12151), .Q (new_AGEMA_signal_12152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4331 ( .C (clk), .D (new_AGEMA_signal_12155), .Q (new_AGEMA_signal_12156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4335 ( .C (clk), .D (new_AGEMA_signal_12159), .Q (new_AGEMA_signal_12160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4339 ( .C (clk), .D (new_AGEMA_signal_12163), .Q (new_AGEMA_signal_12164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4343 ( .C (clk), .D (new_AGEMA_signal_12167), .Q (new_AGEMA_signal_12168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4347 ( .C (clk), .D (new_AGEMA_signal_12171), .Q (new_AGEMA_signal_12172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4351 ( .C (clk), .D (new_AGEMA_signal_12175), .Q (new_AGEMA_signal_12176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4355 ( .C (clk), .D (new_AGEMA_signal_12179), .Q (new_AGEMA_signal_12180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4359 ( .C (clk), .D (new_AGEMA_signal_12183), .Q (new_AGEMA_signal_12184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4363 ( .C (clk), .D (new_AGEMA_signal_12187), .Q (new_AGEMA_signal_12188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4367 ( .C (clk), .D (new_AGEMA_signal_12191), .Q (new_AGEMA_signal_12192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4371 ( .C (clk), .D (new_AGEMA_signal_12195), .Q (new_AGEMA_signal_12196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4375 ( .C (clk), .D (new_AGEMA_signal_12199), .Q (new_AGEMA_signal_12200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4379 ( .C (clk), .D (new_AGEMA_signal_12203), .Q (new_AGEMA_signal_12204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4383 ( .C (clk), .D (new_AGEMA_signal_12207), .Q (new_AGEMA_signal_12208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4387 ( .C (clk), .D (new_AGEMA_signal_12211), .Q (new_AGEMA_signal_12212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4391 ( .C (clk), .D (new_AGEMA_signal_12215), .Q (new_AGEMA_signal_12216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4395 ( .C (clk), .D (new_AGEMA_signal_12219), .Q (new_AGEMA_signal_12220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4399 ( .C (clk), .D (new_AGEMA_signal_12223), .Q (new_AGEMA_signal_12224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4403 ( .C (clk), .D (new_AGEMA_signal_12227), .Q (new_AGEMA_signal_12228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4407 ( .C (clk), .D (new_AGEMA_signal_12231), .Q (new_AGEMA_signal_12232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4411 ( .C (clk), .D (new_AGEMA_signal_12235), .Q (new_AGEMA_signal_12236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4415 ( .C (clk), .D (new_AGEMA_signal_12239), .Q (new_AGEMA_signal_12240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4419 ( .C (clk), .D (new_AGEMA_signal_12243), .Q (new_AGEMA_signal_12244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4423 ( .C (clk), .D (new_AGEMA_signal_12247), .Q (new_AGEMA_signal_12248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4427 ( .C (clk), .D (new_AGEMA_signal_12251), .Q (new_AGEMA_signal_12252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4431 ( .C (clk), .D (new_AGEMA_signal_12255), .Q (new_AGEMA_signal_12256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4435 ( .C (clk), .D (new_AGEMA_signal_12259), .Q (new_AGEMA_signal_12260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4439 ( .C (clk), .D (new_AGEMA_signal_12263), .Q (new_AGEMA_signal_12264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4443 ( .C (clk), .D (new_AGEMA_signal_12267), .Q (new_AGEMA_signal_12268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4447 ( .C (clk), .D (new_AGEMA_signal_12271), .Q (new_AGEMA_signal_12272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4451 ( .C (clk), .D (new_AGEMA_signal_12275), .Q (new_AGEMA_signal_12276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4455 ( .C (clk), .D (new_AGEMA_signal_12279), .Q (new_AGEMA_signal_12280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4459 ( .C (clk), .D (new_AGEMA_signal_12283), .Q (new_AGEMA_signal_12284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4463 ( .C (clk), .D (new_AGEMA_signal_12287), .Q (new_AGEMA_signal_12288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4467 ( .C (clk), .D (new_AGEMA_signal_12291), .Q (new_AGEMA_signal_12292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4471 ( .C (clk), .D (new_AGEMA_signal_12295), .Q (new_AGEMA_signal_12296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4475 ( .C (clk), .D (new_AGEMA_signal_12299), .Q (new_AGEMA_signal_12300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4479 ( .C (clk), .D (new_AGEMA_signal_12303), .Q (new_AGEMA_signal_12304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4483 ( .C (clk), .D (new_AGEMA_signal_12307), .Q (new_AGEMA_signal_12308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4487 ( .C (clk), .D (new_AGEMA_signal_12311), .Q (new_AGEMA_signal_12312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4491 ( .C (clk), .D (new_AGEMA_signal_12315), .Q (new_AGEMA_signal_12316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4495 ( .C (clk), .D (new_AGEMA_signal_12319), .Q (new_AGEMA_signal_12320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4499 ( .C (clk), .D (new_AGEMA_signal_12323), .Q (new_AGEMA_signal_12324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4503 ( .C (clk), .D (new_AGEMA_signal_12327), .Q (new_AGEMA_signal_12328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4507 ( .C (clk), .D (new_AGEMA_signal_12331), .Q (new_AGEMA_signal_12332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4511 ( .C (clk), .D (new_AGEMA_signal_12335), .Q (new_AGEMA_signal_12336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4515 ( .C (clk), .D (new_AGEMA_signal_12339), .Q (new_AGEMA_signal_12340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4519 ( .C (clk), .D (new_AGEMA_signal_12343), .Q (new_AGEMA_signal_12344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4523 ( .C (clk), .D (new_AGEMA_signal_12347), .Q (new_AGEMA_signal_12348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4527 ( .C (clk), .D (new_AGEMA_signal_12351), .Q (new_AGEMA_signal_12352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4531 ( .C (clk), .D (new_AGEMA_signal_12355), .Q (new_AGEMA_signal_12356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4535 ( .C (clk), .D (new_AGEMA_signal_12359), .Q (new_AGEMA_signal_12360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4539 ( .C (clk), .D (new_AGEMA_signal_12363), .Q (new_AGEMA_signal_12364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4543 ( .C (clk), .D (new_AGEMA_signal_12367), .Q (new_AGEMA_signal_12368) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4547 ( .C (clk), .D (new_AGEMA_signal_12371), .Q (new_AGEMA_signal_12372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4551 ( .C (clk), .D (new_AGEMA_signal_12375), .Q (new_AGEMA_signal_12376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4555 ( .C (clk), .D (new_AGEMA_signal_12379), .Q (new_AGEMA_signal_12380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4559 ( .C (clk), .D (new_AGEMA_signal_12383), .Q (new_AGEMA_signal_12384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4563 ( .C (clk), .D (new_AGEMA_signal_12387), .Q (new_AGEMA_signal_12388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4567 ( .C (clk), .D (new_AGEMA_signal_12391), .Q (new_AGEMA_signal_12392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4571 ( .C (clk), .D (new_AGEMA_signal_12395), .Q (new_AGEMA_signal_12396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4575 ( .C (clk), .D (new_AGEMA_signal_12399), .Q (new_AGEMA_signal_12400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4579 ( .C (clk), .D (new_AGEMA_signal_12403), .Q (new_AGEMA_signal_12404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4583 ( .C (clk), .D (new_AGEMA_signal_12407), .Q (new_AGEMA_signal_12408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4587 ( .C (clk), .D (new_AGEMA_signal_12411), .Q (new_AGEMA_signal_12412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4591 ( .C (clk), .D (new_AGEMA_signal_12415), .Q (new_AGEMA_signal_12416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4595 ( .C (clk), .D (new_AGEMA_signal_12419), .Q (new_AGEMA_signal_12420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4599 ( .C (clk), .D (new_AGEMA_signal_12423), .Q (new_AGEMA_signal_12424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4603 ( .C (clk), .D (new_AGEMA_signal_12427), .Q (new_AGEMA_signal_12428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4607 ( .C (clk), .D (new_AGEMA_signal_12431), .Q (new_AGEMA_signal_12432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4611 ( .C (clk), .D (new_AGEMA_signal_12435), .Q (new_AGEMA_signal_12436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4615 ( .C (clk), .D (new_AGEMA_signal_12439), .Q (new_AGEMA_signal_12440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4619 ( .C (clk), .D (new_AGEMA_signal_12443), .Q (new_AGEMA_signal_12444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4623 ( .C (clk), .D (new_AGEMA_signal_12447), .Q (new_AGEMA_signal_12448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4627 ( .C (clk), .D (new_AGEMA_signal_12451), .Q (new_AGEMA_signal_12452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4631 ( .C (clk), .D (new_AGEMA_signal_12455), .Q (new_AGEMA_signal_12456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4635 ( .C (clk), .D (new_AGEMA_signal_12459), .Q (new_AGEMA_signal_12460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4639 ( .C (clk), .D (new_AGEMA_signal_12463), .Q (new_AGEMA_signal_12464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4643 ( .C (clk), .D (new_AGEMA_signal_12467), .Q (new_AGEMA_signal_12468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4647 ( .C (clk), .D (new_AGEMA_signal_12471), .Q (new_AGEMA_signal_12472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4651 ( .C (clk), .D (new_AGEMA_signal_12475), .Q (new_AGEMA_signal_12476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4655 ( .C (clk), .D (new_AGEMA_signal_12479), .Q (new_AGEMA_signal_12480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4659 ( .C (clk), .D (new_AGEMA_signal_12483), .Q (new_AGEMA_signal_12484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4663 ( .C (clk), .D (new_AGEMA_signal_12487), .Q (new_AGEMA_signal_12488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4667 ( .C (clk), .D (new_AGEMA_signal_12491), .Q (new_AGEMA_signal_12492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4671 ( .C (clk), .D (new_AGEMA_signal_12495), .Q (new_AGEMA_signal_12496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4675 ( .C (clk), .D (new_AGEMA_signal_12499), .Q (new_AGEMA_signal_12500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4679 ( .C (clk), .D (new_AGEMA_signal_12503), .Q (new_AGEMA_signal_12504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4683 ( .C (clk), .D (new_AGEMA_signal_12507), .Q (new_AGEMA_signal_12508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4687 ( .C (clk), .D (new_AGEMA_signal_12511), .Q (new_AGEMA_signal_12512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4691 ( .C (clk), .D (new_AGEMA_signal_12515), .Q (new_AGEMA_signal_12516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4695 ( .C (clk), .D (new_AGEMA_signal_12519), .Q (new_AGEMA_signal_12520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4699 ( .C (clk), .D (new_AGEMA_signal_12523), .Q (new_AGEMA_signal_12524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4703 ( .C (clk), .D (new_AGEMA_signal_12527), .Q (new_AGEMA_signal_12528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4707 ( .C (clk), .D (new_AGEMA_signal_12531), .Q (new_AGEMA_signal_12532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4711 ( .C (clk), .D (new_AGEMA_signal_12535), .Q (new_AGEMA_signal_12536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4715 ( .C (clk), .D (new_AGEMA_signal_12539), .Q (new_AGEMA_signal_12540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4719 ( .C (clk), .D (new_AGEMA_signal_12543), .Q (new_AGEMA_signal_12544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4723 ( .C (clk), .D (new_AGEMA_signal_12547), .Q (new_AGEMA_signal_12548) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4727 ( .C (clk), .D (new_AGEMA_signal_12551), .Q (new_AGEMA_signal_12552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4731 ( .C (clk), .D (new_AGEMA_signal_12555), .Q (new_AGEMA_signal_12556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4735 ( .C (clk), .D (new_AGEMA_signal_12559), .Q (new_AGEMA_signal_12560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4739 ( .C (clk), .D (new_AGEMA_signal_12563), .Q (new_AGEMA_signal_12564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4743 ( .C (clk), .D (new_AGEMA_signal_12567), .Q (new_AGEMA_signal_12568) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4747 ( .C (clk), .D (new_AGEMA_signal_12571), .Q (new_AGEMA_signal_12572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4751 ( .C (clk), .D (new_AGEMA_signal_12575), .Q (new_AGEMA_signal_12576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4755 ( .C (clk), .D (new_AGEMA_signal_12579), .Q (new_AGEMA_signal_12580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4759 ( .C (clk), .D (new_AGEMA_signal_12583), .Q (new_AGEMA_signal_12584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4763 ( .C (clk), .D (new_AGEMA_signal_12587), .Q (new_AGEMA_signal_12588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4767 ( .C (clk), .D (new_AGEMA_signal_12591), .Q (new_AGEMA_signal_12592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4771 ( .C (clk), .D (new_AGEMA_signal_12595), .Q (new_AGEMA_signal_12596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4775 ( .C (clk), .D (new_AGEMA_signal_12599), .Q (new_AGEMA_signal_12600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4779 ( .C (clk), .D (new_AGEMA_signal_12603), .Q (new_AGEMA_signal_12604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4783 ( .C (clk), .D (new_AGEMA_signal_12607), .Q (new_AGEMA_signal_12608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4787 ( .C (clk), .D (new_AGEMA_signal_12611), .Q (new_AGEMA_signal_12612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4791 ( .C (clk), .D (new_AGEMA_signal_12615), .Q (new_AGEMA_signal_12616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4795 ( .C (clk), .D (new_AGEMA_signal_12619), .Q (new_AGEMA_signal_12620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4799 ( .C (clk), .D (new_AGEMA_signal_12623), .Q (new_AGEMA_signal_12624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4803 ( .C (clk), .D (new_AGEMA_signal_12627), .Q (new_AGEMA_signal_12628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4807 ( .C (clk), .D (new_AGEMA_signal_12631), .Q (new_AGEMA_signal_12632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4811 ( .C (clk), .D (new_AGEMA_signal_12635), .Q (new_AGEMA_signal_12636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4815 ( .C (clk), .D (new_AGEMA_signal_12639), .Q (new_AGEMA_signal_12640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4819 ( .C (clk), .D (new_AGEMA_signal_12643), .Q (new_AGEMA_signal_12644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4823 ( .C (clk), .D (new_AGEMA_signal_12647), .Q (new_AGEMA_signal_12648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4827 ( .C (clk), .D (new_AGEMA_signal_12651), .Q (new_AGEMA_signal_12652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4831 ( .C (clk), .D (new_AGEMA_signal_12655), .Q (new_AGEMA_signal_12656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4835 ( .C (clk), .D (new_AGEMA_signal_12659), .Q (new_AGEMA_signal_12660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4839 ( .C (clk), .D (new_AGEMA_signal_12663), .Q (new_AGEMA_signal_12664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4843 ( .C (clk), .D (new_AGEMA_signal_12667), .Q (new_AGEMA_signal_12668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4847 ( .C (clk), .D (new_AGEMA_signal_12671), .Q (new_AGEMA_signal_12672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4851 ( .C (clk), .D (new_AGEMA_signal_12675), .Q (new_AGEMA_signal_12676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4855 ( .C (clk), .D (new_AGEMA_signal_12679), .Q (new_AGEMA_signal_12680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4859 ( .C (clk), .D (new_AGEMA_signal_12683), .Q (new_AGEMA_signal_12684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4863 ( .C (clk), .D (new_AGEMA_signal_12687), .Q (new_AGEMA_signal_12688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4867 ( .C (clk), .D (new_AGEMA_signal_12691), .Q (new_AGEMA_signal_12692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4871 ( .C (clk), .D (new_AGEMA_signal_12695), .Q (new_AGEMA_signal_12696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4875 ( .C (clk), .D (new_AGEMA_signal_12699), .Q (new_AGEMA_signal_12700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4879 ( .C (clk), .D (new_AGEMA_signal_12703), .Q (new_AGEMA_signal_12704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4883 ( .C (clk), .D (new_AGEMA_signal_12707), .Q (new_AGEMA_signal_12708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4887 ( .C (clk), .D (new_AGEMA_signal_12711), .Q (new_AGEMA_signal_12712) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4891 ( .C (clk), .D (new_AGEMA_signal_12715), .Q (new_AGEMA_signal_12716) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4895 ( .C (clk), .D (new_AGEMA_signal_12719), .Q (new_AGEMA_signal_12720) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4899 ( .C (clk), .D (new_AGEMA_signal_12723), .Q (new_AGEMA_signal_12724) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4903 ( .C (clk), .D (new_AGEMA_signal_12727), .Q (new_AGEMA_signal_12728) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4907 ( .C (clk), .D (new_AGEMA_signal_12731), .Q (new_AGEMA_signal_12732) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4911 ( .C (clk), .D (new_AGEMA_signal_12735), .Q (new_AGEMA_signal_12736) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4915 ( .C (clk), .D (new_AGEMA_signal_12739), .Q (new_AGEMA_signal_12740) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4919 ( .C (clk), .D (new_AGEMA_signal_12743), .Q (new_AGEMA_signal_12744) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4923 ( .C (clk), .D (new_AGEMA_signal_12747), .Q (new_AGEMA_signal_12748) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4927 ( .C (clk), .D (new_AGEMA_signal_12751), .Q (new_AGEMA_signal_12752) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4931 ( .C (clk), .D (new_AGEMA_signal_12755), .Q (new_AGEMA_signal_12756) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4935 ( .C (clk), .D (new_AGEMA_signal_12759), .Q (new_AGEMA_signal_12760) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4939 ( .C (clk), .D (new_AGEMA_signal_12763), .Q (new_AGEMA_signal_12764) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4943 ( .C (clk), .D (new_AGEMA_signal_12767), .Q (new_AGEMA_signal_12768) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4947 ( .C (clk), .D (new_AGEMA_signal_12771), .Q (new_AGEMA_signal_12772) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4951 ( .C (clk), .D (new_AGEMA_signal_12775), .Q (new_AGEMA_signal_12776) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4955 ( .C (clk), .D (new_AGEMA_signal_12779), .Q (new_AGEMA_signal_12780) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4959 ( .C (clk), .D (new_AGEMA_signal_12783), .Q (new_AGEMA_signal_12784) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4963 ( .C (clk), .D (new_AGEMA_signal_12787), .Q (new_AGEMA_signal_12788) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4967 ( .C (clk), .D (new_AGEMA_signal_12791), .Q (new_AGEMA_signal_12792) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4971 ( .C (clk), .D (new_AGEMA_signal_12795), .Q (new_AGEMA_signal_12796) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4975 ( .C (clk), .D (new_AGEMA_signal_12799), .Q (new_AGEMA_signal_12800) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4979 ( .C (clk), .D (new_AGEMA_signal_12803), .Q (new_AGEMA_signal_12804) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4983 ( .C (clk), .D (new_AGEMA_signal_12807), .Q (new_AGEMA_signal_12808) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4987 ( .C (clk), .D (new_AGEMA_signal_12811), .Q (new_AGEMA_signal_12812) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4991 ( .C (clk), .D (new_AGEMA_signal_12815), .Q (new_AGEMA_signal_12816) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4995 ( .C (clk), .D (new_AGEMA_signal_12819), .Q (new_AGEMA_signal_12820) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4999 ( .C (clk), .D (new_AGEMA_signal_12823), .Q (new_AGEMA_signal_12824) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5003 ( .C (clk), .D (new_AGEMA_signal_12827), .Q (new_AGEMA_signal_12828) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5007 ( .C (clk), .D (new_AGEMA_signal_12831), .Q (new_AGEMA_signal_12832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5011 ( .C (clk), .D (new_AGEMA_signal_12835), .Q (new_AGEMA_signal_12836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5015 ( .C (clk), .D (new_AGEMA_signal_12839), .Q (new_AGEMA_signal_12840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5019 ( .C (clk), .D (new_AGEMA_signal_12843), .Q (new_AGEMA_signal_12844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5023 ( .C (clk), .D (new_AGEMA_signal_12847), .Q (new_AGEMA_signal_12848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5027 ( .C (clk), .D (new_AGEMA_signal_12851), .Q (new_AGEMA_signal_12852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5031 ( .C (clk), .D (new_AGEMA_signal_12855), .Q (new_AGEMA_signal_12856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5035 ( .C (clk), .D (new_AGEMA_signal_12859), .Q (new_AGEMA_signal_12860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5039 ( .C (clk), .D (new_AGEMA_signal_12863), .Q (new_AGEMA_signal_12864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5043 ( .C (clk), .D (new_AGEMA_signal_12867), .Q (new_AGEMA_signal_12868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5047 ( .C (clk), .D (new_AGEMA_signal_12871), .Q (new_AGEMA_signal_12872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5051 ( .C (clk), .D (new_AGEMA_signal_12875), .Q (new_AGEMA_signal_12876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5055 ( .C (clk), .D (new_AGEMA_signal_12879), .Q (new_AGEMA_signal_12880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5059 ( .C (clk), .D (new_AGEMA_signal_12883), .Q (new_AGEMA_signal_12884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5063 ( .C (clk), .D (new_AGEMA_signal_12887), .Q (new_AGEMA_signal_12888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5067 ( .C (clk), .D (new_AGEMA_signal_12891), .Q (new_AGEMA_signal_12892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5071 ( .C (clk), .D (new_AGEMA_signal_12895), .Q (new_AGEMA_signal_12896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5075 ( .C (clk), .D (new_AGEMA_signal_12899), .Q (new_AGEMA_signal_12900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5079 ( .C (clk), .D (new_AGEMA_signal_12903), .Q (new_AGEMA_signal_12904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5083 ( .C (clk), .D (new_AGEMA_signal_12907), .Q (new_AGEMA_signal_12908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5087 ( .C (clk), .D (new_AGEMA_signal_12911), .Q (new_AGEMA_signal_12912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5091 ( .C (clk), .D (new_AGEMA_signal_12915), .Q (new_AGEMA_signal_12916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5095 ( .C (clk), .D (new_AGEMA_signal_12919), .Q (new_AGEMA_signal_12920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5099 ( .C (clk), .D (new_AGEMA_signal_12923), .Q (new_AGEMA_signal_12924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5103 ( .C (clk), .D (new_AGEMA_signal_12927), .Q (new_AGEMA_signal_12928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5107 ( .C (clk), .D (new_AGEMA_signal_12931), .Q (new_AGEMA_signal_12932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5111 ( .C (clk), .D (new_AGEMA_signal_12935), .Q (new_AGEMA_signal_12936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5115 ( .C (clk), .D (new_AGEMA_signal_12939), .Q (new_AGEMA_signal_12940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5119 ( .C (clk), .D (new_AGEMA_signal_12943), .Q (new_AGEMA_signal_12944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5123 ( .C (clk), .D (new_AGEMA_signal_12947), .Q (new_AGEMA_signal_12948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5127 ( .C (clk), .D (new_AGEMA_signal_12951), .Q (new_AGEMA_signal_12952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5131 ( .C (clk), .D (new_AGEMA_signal_12955), .Q (new_AGEMA_signal_12956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5135 ( .C (clk), .D (new_AGEMA_signal_12959), .Q (new_AGEMA_signal_12960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5139 ( .C (clk), .D (new_AGEMA_signal_12963), .Q (new_AGEMA_signal_12964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5143 ( .C (clk), .D (new_AGEMA_signal_12967), .Q (new_AGEMA_signal_12968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5147 ( .C (clk), .D (new_AGEMA_signal_12971), .Q (new_AGEMA_signal_12972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5151 ( .C (clk), .D (new_AGEMA_signal_12975), .Q (new_AGEMA_signal_12976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5155 ( .C (clk), .D (new_AGEMA_signal_12979), .Q (new_AGEMA_signal_12980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5159 ( .C (clk), .D (new_AGEMA_signal_12983), .Q (new_AGEMA_signal_12984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5163 ( .C (clk), .D (new_AGEMA_signal_12987), .Q (new_AGEMA_signal_12988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5167 ( .C (clk), .D (new_AGEMA_signal_12991), .Q (new_AGEMA_signal_12992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5171 ( .C (clk), .D (new_AGEMA_signal_12995), .Q (new_AGEMA_signal_12996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5175 ( .C (clk), .D (new_AGEMA_signal_12999), .Q (new_AGEMA_signal_13000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5179 ( .C (clk), .D (new_AGEMA_signal_13003), .Q (new_AGEMA_signal_13004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5183 ( .C (clk), .D (new_AGEMA_signal_13007), .Q (new_AGEMA_signal_13008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5187 ( .C (clk), .D (new_AGEMA_signal_13011), .Q (new_AGEMA_signal_13012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5191 ( .C (clk), .D (new_AGEMA_signal_13015), .Q (new_AGEMA_signal_13016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5195 ( .C (clk), .D (new_AGEMA_signal_13019), .Q (new_AGEMA_signal_13020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5199 ( .C (clk), .D (new_AGEMA_signal_13023), .Q (new_AGEMA_signal_13024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5203 ( .C (clk), .D (new_AGEMA_signal_13027), .Q (new_AGEMA_signal_13028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5207 ( .C (clk), .D (new_AGEMA_signal_13031), .Q (new_AGEMA_signal_13032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5211 ( .C (clk), .D (new_AGEMA_signal_13035), .Q (new_AGEMA_signal_13036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5215 ( .C (clk), .D (new_AGEMA_signal_13039), .Q (new_AGEMA_signal_13040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5219 ( .C (clk), .D (new_AGEMA_signal_13043), .Q (new_AGEMA_signal_13044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5223 ( .C (clk), .D (new_AGEMA_signal_13047), .Q (new_AGEMA_signal_13048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5227 ( .C (clk), .D (new_AGEMA_signal_13051), .Q (new_AGEMA_signal_13052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5231 ( .C (clk), .D (new_AGEMA_signal_13055), .Q (new_AGEMA_signal_13056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5235 ( .C (clk), .D (new_AGEMA_signal_13059), .Q (new_AGEMA_signal_13060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5239 ( .C (clk), .D (new_AGEMA_signal_13063), .Q (new_AGEMA_signal_13064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5243 ( .C (clk), .D (new_AGEMA_signal_13067), .Q (new_AGEMA_signal_13068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5247 ( .C (clk), .D (new_AGEMA_signal_13071), .Q (new_AGEMA_signal_13072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5251 ( .C (clk), .D (new_AGEMA_signal_13075), .Q (new_AGEMA_signal_13076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5255 ( .C (clk), .D (new_AGEMA_signal_13079), .Q (new_AGEMA_signal_13080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5259 ( .C (clk), .D (new_AGEMA_signal_13083), .Q (new_AGEMA_signal_13084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5263 ( .C (clk), .D (new_AGEMA_signal_13087), .Q (new_AGEMA_signal_13088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5267 ( .C (clk), .D (new_AGEMA_signal_13091), .Q (new_AGEMA_signal_13092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5271 ( .C (clk), .D (new_AGEMA_signal_13095), .Q (new_AGEMA_signal_13096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5275 ( .C (clk), .D (new_AGEMA_signal_13099), .Q (new_AGEMA_signal_13100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5279 ( .C (clk), .D (new_AGEMA_signal_13103), .Q (new_AGEMA_signal_13104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5283 ( .C (clk), .D (new_AGEMA_signal_13107), .Q (new_AGEMA_signal_13108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5287 ( .C (clk), .D (new_AGEMA_signal_13111), .Q (new_AGEMA_signal_13112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5291 ( .C (clk), .D (new_AGEMA_signal_13115), .Q (new_AGEMA_signal_13116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5295 ( .C (clk), .D (new_AGEMA_signal_13119), .Q (new_AGEMA_signal_13120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5299 ( .C (clk), .D (new_AGEMA_signal_13123), .Q (new_AGEMA_signal_13124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5303 ( .C (clk), .D (new_AGEMA_signal_13127), .Q (new_AGEMA_signal_13128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5307 ( .C (clk), .D (new_AGEMA_signal_13131), .Q (new_AGEMA_signal_13132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5311 ( .C (clk), .D (new_AGEMA_signal_13135), .Q (new_AGEMA_signal_13136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5315 ( .C (clk), .D (new_AGEMA_signal_13139), .Q (new_AGEMA_signal_13140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5319 ( .C (clk), .D (new_AGEMA_signal_13143), .Q (new_AGEMA_signal_13144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5323 ( .C (clk), .D (new_AGEMA_signal_13147), .Q (new_AGEMA_signal_13148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5327 ( .C (clk), .D (new_AGEMA_signal_13151), .Q (new_AGEMA_signal_13152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5331 ( .C (clk), .D (new_AGEMA_signal_13155), .Q (new_AGEMA_signal_13156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5335 ( .C (clk), .D (new_AGEMA_signal_13159), .Q (new_AGEMA_signal_13160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5339 ( .C (clk), .D (new_AGEMA_signal_13163), .Q (new_AGEMA_signal_13164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5343 ( .C (clk), .D (new_AGEMA_signal_13167), .Q (new_AGEMA_signal_13168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5347 ( .C (clk), .D (new_AGEMA_signal_13171), .Q (new_AGEMA_signal_13172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5351 ( .C (clk), .D (new_AGEMA_signal_13175), .Q (new_AGEMA_signal_13176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5355 ( .C (clk), .D (new_AGEMA_signal_13179), .Q (new_AGEMA_signal_13180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5359 ( .C (clk), .D (new_AGEMA_signal_13183), .Q (new_AGEMA_signal_13184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5363 ( .C (clk), .D (new_AGEMA_signal_13187), .Q (new_AGEMA_signal_13188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5367 ( .C (clk), .D (new_AGEMA_signal_13191), .Q (new_AGEMA_signal_13192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5371 ( .C (clk), .D (new_AGEMA_signal_13195), .Q (new_AGEMA_signal_13196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5375 ( .C (clk), .D (new_AGEMA_signal_13199), .Q (new_AGEMA_signal_13200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5379 ( .C (clk), .D (new_AGEMA_signal_13203), .Q (new_AGEMA_signal_13204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5383 ( .C (clk), .D (new_AGEMA_signal_13207), .Q (new_AGEMA_signal_13208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5387 ( .C (clk), .D (new_AGEMA_signal_13211), .Q (new_AGEMA_signal_13212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5391 ( .C (clk), .D (new_AGEMA_signal_13215), .Q (new_AGEMA_signal_13216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5395 ( .C (clk), .D (new_AGEMA_signal_13219), .Q (new_AGEMA_signal_13220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5399 ( .C (clk), .D (new_AGEMA_signal_13223), .Q (new_AGEMA_signal_13224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5403 ( .C (clk), .D (new_AGEMA_signal_13227), .Q (new_AGEMA_signal_13228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5407 ( .C (clk), .D (new_AGEMA_signal_13231), .Q (new_AGEMA_signal_13232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5411 ( .C (clk), .D (new_AGEMA_signal_13235), .Q (new_AGEMA_signal_13236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5415 ( .C (clk), .D (new_AGEMA_signal_13239), .Q (new_AGEMA_signal_13240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5419 ( .C (clk), .D (new_AGEMA_signal_13243), .Q (new_AGEMA_signal_13244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5423 ( .C (clk), .D (new_AGEMA_signal_13247), .Q (new_AGEMA_signal_13248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5427 ( .C (clk), .D (new_AGEMA_signal_13251), .Q (new_AGEMA_signal_13252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5431 ( .C (clk), .D (new_AGEMA_signal_13255), .Q (new_AGEMA_signal_13256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5435 ( .C (clk), .D (new_AGEMA_signal_13259), .Q (new_AGEMA_signal_13260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5439 ( .C (clk), .D (new_AGEMA_signal_13263), .Q (new_AGEMA_signal_13264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5443 ( .C (clk), .D (new_AGEMA_signal_13267), .Q (new_AGEMA_signal_13268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5447 ( .C (clk), .D (new_AGEMA_signal_13271), .Q (new_AGEMA_signal_13272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5451 ( .C (clk), .D (new_AGEMA_signal_13275), .Q (new_AGEMA_signal_13276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5455 ( .C (clk), .D (new_AGEMA_signal_13279), .Q (new_AGEMA_signal_13280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5459 ( .C (clk), .D (new_AGEMA_signal_13283), .Q (new_AGEMA_signal_13284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5463 ( .C (clk), .D (new_AGEMA_signal_13287), .Q (new_AGEMA_signal_13288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5467 ( .C (clk), .D (new_AGEMA_signal_13291), .Q (new_AGEMA_signal_13292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5471 ( .C (clk), .D (new_AGEMA_signal_13295), .Q (new_AGEMA_signal_13296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5475 ( .C (clk), .D (new_AGEMA_signal_13299), .Q (new_AGEMA_signal_13300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5479 ( .C (clk), .D (new_AGEMA_signal_13303), .Q (new_AGEMA_signal_13304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5483 ( .C (clk), .D (new_AGEMA_signal_13307), .Q (new_AGEMA_signal_13308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5487 ( .C (clk), .D (new_AGEMA_signal_13311), .Q (new_AGEMA_signal_13312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5491 ( .C (clk), .D (new_AGEMA_signal_13315), .Q (new_AGEMA_signal_13316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5495 ( .C (clk), .D (new_AGEMA_signal_13319), .Q (new_AGEMA_signal_13320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5499 ( .C (clk), .D (new_AGEMA_signal_13323), .Q (new_AGEMA_signal_13324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5503 ( .C (clk), .D (new_AGEMA_signal_13327), .Q (new_AGEMA_signal_13328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5507 ( .C (clk), .D (new_AGEMA_signal_13331), .Q (new_AGEMA_signal_13332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5511 ( .C (clk), .D (new_AGEMA_signal_13335), .Q (new_AGEMA_signal_13336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5515 ( .C (clk), .D (new_AGEMA_signal_13339), .Q (new_AGEMA_signal_13340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5519 ( .C (clk), .D (new_AGEMA_signal_13343), .Q (new_AGEMA_signal_13344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5523 ( .C (clk), .D (new_AGEMA_signal_13347), .Q (new_AGEMA_signal_13348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5527 ( .C (clk), .D (new_AGEMA_signal_13351), .Q (new_AGEMA_signal_13352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5531 ( .C (clk), .D (new_AGEMA_signal_13355), .Q (new_AGEMA_signal_13356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5535 ( .C (clk), .D (new_AGEMA_signal_13359), .Q (new_AGEMA_signal_13360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5539 ( .C (clk), .D (new_AGEMA_signal_13363), .Q (new_AGEMA_signal_13364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5543 ( .C (clk), .D (new_AGEMA_signal_13367), .Q (new_AGEMA_signal_13368) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5547 ( .C (clk), .D (new_AGEMA_signal_13371), .Q (new_AGEMA_signal_13372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5551 ( .C (clk), .D (new_AGEMA_signal_13375), .Q (new_AGEMA_signal_13376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5555 ( .C (clk), .D (new_AGEMA_signal_13379), .Q (new_AGEMA_signal_13380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5559 ( .C (clk), .D (new_AGEMA_signal_13383), .Q (new_AGEMA_signal_13384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5563 ( .C (clk), .D (new_AGEMA_signal_13387), .Q (new_AGEMA_signal_13388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5567 ( .C (clk), .D (new_AGEMA_signal_13391), .Q (new_AGEMA_signal_13392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5571 ( .C (clk), .D (new_AGEMA_signal_13395), .Q (new_AGEMA_signal_13396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5575 ( .C (clk), .D (new_AGEMA_signal_13399), .Q (new_AGEMA_signal_13400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5579 ( .C (clk), .D (new_AGEMA_signal_13403), .Q (new_AGEMA_signal_13404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5583 ( .C (clk), .D (new_AGEMA_signal_13407), .Q (new_AGEMA_signal_13408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5587 ( .C (clk), .D (new_AGEMA_signal_13411), .Q (new_AGEMA_signal_13412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5591 ( .C (clk), .D (new_AGEMA_signal_13415), .Q (new_AGEMA_signal_13416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5595 ( .C (clk), .D (new_AGEMA_signal_13419), .Q (new_AGEMA_signal_13420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5599 ( .C (clk), .D (new_AGEMA_signal_13423), .Q (new_AGEMA_signal_13424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5603 ( .C (clk), .D (new_AGEMA_signal_13427), .Q (new_AGEMA_signal_13428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5607 ( .C (clk), .D (new_AGEMA_signal_13431), .Q (new_AGEMA_signal_13432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5611 ( .C (clk), .D (new_AGEMA_signal_13435), .Q (new_AGEMA_signal_13436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5615 ( .C (clk), .D (new_AGEMA_signal_13439), .Q (new_AGEMA_signal_13440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5619 ( .C (clk), .D (new_AGEMA_signal_13443), .Q (new_AGEMA_signal_13444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5623 ( .C (clk), .D (new_AGEMA_signal_13447), .Q (new_AGEMA_signal_13448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5627 ( .C (clk), .D (new_AGEMA_signal_13451), .Q (new_AGEMA_signal_13452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5631 ( .C (clk), .D (new_AGEMA_signal_13455), .Q (new_AGEMA_signal_13456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5635 ( .C (clk), .D (new_AGEMA_signal_13459), .Q (new_AGEMA_signal_13460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5639 ( .C (clk), .D (new_AGEMA_signal_13463), .Q (new_AGEMA_signal_13464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5643 ( .C (clk), .D (new_AGEMA_signal_13467), .Q (new_AGEMA_signal_13468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5647 ( .C (clk), .D (new_AGEMA_signal_13471), .Q (new_AGEMA_signal_13472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5651 ( .C (clk), .D (new_AGEMA_signal_13475), .Q (new_AGEMA_signal_13476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5655 ( .C (clk), .D (new_AGEMA_signal_13479), .Q (new_AGEMA_signal_13480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5659 ( .C (clk), .D (new_AGEMA_signal_13483), .Q (new_AGEMA_signal_13484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5663 ( .C (clk), .D (new_AGEMA_signal_13487), .Q (new_AGEMA_signal_13488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5667 ( .C (clk), .D (new_AGEMA_signal_13491), .Q (new_AGEMA_signal_13492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5671 ( .C (clk), .D (new_AGEMA_signal_13495), .Q (new_AGEMA_signal_13496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5675 ( .C (clk), .D (new_AGEMA_signal_13499), .Q (new_AGEMA_signal_13500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5679 ( .C (clk), .D (new_AGEMA_signal_13503), .Q (new_AGEMA_signal_13504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5683 ( .C (clk), .D (new_AGEMA_signal_13507), .Q (new_AGEMA_signal_13508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5687 ( .C (clk), .D (new_AGEMA_signal_13511), .Q (new_AGEMA_signal_13512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5691 ( .C (clk), .D (new_AGEMA_signal_13515), .Q (new_AGEMA_signal_13516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5695 ( .C (clk), .D (new_AGEMA_signal_13519), .Q (new_AGEMA_signal_13520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5699 ( .C (clk), .D (new_AGEMA_signal_13523), .Q (new_AGEMA_signal_13524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5703 ( .C (clk), .D (new_AGEMA_signal_13527), .Q (new_AGEMA_signal_13528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5707 ( .C (clk), .D (new_AGEMA_signal_13531), .Q (new_AGEMA_signal_13532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5711 ( .C (clk), .D (new_AGEMA_signal_13535), .Q (new_AGEMA_signal_13536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5715 ( .C (clk), .D (new_AGEMA_signal_13539), .Q (new_AGEMA_signal_13540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5719 ( .C (clk), .D (new_AGEMA_signal_13543), .Q (new_AGEMA_signal_13544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5723 ( .C (clk), .D (new_AGEMA_signal_13547), .Q (new_AGEMA_signal_13548) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5727 ( .C (clk), .D (new_AGEMA_signal_13551), .Q (new_AGEMA_signal_13552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5731 ( .C (clk), .D (new_AGEMA_signal_13555), .Q (new_AGEMA_signal_13556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5735 ( .C (clk), .D (new_AGEMA_signal_13559), .Q (new_AGEMA_signal_13560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5739 ( .C (clk), .D (new_AGEMA_signal_13563), .Q (new_AGEMA_signal_13564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5743 ( .C (clk), .D (new_AGEMA_signal_13567), .Q (new_AGEMA_signal_13568) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5747 ( .C (clk), .D (new_AGEMA_signal_13571), .Q (new_AGEMA_signal_13572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5751 ( .C (clk), .D (new_AGEMA_signal_13575), .Q (new_AGEMA_signal_13576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5755 ( .C (clk), .D (new_AGEMA_signal_13579), .Q (new_AGEMA_signal_13580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5759 ( .C (clk), .D (new_AGEMA_signal_13583), .Q (new_AGEMA_signal_13584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5763 ( .C (clk), .D (new_AGEMA_signal_13587), .Q (new_AGEMA_signal_13588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5767 ( .C (clk), .D (new_AGEMA_signal_13591), .Q (new_AGEMA_signal_13592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5771 ( .C (clk), .D (new_AGEMA_signal_13595), .Q (new_AGEMA_signal_13596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5775 ( .C (clk), .D (new_AGEMA_signal_13599), .Q (new_AGEMA_signal_13600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5779 ( .C (clk), .D (new_AGEMA_signal_13603), .Q (new_AGEMA_signal_13604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5783 ( .C (clk), .D (new_AGEMA_signal_13607), .Q (new_AGEMA_signal_13608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5787 ( .C (clk), .D (new_AGEMA_signal_13611), .Q (new_AGEMA_signal_13612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5791 ( .C (clk), .D (new_AGEMA_signal_13615), .Q (new_AGEMA_signal_13616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5795 ( .C (clk), .D (new_AGEMA_signal_13619), .Q (new_AGEMA_signal_13620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5799 ( .C (clk), .D (new_AGEMA_signal_13623), .Q (new_AGEMA_signal_13624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5803 ( .C (clk), .D (new_AGEMA_signal_13627), .Q (new_AGEMA_signal_13628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5807 ( .C (clk), .D (new_AGEMA_signal_13631), .Q (new_AGEMA_signal_13632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5811 ( .C (clk), .D (new_AGEMA_signal_13635), .Q (new_AGEMA_signal_13636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5815 ( .C (clk), .D (new_AGEMA_signal_13639), .Q (new_AGEMA_signal_13640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5819 ( .C (clk), .D (new_AGEMA_signal_13643), .Q (new_AGEMA_signal_13644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5823 ( .C (clk), .D (new_AGEMA_signal_13647), .Q (new_AGEMA_signal_13648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5827 ( .C (clk), .D (new_AGEMA_signal_13651), .Q (new_AGEMA_signal_13652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5831 ( .C (clk), .D (new_AGEMA_signal_13655), .Q (new_AGEMA_signal_13656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5835 ( .C (clk), .D (new_AGEMA_signal_13659), .Q (new_AGEMA_signal_13660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5839 ( .C (clk), .D (new_AGEMA_signal_13663), .Q (new_AGEMA_signal_13664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5843 ( .C (clk), .D (new_AGEMA_signal_13667), .Q (new_AGEMA_signal_13668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5847 ( .C (clk), .D (new_AGEMA_signal_13671), .Q (new_AGEMA_signal_13672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5851 ( .C (clk), .D (new_AGEMA_signal_13675), .Q (new_AGEMA_signal_13676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5855 ( .C (clk), .D (new_AGEMA_signal_13679), .Q (new_AGEMA_signal_13680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5859 ( .C (clk), .D (new_AGEMA_signal_13683), .Q (new_AGEMA_signal_13684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5863 ( .C (clk), .D (new_AGEMA_signal_13687), .Q (new_AGEMA_signal_13688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5867 ( .C (clk), .D (new_AGEMA_signal_13691), .Q (new_AGEMA_signal_13692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5871 ( .C (clk), .D (new_AGEMA_signal_13695), .Q (new_AGEMA_signal_13696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5875 ( .C (clk), .D (new_AGEMA_signal_13699), .Q (new_AGEMA_signal_13700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5879 ( .C (clk), .D (new_AGEMA_signal_13703), .Q (new_AGEMA_signal_13704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5883 ( .C (clk), .D (new_AGEMA_signal_13707), .Q (new_AGEMA_signal_13708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5887 ( .C (clk), .D (new_AGEMA_signal_13711), .Q (new_AGEMA_signal_13712) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5891 ( .C (clk), .D (new_AGEMA_signal_13715), .Q (new_AGEMA_signal_13716) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5895 ( .C (clk), .D (new_AGEMA_signal_13719), .Q (new_AGEMA_signal_13720) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5899 ( .C (clk), .D (new_AGEMA_signal_13723), .Q (new_AGEMA_signal_13724) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5903 ( .C (clk), .D (new_AGEMA_signal_13727), .Q (new_AGEMA_signal_13728) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5907 ( .C (clk), .D (new_AGEMA_signal_13731), .Q (new_AGEMA_signal_13732) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5911 ( .C (clk), .D (new_AGEMA_signal_13735), .Q (new_AGEMA_signal_13736) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5915 ( .C (clk), .D (new_AGEMA_signal_13739), .Q (new_AGEMA_signal_13740) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5919 ( .C (clk), .D (new_AGEMA_signal_13743), .Q (new_AGEMA_signal_13744) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5923 ( .C (clk), .D (new_AGEMA_signal_13747), .Q (new_AGEMA_signal_13748) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5927 ( .C (clk), .D (new_AGEMA_signal_13751), .Q (new_AGEMA_signal_13752) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5931 ( .C (clk), .D (new_AGEMA_signal_13755), .Q (new_AGEMA_signal_13756) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5935 ( .C (clk), .D (new_AGEMA_signal_13759), .Q (new_AGEMA_signal_13760) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5939 ( .C (clk), .D (new_AGEMA_signal_13763), .Q (new_AGEMA_signal_13764) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5943 ( .C (clk), .D (new_AGEMA_signal_13767), .Q (new_AGEMA_signal_13768) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5947 ( .C (clk), .D (new_AGEMA_signal_13771), .Q (new_AGEMA_signal_13772) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5951 ( .C (clk), .D (new_AGEMA_signal_13775), .Q (new_AGEMA_signal_13776) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5955 ( .C (clk), .D (new_AGEMA_signal_13779), .Q (new_AGEMA_signal_13780) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5959 ( .C (clk), .D (new_AGEMA_signal_13783), .Q (new_AGEMA_signal_13784) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5963 ( .C (clk), .D (new_AGEMA_signal_13787), .Q (new_AGEMA_signal_13788) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5967 ( .C (clk), .D (new_AGEMA_signal_13791), .Q (new_AGEMA_signal_13792) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5971 ( .C (clk), .D (new_AGEMA_signal_13795), .Q (new_AGEMA_signal_13796) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5975 ( .C (clk), .D (new_AGEMA_signal_13799), .Q (new_AGEMA_signal_13800) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5979 ( .C (clk), .D (new_AGEMA_signal_13803), .Q (new_AGEMA_signal_13804) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5983 ( .C (clk), .D (new_AGEMA_signal_13807), .Q (new_AGEMA_signal_13808) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5987 ( .C (clk), .D (new_AGEMA_signal_13811), .Q (new_AGEMA_signal_13812) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5991 ( .C (clk), .D (new_AGEMA_signal_13815), .Q (new_AGEMA_signal_13816) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5995 ( .C (clk), .D (new_AGEMA_signal_13819), .Q (new_AGEMA_signal_13820) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5999 ( .C (clk), .D (new_AGEMA_signal_13823), .Q (new_AGEMA_signal_13824) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6003 ( .C (clk), .D (new_AGEMA_signal_13827), .Q (new_AGEMA_signal_13828) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6007 ( .C (clk), .D (new_AGEMA_signal_13831), .Q (new_AGEMA_signal_13832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6011 ( .C (clk), .D (new_AGEMA_signal_13835), .Q (new_AGEMA_signal_13836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6015 ( .C (clk), .D (new_AGEMA_signal_13839), .Q (new_AGEMA_signal_13840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6019 ( .C (clk), .D (new_AGEMA_signal_13843), .Q (new_AGEMA_signal_13844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6023 ( .C (clk), .D (new_AGEMA_signal_13847), .Q (new_AGEMA_signal_13848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6027 ( .C (clk), .D (new_AGEMA_signal_13851), .Q (new_AGEMA_signal_13852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6031 ( .C (clk), .D (new_AGEMA_signal_13855), .Q (new_AGEMA_signal_13856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6035 ( .C (clk), .D (new_AGEMA_signal_13859), .Q (new_AGEMA_signal_13860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6039 ( .C (clk), .D (new_AGEMA_signal_13863), .Q (new_AGEMA_signal_13864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6043 ( .C (clk), .D (new_AGEMA_signal_13867), .Q (new_AGEMA_signal_13868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6047 ( .C (clk), .D (new_AGEMA_signal_13871), .Q (new_AGEMA_signal_13872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6051 ( .C (clk), .D (new_AGEMA_signal_13875), .Q (new_AGEMA_signal_13876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6055 ( .C (clk), .D (new_AGEMA_signal_13879), .Q (new_AGEMA_signal_13880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6059 ( .C (clk), .D (new_AGEMA_signal_13883), .Q (new_AGEMA_signal_13884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6063 ( .C (clk), .D (new_AGEMA_signal_13887), .Q (new_AGEMA_signal_13888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6067 ( .C (clk), .D (new_AGEMA_signal_13891), .Q (new_AGEMA_signal_13892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6071 ( .C (clk), .D (new_AGEMA_signal_13895), .Q (new_AGEMA_signal_13896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6075 ( .C (clk), .D (new_AGEMA_signal_13899), .Q (new_AGEMA_signal_13900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6079 ( .C (clk), .D (new_AGEMA_signal_13903), .Q (new_AGEMA_signal_13904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6083 ( .C (clk), .D (new_AGEMA_signal_13907), .Q (new_AGEMA_signal_13908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6087 ( .C (clk), .D (new_AGEMA_signal_13911), .Q (new_AGEMA_signal_13912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6091 ( .C (clk), .D (new_AGEMA_signal_13915), .Q (new_AGEMA_signal_13916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6095 ( .C (clk), .D (new_AGEMA_signal_13919), .Q (new_AGEMA_signal_13920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6099 ( .C (clk), .D (new_AGEMA_signal_13923), .Q (new_AGEMA_signal_13924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6103 ( .C (clk), .D (new_AGEMA_signal_13927), .Q (new_AGEMA_signal_13928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6107 ( .C (clk), .D (new_AGEMA_signal_13931), .Q (new_AGEMA_signal_13932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6111 ( .C (clk), .D (new_AGEMA_signal_13935), .Q (new_AGEMA_signal_13936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6115 ( .C (clk), .D (new_AGEMA_signal_13939), .Q (new_AGEMA_signal_13940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6119 ( .C (clk), .D (new_AGEMA_signal_13943), .Q (new_AGEMA_signal_13944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6123 ( .C (clk), .D (new_AGEMA_signal_13947), .Q (new_AGEMA_signal_13948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6127 ( .C (clk), .D (new_AGEMA_signal_13951), .Q (new_AGEMA_signal_13952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6131 ( .C (clk), .D (new_AGEMA_signal_13955), .Q (new_AGEMA_signal_13956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6135 ( .C (clk), .D (new_AGEMA_signal_13959), .Q (new_AGEMA_signal_13960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6139 ( .C (clk), .D (new_AGEMA_signal_13963), .Q (new_AGEMA_signal_13964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6143 ( .C (clk), .D (new_AGEMA_signal_13967), .Q (new_AGEMA_signal_13968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6147 ( .C (clk), .D (new_AGEMA_signal_13971), .Q (new_AGEMA_signal_13972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6151 ( .C (clk), .D (new_AGEMA_signal_13975), .Q (new_AGEMA_signal_13976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6155 ( .C (clk), .D (new_AGEMA_signal_13979), .Q (new_AGEMA_signal_13980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6159 ( .C (clk), .D (new_AGEMA_signal_13983), .Q (new_AGEMA_signal_13984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6163 ( .C (clk), .D (new_AGEMA_signal_13987), .Q (new_AGEMA_signal_13988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6167 ( .C (clk), .D (new_AGEMA_signal_13991), .Q (new_AGEMA_signal_13992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6171 ( .C (clk), .D (new_AGEMA_signal_13995), .Q (new_AGEMA_signal_13996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6175 ( .C (clk), .D (new_AGEMA_signal_13999), .Q (new_AGEMA_signal_14000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6179 ( .C (clk), .D (new_AGEMA_signal_14003), .Q (new_AGEMA_signal_14004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6183 ( .C (clk), .D (new_AGEMA_signal_14007), .Q (new_AGEMA_signal_14008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6187 ( .C (clk), .D (new_AGEMA_signal_14011), .Q (new_AGEMA_signal_14012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6191 ( .C (clk), .D (new_AGEMA_signal_14015), .Q (new_AGEMA_signal_14016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6195 ( .C (clk), .D (new_AGEMA_signal_14019), .Q (new_AGEMA_signal_14020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6199 ( .C (clk), .D (new_AGEMA_signal_14023), .Q (new_AGEMA_signal_14024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6203 ( .C (clk), .D (new_AGEMA_signal_14027), .Q (new_AGEMA_signal_14028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6207 ( .C (clk), .D (new_AGEMA_signal_14031), .Q (new_AGEMA_signal_14032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6211 ( .C (clk), .D (new_AGEMA_signal_14035), .Q (new_AGEMA_signal_14036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6215 ( .C (clk), .D (new_AGEMA_signal_14039), .Q (new_AGEMA_signal_14040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6219 ( .C (clk), .D (new_AGEMA_signal_14043), .Q (new_AGEMA_signal_14044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6223 ( .C (clk), .D (new_AGEMA_signal_14047), .Q (new_AGEMA_signal_14048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6227 ( .C (clk), .D (new_AGEMA_signal_14051), .Q (new_AGEMA_signal_14052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6231 ( .C (clk), .D (new_AGEMA_signal_14055), .Q (new_AGEMA_signal_14056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6235 ( .C (clk), .D (new_AGEMA_signal_14059), .Q (new_AGEMA_signal_14060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6239 ( .C (clk), .D (new_AGEMA_signal_14063), .Q (new_AGEMA_signal_14064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6243 ( .C (clk), .D (new_AGEMA_signal_14067), .Q (new_AGEMA_signal_14068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6247 ( .C (clk), .D (new_AGEMA_signal_14071), .Q (new_AGEMA_signal_14072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6251 ( .C (clk), .D (new_AGEMA_signal_14075), .Q (new_AGEMA_signal_14076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6255 ( .C (clk), .D (new_AGEMA_signal_14079), .Q (new_AGEMA_signal_14080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6259 ( .C (clk), .D (new_AGEMA_signal_14083), .Q (new_AGEMA_signal_14084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6263 ( .C (clk), .D (new_AGEMA_signal_14087), .Q (new_AGEMA_signal_14088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6267 ( .C (clk), .D (new_AGEMA_signal_14091), .Q (new_AGEMA_signal_14092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6271 ( .C (clk), .D (new_AGEMA_signal_14095), .Q (new_AGEMA_signal_14096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6275 ( .C (clk), .D (new_AGEMA_signal_14099), .Q (new_AGEMA_signal_14100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6279 ( .C (clk), .D (new_AGEMA_signal_14103), .Q (new_AGEMA_signal_14104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6283 ( .C (clk), .D (new_AGEMA_signal_14107), .Q (new_AGEMA_signal_14108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6287 ( .C (clk), .D (new_AGEMA_signal_14111), .Q (new_AGEMA_signal_14112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6291 ( .C (clk), .D (new_AGEMA_signal_14115), .Q (new_AGEMA_signal_14116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6295 ( .C (clk), .D (new_AGEMA_signal_14119), .Q (new_AGEMA_signal_14120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6299 ( .C (clk), .D (new_AGEMA_signal_14123), .Q (new_AGEMA_signal_14124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6303 ( .C (clk), .D (new_AGEMA_signal_14127), .Q (new_AGEMA_signal_14128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6307 ( .C (clk), .D (new_AGEMA_signal_14131), .Q (new_AGEMA_signal_14132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6311 ( .C (clk), .D (new_AGEMA_signal_14135), .Q (new_AGEMA_signal_14136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6315 ( .C (clk), .D (new_AGEMA_signal_14139), .Q (new_AGEMA_signal_14140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6319 ( .C (clk), .D (new_AGEMA_signal_14143), .Q (new_AGEMA_signal_14144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6323 ( .C (clk), .D (new_AGEMA_signal_14147), .Q (new_AGEMA_signal_14148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6327 ( .C (clk), .D (new_AGEMA_signal_14151), .Q (new_AGEMA_signal_14152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6331 ( .C (clk), .D (new_AGEMA_signal_14155), .Q (new_AGEMA_signal_14156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6335 ( .C (clk), .D (new_AGEMA_signal_14159), .Q (new_AGEMA_signal_14160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6339 ( .C (clk), .D (new_AGEMA_signal_14163), .Q (new_AGEMA_signal_14164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6343 ( .C (clk), .D (new_AGEMA_signal_14167), .Q (new_AGEMA_signal_14168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6347 ( .C (clk), .D (new_AGEMA_signal_14171), .Q (new_AGEMA_signal_14172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6351 ( .C (clk), .D (new_AGEMA_signal_14175), .Q (new_AGEMA_signal_14176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6355 ( .C (clk), .D (new_AGEMA_signal_14179), .Q (new_AGEMA_signal_14180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6359 ( .C (clk), .D (new_AGEMA_signal_14183), .Q (new_AGEMA_signal_14184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6363 ( .C (clk), .D (new_AGEMA_signal_14187), .Q (new_AGEMA_signal_14188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6367 ( .C (clk), .D (new_AGEMA_signal_14191), .Q (new_AGEMA_signal_14192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6371 ( .C (clk), .D (new_AGEMA_signal_14195), .Q (new_AGEMA_signal_14196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6375 ( .C (clk), .D (new_AGEMA_signal_14199), .Q (new_AGEMA_signal_14200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6379 ( .C (clk), .D (new_AGEMA_signal_14203), .Q (new_AGEMA_signal_14204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6383 ( .C (clk), .D (new_AGEMA_signal_14207), .Q (new_AGEMA_signal_14208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6387 ( .C (clk), .D (new_AGEMA_signal_14211), .Q (new_AGEMA_signal_14212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6391 ( .C (clk), .D (new_AGEMA_signal_14215), .Q (new_AGEMA_signal_14216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6395 ( .C (clk), .D (new_AGEMA_signal_14219), .Q (new_AGEMA_signal_14220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6399 ( .C (clk), .D (new_AGEMA_signal_14223), .Q (new_AGEMA_signal_14224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6403 ( .C (clk), .D (new_AGEMA_signal_14227), .Q (new_AGEMA_signal_14228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6407 ( .C (clk), .D (new_AGEMA_signal_14231), .Q (new_AGEMA_signal_14232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6411 ( .C (clk), .D (new_AGEMA_signal_14235), .Q (new_AGEMA_signal_14236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6415 ( .C (clk), .D (new_AGEMA_signal_14239), .Q (new_AGEMA_signal_14240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6419 ( .C (clk), .D (new_AGEMA_signal_14243), .Q (new_AGEMA_signal_14244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6423 ( .C (clk), .D (new_AGEMA_signal_14247), .Q (new_AGEMA_signal_14248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6427 ( .C (clk), .D (new_AGEMA_signal_14251), .Q (new_AGEMA_signal_14252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6431 ( .C (clk), .D (new_AGEMA_signal_14255), .Q (new_AGEMA_signal_14256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6435 ( .C (clk), .D (new_AGEMA_signal_14259), .Q (new_AGEMA_signal_14260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6439 ( .C (clk), .D (new_AGEMA_signal_14263), .Q (new_AGEMA_signal_14264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6443 ( .C (clk), .D (new_AGEMA_signal_14267), .Q (new_AGEMA_signal_14268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6447 ( .C (clk), .D (new_AGEMA_signal_14271), .Q (new_AGEMA_signal_14272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6451 ( .C (clk), .D (new_AGEMA_signal_14275), .Q (new_AGEMA_signal_14276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6455 ( .C (clk), .D (new_AGEMA_signal_14279), .Q (new_AGEMA_signal_14280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6459 ( .C (clk), .D (new_AGEMA_signal_14283), .Q (new_AGEMA_signal_14284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6463 ( .C (clk), .D (new_AGEMA_signal_14287), .Q (new_AGEMA_signal_14288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6467 ( .C (clk), .D (new_AGEMA_signal_14291), .Q (new_AGEMA_signal_14292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6471 ( .C (clk), .D (new_AGEMA_signal_14295), .Q (new_AGEMA_signal_14296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6475 ( .C (clk), .D (new_AGEMA_signal_14299), .Q (new_AGEMA_signal_14300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6479 ( .C (clk), .D (new_AGEMA_signal_14303), .Q (new_AGEMA_signal_14304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6483 ( .C (clk), .D (new_AGEMA_signal_14307), .Q (new_AGEMA_signal_14308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6487 ( .C (clk), .D (new_AGEMA_signal_14311), .Q (new_AGEMA_signal_14312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6491 ( .C (clk), .D (new_AGEMA_signal_14315), .Q (new_AGEMA_signal_14316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6495 ( .C (clk), .D (new_AGEMA_signal_14319), .Q (new_AGEMA_signal_14320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6499 ( .C (clk), .D (new_AGEMA_signal_14323), .Q (new_AGEMA_signal_14324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6503 ( .C (clk), .D (new_AGEMA_signal_14327), .Q (new_AGEMA_signal_14328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6507 ( .C (clk), .D (new_AGEMA_signal_14331), .Q (new_AGEMA_signal_14332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6511 ( .C (clk), .D (new_AGEMA_signal_14335), .Q (new_AGEMA_signal_14336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6515 ( .C (clk), .D (new_AGEMA_signal_14339), .Q (new_AGEMA_signal_14340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6519 ( .C (clk), .D (new_AGEMA_signal_14343), .Q (new_AGEMA_signal_14344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6523 ( .C (clk), .D (new_AGEMA_signal_14347), .Q (new_AGEMA_signal_14348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6527 ( .C (clk), .D (new_AGEMA_signal_14351), .Q (new_AGEMA_signal_14352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6531 ( .C (clk), .D (new_AGEMA_signal_14355), .Q (new_AGEMA_signal_14356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6535 ( .C (clk), .D (new_AGEMA_signal_14359), .Q (new_AGEMA_signal_14360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6539 ( .C (clk), .D (new_AGEMA_signal_14363), .Q (new_AGEMA_signal_14364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6543 ( .C (clk), .D (new_AGEMA_signal_14367), .Q (new_AGEMA_signal_14368) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6547 ( .C (clk), .D (new_AGEMA_signal_14371), .Q (new_AGEMA_signal_14372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6551 ( .C (clk), .D (new_AGEMA_signal_14375), .Q (new_AGEMA_signal_14376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6555 ( .C (clk), .D (new_AGEMA_signal_14379), .Q (new_AGEMA_signal_14380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6559 ( .C (clk), .D (new_AGEMA_signal_14383), .Q (new_AGEMA_signal_14384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6563 ( .C (clk), .D (new_AGEMA_signal_14387), .Q (new_AGEMA_signal_14388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6567 ( .C (clk), .D (new_AGEMA_signal_14391), .Q (new_AGEMA_signal_14392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6571 ( .C (clk), .D (new_AGEMA_signal_14395), .Q (new_AGEMA_signal_14396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6575 ( .C (clk), .D (new_AGEMA_signal_14399), .Q (new_AGEMA_signal_14400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6579 ( .C (clk), .D (new_AGEMA_signal_14403), .Q (new_AGEMA_signal_14404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6583 ( .C (clk), .D (new_AGEMA_signal_14407), .Q (new_AGEMA_signal_14408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6587 ( .C (clk), .D (new_AGEMA_signal_14411), .Q (new_AGEMA_signal_14412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6591 ( .C (clk), .D (new_AGEMA_signal_14415), .Q (new_AGEMA_signal_14416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6595 ( .C (clk), .D (new_AGEMA_signal_14419), .Q (new_AGEMA_signal_14420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6599 ( .C (clk), .D (new_AGEMA_signal_14423), .Q (new_AGEMA_signal_14424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6603 ( .C (clk), .D (new_AGEMA_signal_14427), .Q (new_AGEMA_signal_14428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6607 ( .C (clk), .D (new_AGEMA_signal_14431), .Q (new_AGEMA_signal_14432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6611 ( .C (clk), .D (new_AGEMA_signal_14435), .Q (new_AGEMA_signal_14436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6615 ( .C (clk), .D (new_AGEMA_signal_14439), .Q (new_AGEMA_signal_14440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6619 ( .C (clk), .D (new_AGEMA_signal_14443), .Q (new_AGEMA_signal_14444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6623 ( .C (clk), .D (new_AGEMA_signal_14447), .Q (new_AGEMA_signal_14448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6627 ( .C (clk), .D (new_AGEMA_signal_14451), .Q (new_AGEMA_signal_14452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6631 ( .C (clk), .D (new_AGEMA_signal_14455), .Q (new_AGEMA_signal_14456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6635 ( .C (clk), .D (new_AGEMA_signal_14459), .Q (new_AGEMA_signal_14460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6639 ( .C (clk), .D (new_AGEMA_signal_14463), .Q (new_AGEMA_signal_14464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6643 ( .C (clk), .D (new_AGEMA_signal_14467), .Q (new_AGEMA_signal_14468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6647 ( .C (clk), .D (new_AGEMA_signal_14471), .Q (new_AGEMA_signal_14472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6651 ( .C (clk), .D (new_AGEMA_signal_14475), .Q (new_AGEMA_signal_14476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6655 ( .C (clk), .D (new_AGEMA_signal_14479), .Q (new_AGEMA_signal_14480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6659 ( .C (clk), .D (new_AGEMA_signal_14483), .Q (new_AGEMA_signal_14484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6663 ( .C (clk), .D (new_AGEMA_signal_14487), .Q (new_AGEMA_signal_14488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6667 ( .C (clk), .D (new_AGEMA_signal_14491), .Q (new_AGEMA_signal_14492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6671 ( .C (clk), .D (new_AGEMA_signal_14495), .Q (new_AGEMA_signal_14496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6675 ( .C (clk), .D (new_AGEMA_signal_14499), .Q (new_AGEMA_signal_14500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6679 ( .C (clk), .D (new_AGEMA_signal_14503), .Q (new_AGEMA_signal_14504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6683 ( .C (clk), .D (new_AGEMA_signal_14507), .Q (new_AGEMA_signal_14508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6687 ( .C (clk), .D (new_AGEMA_signal_14511), .Q (new_AGEMA_signal_14512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6691 ( .C (clk), .D (new_AGEMA_signal_14515), .Q (new_AGEMA_signal_14516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6695 ( .C (clk), .D (new_AGEMA_signal_14519), .Q (new_AGEMA_signal_14520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6699 ( .C (clk), .D (new_AGEMA_signal_14523), .Q (new_AGEMA_signal_14524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6703 ( .C (clk), .D (new_AGEMA_signal_14527), .Q (new_AGEMA_signal_14528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6707 ( .C (clk), .D (new_AGEMA_signal_14531), .Q (new_AGEMA_signal_14532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6711 ( .C (clk), .D (new_AGEMA_signal_14535), .Q (new_AGEMA_signal_14536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6715 ( .C (clk), .D (new_AGEMA_signal_14539), .Q (new_AGEMA_signal_14540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6719 ( .C (clk), .D (new_AGEMA_signal_14543), .Q (new_AGEMA_signal_14544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6723 ( .C (clk), .D (new_AGEMA_signal_14547), .Q (new_AGEMA_signal_14548) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6727 ( .C (clk), .D (new_AGEMA_signal_14551), .Q (new_AGEMA_signal_14552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6731 ( .C (clk), .D (new_AGEMA_signal_14555), .Q (new_AGEMA_signal_14556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6735 ( .C (clk), .D (new_AGEMA_signal_14559), .Q (new_AGEMA_signal_14560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6739 ( .C (clk), .D (new_AGEMA_signal_14563), .Q (new_AGEMA_signal_14564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6743 ( .C (clk), .D (new_AGEMA_signal_14567), .Q (new_AGEMA_signal_14568) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6747 ( .C (clk), .D (new_AGEMA_signal_14571), .Q (new_AGEMA_signal_14572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6751 ( .C (clk), .D (new_AGEMA_signal_14575), .Q (new_AGEMA_signal_14576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6755 ( .C (clk), .D (new_AGEMA_signal_14579), .Q (new_AGEMA_signal_14580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6759 ( .C (clk), .D (new_AGEMA_signal_14583), .Q (new_AGEMA_signal_14584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6763 ( .C (clk), .D (new_AGEMA_signal_14587), .Q (new_AGEMA_signal_14588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6767 ( .C (clk), .D (new_AGEMA_signal_14591), .Q (new_AGEMA_signal_14592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6771 ( .C (clk), .D (new_AGEMA_signal_14595), .Q (new_AGEMA_signal_14596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6775 ( .C (clk), .D (new_AGEMA_signal_14599), .Q (new_AGEMA_signal_14600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6779 ( .C (clk), .D (new_AGEMA_signal_14603), .Q (new_AGEMA_signal_14604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6783 ( .C (clk), .D (new_AGEMA_signal_14607), .Q (new_AGEMA_signal_14608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6787 ( .C (clk), .D (new_AGEMA_signal_14611), .Q (new_AGEMA_signal_14612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6791 ( .C (clk), .D (new_AGEMA_signal_14615), .Q (new_AGEMA_signal_14616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6795 ( .C (clk), .D (new_AGEMA_signal_14619), .Q (new_AGEMA_signal_14620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6799 ( .C (clk), .D (new_AGEMA_signal_14623), .Q (new_AGEMA_signal_14624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6803 ( .C (clk), .D (new_AGEMA_signal_14627), .Q (new_AGEMA_signal_14628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6807 ( .C (clk), .D (new_AGEMA_signal_14631), .Q (new_AGEMA_signal_14632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6811 ( .C (clk), .D (new_AGEMA_signal_14635), .Q (new_AGEMA_signal_14636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6815 ( .C (clk), .D (new_AGEMA_signal_14639), .Q (new_AGEMA_signal_14640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6819 ( .C (clk), .D (new_AGEMA_signal_14643), .Q (new_AGEMA_signal_14644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6823 ( .C (clk), .D (new_AGEMA_signal_14647), .Q (new_AGEMA_signal_14648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6827 ( .C (clk), .D (new_AGEMA_signal_14651), .Q (new_AGEMA_signal_14652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6831 ( .C (clk), .D (new_AGEMA_signal_14655), .Q (new_AGEMA_signal_14656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6835 ( .C (clk), .D (new_AGEMA_signal_14659), .Q (new_AGEMA_signal_14660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6839 ( .C (clk), .D (new_AGEMA_signal_14663), .Q (new_AGEMA_signal_14664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6843 ( .C (clk), .D (new_AGEMA_signal_14667), .Q (new_AGEMA_signal_14668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6847 ( .C (clk), .D (new_AGEMA_signal_14671), .Q (new_AGEMA_signal_14672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6851 ( .C (clk), .D (new_AGEMA_signal_14675), .Q (new_AGEMA_signal_14676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6855 ( .C (clk), .D (new_AGEMA_signal_14679), .Q (new_AGEMA_signal_14680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6859 ( .C (clk), .D (new_AGEMA_signal_14683), .Q (new_AGEMA_signal_14684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6863 ( .C (clk), .D (new_AGEMA_signal_14687), .Q (new_AGEMA_signal_14688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6867 ( .C (clk), .D (new_AGEMA_signal_14691), .Q (new_AGEMA_signal_14692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6871 ( .C (clk), .D (new_AGEMA_signal_14695), .Q (new_AGEMA_signal_14696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6875 ( .C (clk), .D (new_AGEMA_signal_14699), .Q (new_AGEMA_signal_14700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6879 ( .C (clk), .D (new_AGEMA_signal_14703), .Q (new_AGEMA_signal_14704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6883 ( .C (clk), .D (new_AGEMA_signal_14707), .Q (new_AGEMA_signal_14708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6887 ( .C (clk), .D (new_AGEMA_signal_14711), .Q (new_AGEMA_signal_14712) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6891 ( .C (clk), .D (new_AGEMA_signal_14715), .Q (new_AGEMA_signal_14716) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6895 ( .C (clk), .D (new_AGEMA_signal_14719), .Q (new_AGEMA_signal_14720) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6899 ( .C (clk), .D (new_AGEMA_signal_14723), .Q (new_AGEMA_signal_14724) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6903 ( .C (clk), .D (new_AGEMA_signal_14727), .Q (new_AGEMA_signal_14728) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6907 ( .C (clk), .D (new_AGEMA_signal_14731), .Q (new_AGEMA_signal_14732) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6911 ( .C (clk), .D (new_AGEMA_signal_14735), .Q (new_AGEMA_signal_14736) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6915 ( .C (clk), .D (new_AGEMA_signal_14739), .Q (new_AGEMA_signal_14740) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6919 ( .C (clk), .D (new_AGEMA_signal_14743), .Q (new_AGEMA_signal_14744) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6923 ( .C (clk), .D (new_AGEMA_signal_14747), .Q (new_AGEMA_signal_14748) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6927 ( .C (clk), .D (new_AGEMA_signal_14751), .Q (new_AGEMA_signal_14752) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6931 ( .C (clk), .D (new_AGEMA_signal_14755), .Q (new_AGEMA_signal_14756) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6935 ( .C (clk), .D (new_AGEMA_signal_14759), .Q (new_AGEMA_signal_14760) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6939 ( .C (clk), .D (new_AGEMA_signal_14763), .Q (new_AGEMA_signal_14764) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6943 ( .C (clk), .D (new_AGEMA_signal_14767), .Q (new_AGEMA_signal_14768) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6947 ( .C (clk), .D (new_AGEMA_signal_14771), .Q (new_AGEMA_signal_14772) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6951 ( .C (clk), .D (new_AGEMA_signal_14775), .Q (new_AGEMA_signal_14776) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6955 ( .C (clk), .D (new_AGEMA_signal_14779), .Q (new_AGEMA_signal_14780) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6959 ( .C (clk), .D (new_AGEMA_signal_14783), .Q (new_AGEMA_signal_14784) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6963 ( .C (clk), .D (new_AGEMA_signal_14787), .Q (new_AGEMA_signal_14788) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6967 ( .C (clk), .D (new_AGEMA_signal_14791), .Q (new_AGEMA_signal_14792) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6971 ( .C (clk), .D (new_AGEMA_signal_14795), .Q (new_AGEMA_signal_14796) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6975 ( .C (clk), .D (new_AGEMA_signal_14799), .Q (new_AGEMA_signal_14800) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6979 ( .C (clk), .D (new_AGEMA_signal_14803), .Q (new_AGEMA_signal_14804) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6983 ( .C (clk), .D (new_AGEMA_signal_14807), .Q (new_AGEMA_signal_14808) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6987 ( .C (clk), .D (new_AGEMA_signal_14811), .Q (new_AGEMA_signal_14812) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6991 ( .C (clk), .D (new_AGEMA_signal_14815), .Q (new_AGEMA_signal_14816) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6995 ( .C (clk), .D (new_AGEMA_signal_14819), .Q (new_AGEMA_signal_14820) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6999 ( .C (clk), .D (new_AGEMA_signal_14823), .Q (new_AGEMA_signal_14824) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7003 ( .C (clk), .D (new_AGEMA_signal_14827), .Q (new_AGEMA_signal_14828) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7007 ( .C (clk), .D (new_AGEMA_signal_14831), .Q (new_AGEMA_signal_14832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7011 ( .C (clk), .D (new_AGEMA_signal_14835), .Q (new_AGEMA_signal_14836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7015 ( .C (clk), .D (new_AGEMA_signal_14839), .Q (new_AGEMA_signal_14840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7019 ( .C (clk), .D (new_AGEMA_signal_14843), .Q (new_AGEMA_signal_14844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7023 ( .C (clk), .D (new_AGEMA_signal_14847), .Q (new_AGEMA_signal_14848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7027 ( .C (clk), .D (new_AGEMA_signal_14851), .Q (new_AGEMA_signal_14852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7031 ( .C (clk), .D (new_AGEMA_signal_14855), .Q (new_AGEMA_signal_14856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7035 ( .C (clk), .D (new_AGEMA_signal_14859), .Q (new_AGEMA_signal_14860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7039 ( .C (clk), .D (new_AGEMA_signal_14863), .Q (new_AGEMA_signal_14864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7043 ( .C (clk), .D (new_AGEMA_signal_14867), .Q (new_AGEMA_signal_14868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7047 ( .C (clk), .D (new_AGEMA_signal_14871), .Q (new_AGEMA_signal_14872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7051 ( .C (clk), .D (new_AGEMA_signal_14875), .Q (new_AGEMA_signal_14876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7055 ( .C (clk), .D (new_AGEMA_signal_14879), .Q (new_AGEMA_signal_14880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7059 ( .C (clk), .D (new_AGEMA_signal_14883), .Q (new_AGEMA_signal_14884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7063 ( .C (clk), .D (new_AGEMA_signal_14887), .Q (new_AGEMA_signal_14888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7067 ( .C (clk), .D (new_AGEMA_signal_14891), .Q (new_AGEMA_signal_14892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7071 ( .C (clk), .D (new_AGEMA_signal_14895), .Q (new_AGEMA_signal_14896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7075 ( .C (clk), .D (new_AGEMA_signal_14899), .Q (new_AGEMA_signal_14900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7079 ( .C (clk), .D (new_AGEMA_signal_14903), .Q (new_AGEMA_signal_14904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7083 ( .C (clk), .D (new_AGEMA_signal_14907), .Q (new_AGEMA_signal_14908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7087 ( .C (clk), .D (new_AGEMA_signal_14911), .Q (new_AGEMA_signal_14912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7091 ( .C (clk), .D (new_AGEMA_signal_14915), .Q (new_AGEMA_signal_14916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7095 ( .C (clk), .D (new_AGEMA_signal_14919), .Q (new_AGEMA_signal_14920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7099 ( .C (clk), .D (new_AGEMA_signal_14923), .Q (new_AGEMA_signal_14924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7103 ( .C (clk), .D (new_AGEMA_signal_14927), .Q (new_AGEMA_signal_14928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7107 ( .C (clk), .D (new_AGEMA_signal_14931), .Q (new_AGEMA_signal_14932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7111 ( .C (clk), .D (new_AGEMA_signal_14935), .Q (new_AGEMA_signal_14936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7115 ( .C (clk), .D (new_AGEMA_signal_14939), .Q (new_AGEMA_signal_14940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7119 ( .C (clk), .D (new_AGEMA_signal_14943), .Q (new_AGEMA_signal_14944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7123 ( .C (clk), .D (new_AGEMA_signal_14947), .Q (new_AGEMA_signal_14948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7127 ( .C (clk), .D (new_AGEMA_signal_14951), .Q (new_AGEMA_signal_14952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7131 ( .C (clk), .D (new_AGEMA_signal_14955), .Q (new_AGEMA_signal_14956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7135 ( .C (clk), .D (new_AGEMA_signal_14959), .Q (new_AGEMA_signal_14960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7139 ( .C (clk), .D (new_AGEMA_signal_14963), .Q (new_AGEMA_signal_14964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7143 ( .C (clk), .D (new_AGEMA_signal_14967), .Q (new_AGEMA_signal_14968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7147 ( .C (clk), .D (new_AGEMA_signal_14971), .Q (new_AGEMA_signal_14972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7151 ( .C (clk), .D (new_AGEMA_signal_14975), .Q (new_AGEMA_signal_14976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7155 ( .C (clk), .D (new_AGEMA_signal_14979), .Q (new_AGEMA_signal_14980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7159 ( .C (clk), .D (new_AGEMA_signal_14983), .Q (new_AGEMA_signal_14984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7163 ( .C (clk), .D (new_AGEMA_signal_14987), .Q (new_AGEMA_signal_14988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7167 ( .C (clk), .D (new_AGEMA_signal_14991), .Q (new_AGEMA_signal_14992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7171 ( .C (clk), .D (new_AGEMA_signal_14995), .Q (new_AGEMA_signal_14996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7175 ( .C (clk), .D (new_AGEMA_signal_14999), .Q (new_AGEMA_signal_15000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7179 ( .C (clk), .D (new_AGEMA_signal_15003), .Q (new_AGEMA_signal_15004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7183 ( .C (clk), .D (new_AGEMA_signal_15007), .Q (new_AGEMA_signal_15008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7187 ( .C (clk), .D (new_AGEMA_signal_15011), .Q (new_AGEMA_signal_15012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7191 ( .C (clk), .D (new_AGEMA_signal_15015), .Q (new_AGEMA_signal_15016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7195 ( .C (clk), .D (new_AGEMA_signal_15019), .Q (new_AGEMA_signal_15020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7199 ( .C (clk), .D (new_AGEMA_signal_15023), .Q (new_AGEMA_signal_15024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7203 ( .C (clk), .D (new_AGEMA_signal_15027), .Q (new_AGEMA_signal_15028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7207 ( .C (clk), .D (new_AGEMA_signal_15031), .Q (new_AGEMA_signal_15032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7211 ( .C (clk), .D (new_AGEMA_signal_15035), .Q (new_AGEMA_signal_15036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7215 ( .C (clk), .D (new_AGEMA_signal_15039), .Q (new_AGEMA_signal_15040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7219 ( .C (clk), .D (new_AGEMA_signal_15043), .Q (new_AGEMA_signal_15044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7223 ( .C (clk), .D (new_AGEMA_signal_15047), .Q (new_AGEMA_signal_15048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7227 ( .C (clk), .D (new_AGEMA_signal_15051), .Q (new_AGEMA_signal_15052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7231 ( .C (clk), .D (new_AGEMA_signal_15055), .Q (new_AGEMA_signal_15056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7235 ( .C (clk), .D (new_AGEMA_signal_15059), .Q (new_AGEMA_signal_15060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7239 ( .C (clk), .D (new_AGEMA_signal_15063), .Q (new_AGEMA_signal_15064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7243 ( .C (clk), .D (new_AGEMA_signal_15067), .Q (new_AGEMA_signal_15068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7247 ( .C (clk), .D (new_AGEMA_signal_15071), .Q (new_AGEMA_signal_15072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7251 ( .C (clk), .D (new_AGEMA_signal_15075), .Q (new_AGEMA_signal_15076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7255 ( .C (clk), .D (new_AGEMA_signal_15079), .Q (new_AGEMA_signal_15080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7259 ( .C (clk), .D (new_AGEMA_signal_15083), .Q (new_AGEMA_signal_15084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7263 ( .C (clk), .D (new_AGEMA_signal_15087), .Q (new_AGEMA_signal_15088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7267 ( .C (clk), .D (new_AGEMA_signal_15091), .Q (new_AGEMA_signal_15092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7271 ( .C (clk), .D (new_AGEMA_signal_15095), .Q (new_AGEMA_signal_15096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7275 ( .C (clk), .D (new_AGEMA_signal_15099), .Q (new_AGEMA_signal_15100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7279 ( .C (clk), .D (new_AGEMA_signal_15103), .Q (new_AGEMA_signal_15104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7283 ( .C (clk), .D (new_AGEMA_signal_15107), .Q (new_AGEMA_signal_15108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7287 ( .C (clk), .D (new_AGEMA_signal_15111), .Q (new_AGEMA_signal_15112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7291 ( .C (clk), .D (new_AGEMA_signal_15115), .Q (new_AGEMA_signal_15116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7295 ( .C (clk), .D (new_AGEMA_signal_15119), .Q (new_AGEMA_signal_15120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7299 ( .C (clk), .D (new_AGEMA_signal_15123), .Q (new_AGEMA_signal_15124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7303 ( .C (clk), .D (new_AGEMA_signal_15127), .Q (new_AGEMA_signal_15128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7307 ( .C (clk), .D (new_AGEMA_signal_15131), .Q (new_AGEMA_signal_15132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7311 ( .C (clk), .D (new_AGEMA_signal_15135), .Q (new_AGEMA_signal_15136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7315 ( .C (clk), .D (new_AGEMA_signal_15139), .Q (new_AGEMA_signal_15140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7319 ( .C (clk), .D (new_AGEMA_signal_15143), .Q (new_AGEMA_signal_15144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7323 ( .C (clk), .D (new_AGEMA_signal_15147), .Q (new_AGEMA_signal_15148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7327 ( .C (clk), .D (new_AGEMA_signal_15151), .Q (new_AGEMA_signal_15152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7331 ( .C (clk), .D (new_AGEMA_signal_15155), .Q (new_AGEMA_signal_15156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7335 ( .C (clk), .D (new_AGEMA_signal_15159), .Q (new_AGEMA_signal_15160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7339 ( .C (clk), .D (new_AGEMA_signal_15163), .Q (new_AGEMA_signal_15164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7343 ( .C (clk), .D (new_AGEMA_signal_15167), .Q (new_AGEMA_signal_15168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7347 ( .C (clk), .D (new_AGEMA_signal_15171), .Q (new_AGEMA_signal_15172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7351 ( .C (clk), .D (new_AGEMA_signal_15175), .Q (new_AGEMA_signal_15176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7355 ( .C (clk), .D (new_AGEMA_signal_15179), .Q (new_AGEMA_signal_15180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7359 ( .C (clk), .D (new_AGEMA_signal_15183), .Q (new_AGEMA_signal_15184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7363 ( .C (clk), .D (new_AGEMA_signal_15187), .Q (new_AGEMA_signal_15188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7367 ( .C (clk), .D (new_AGEMA_signal_15191), .Q (new_AGEMA_signal_15192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7371 ( .C (clk), .D (new_AGEMA_signal_15195), .Q (new_AGEMA_signal_15196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7375 ( .C (clk), .D (new_AGEMA_signal_15199), .Q (new_AGEMA_signal_15200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7379 ( .C (clk), .D (new_AGEMA_signal_15203), .Q (new_AGEMA_signal_15204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7383 ( .C (clk), .D (new_AGEMA_signal_15207), .Q (new_AGEMA_signal_15208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7387 ( .C (clk), .D (new_AGEMA_signal_15211), .Q (new_AGEMA_signal_15212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7391 ( .C (clk), .D (new_AGEMA_signal_15215), .Q (new_AGEMA_signal_15216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7395 ( .C (clk), .D (new_AGEMA_signal_15219), .Q (new_AGEMA_signal_15220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7399 ( .C (clk), .D (new_AGEMA_signal_15223), .Q (new_AGEMA_signal_15224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7403 ( .C (clk), .D (new_AGEMA_signal_15227), .Q (new_AGEMA_signal_15228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7407 ( .C (clk), .D (new_AGEMA_signal_15231), .Q (new_AGEMA_signal_15232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7411 ( .C (clk), .D (new_AGEMA_signal_15235), .Q (new_AGEMA_signal_15236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7415 ( .C (clk), .D (new_AGEMA_signal_15239), .Q (new_AGEMA_signal_15240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7419 ( .C (clk), .D (new_AGEMA_signal_15243), .Q (new_AGEMA_signal_15244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7423 ( .C (clk), .D (new_AGEMA_signal_15247), .Q (new_AGEMA_signal_15248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7427 ( .C (clk), .D (new_AGEMA_signal_15251), .Q (new_AGEMA_signal_15252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7431 ( .C (clk), .D (new_AGEMA_signal_15255), .Q (new_AGEMA_signal_15256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7435 ( .C (clk), .D (new_AGEMA_signal_15259), .Q (new_AGEMA_signal_15260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7439 ( .C (clk), .D (new_AGEMA_signal_15263), .Q (new_AGEMA_signal_15264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7443 ( .C (clk), .D (new_AGEMA_signal_15267), .Q (new_AGEMA_signal_15268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7447 ( .C (clk), .D (new_AGEMA_signal_15271), .Q (new_AGEMA_signal_15272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7451 ( .C (clk), .D (new_AGEMA_signal_15275), .Q (new_AGEMA_signal_15276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7455 ( .C (clk), .D (new_AGEMA_signal_15279), .Q (new_AGEMA_signal_15280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7459 ( .C (clk), .D (new_AGEMA_signal_15283), .Q (new_AGEMA_signal_15284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7463 ( .C (clk), .D (new_AGEMA_signal_15287), .Q (new_AGEMA_signal_15288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7467 ( .C (clk), .D (new_AGEMA_signal_15291), .Q (new_AGEMA_signal_15292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7471 ( .C (clk), .D (new_AGEMA_signal_15295), .Q (new_AGEMA_signal_15296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7475 ( .C (clk), .D (new_AGEMA_signal_15299), .Q (new_AGEMA_signal_15300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7479 ( .C (clk), .D (new_AGEMA_signal_15303), .Q (new_AGEMA_signal_15304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7483 ( .C (clk), .D (new_AGEMA_signal_15307), .Q (new_AGEMA_signal_15308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7487 ( .C (clk), .D (new_AGEMA_signal_15311), .Q (new_AGEMA_signal_15312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7491 ( .C (clk), .D (new_AGEMA_signal_15315), .Q (new_AGEMA_signal_15316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7495 ( .C (clk), .D (new_AGEMA_signal_15319), .Q (new_AGEMA_signal_15320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7499 ( .C (clk), .D (new_AGEMA_signal_15323), .Q (new_AGEMA_signal_15324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7503 ( .C (clk), .D (new_AGEMA_signal_15327), .Q (new_AGEMA_signal_15328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7507 ( .C (clk), .D (new_AGEMA_signal_15331), .Q (new_AGEMA_signal_15332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7511 ( .C (clk), .D (new_AGEMA_signal_15335), .Q (new_AGEMA_signal_15336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7515 ( .C (clk), .D (new_AGEMA_signal_15339), .Q (new_AGEMA_signal_15340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7519 ( .C (clk), .D (new_AGEMA_signal_15343), .Q (new_AGEMA_signal_15344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7523 ( .C (clk), .D (new_AGEMA_signal_15347), .Q (new_AGEMA_signal_15348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7527 ( .C (clk), .D (new_AGEMA_signal_15351), .Q (new_AGEMA_signal_15352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7531 ( .C (clk), .D (new_AGEMA_signal_15355), .Q (new_AGEMA_signal_15356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7535 ( .C (clk), .D (new_AGEMA_signal_15359), .Q (new_AGEMA_signal_15360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7539 ( .C (clk), .D (new_AGEMA_signal_15363), .Q (new_AGEMA_signal_15364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7543 ( .C (clk), .D (new_AGEMA_signal_15367), .Q (new_AGEMA_signal_15368) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7547 ( .C (clk), .D (new_AGEMA_signal_15371), .Q (new_AGEMA_signal_15372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7551 ( .C (clk), .D (new_AGEMA_signal_15375), .Q (new_AGEMA_signal_15376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7555 ( .C (clk), .D (new_AGEMA_signal_15379), .Q (new_AGEMA_signal_15380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7559 ( .C (clk), .D (new_AGEMA_signal_15383), .Q (new_AGEMA_signal_15384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7563 ( .C (clk), .D (new_AGEMA_signal_15387), .Q (new_AGEMA_signal_15388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7567 ( .C (clk), .D (new_AGEMA_signal_15391), .Q (new_AGEMA_signal_15392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7571 ( .C (clk), .D (new_AGEMA_signal_15395), .Q (new_AGEMA_signal_15396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7575 ( .C (clk), .D (new_AGEMA_signal_15399), .Q (new_AGEMA_signal_15400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7579 ( .C (clk), .D (new_AGEMA_signal_15403), .Q (new_AGEMA_signal_15404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7583 ( .C (clk), .D (new_AGEMA_signal_15407), .Q (new_AGEMA_signal_15408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7587 ( .C (clk), .D (new_AGEMA_signal_15411), .Q (new_AGEMA_signal_15412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7591 ( .C (clk), .D (new_AGEMA_signal_15415), .Q (new_AGEMA_signal_15416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7595 ( .C (clk), .D (new_AGEMA_signal_15419), .Q (new_AGEMA_signal_15420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7599 ( .C (clk), .D (new_AGEMA_signal_15423), .Q (new_AGEMA_signal_15424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7603 ( .C (clk), .D (new_AGEMA_signal_15427), .Q (new_AGEMA_signal_15428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7607 ( .C (clk), .D (new_AGEMA_signal_15431), .Q (new_AGEMA_signal_15432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7611 ( .C (clk), .D (new_AGEMA_signal_15435), .Q (new_AGEMA_signal_15436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7615 ( .C (clk), .D (new_AGEMA_signal_15439), .Q (new_AGEMA_signal_15440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7619 ( .C (clk), .D (new_AGEMA_signal_15443), .Q (new_AGEMA_signal_15444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7623 ( .C (clk), .D (new_AGEMA_signal_15447), .Q (new_AGEMA_signal_15448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7627 ( .C (clk), .D (new_AGEMA_signal_15451), .Q (new_AGEMA_signal_15452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7631 ( .C (clk), .D (new_AGEMA_signal_15455), .Q (new_AGEMA_signal_15456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7635 ( .C (clk), .D (new_AGEMA_signal_15459), .Q (new_AGEMA_signal_15460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7639 ( .C (clk), .D (new_AGEMA_signal_15463), .Q (new_AGEMA_signal_15464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7643 ( .C (clk), .D (new_AGEMA_signal_15467), .Q (new_AGEMA_signal_15468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7647 ( .C (clk), .D (new_AGEMA_signal_15471), .Q (new_AGEMA_signal_15472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7651 ( .C (clk), .D (new_AGEMA_signal_15475), .Q (new_AGEMA_signal_15476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7655 ( .C (clk), .D (new_AGEMA_signal_15479), .Q (new_AGEMA_signal_15480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7659 ( .C (clk), .D (new_AGEMA_signal_15483), .Q (new_AGEMA_signal_15484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7663 ( .C (clk), .D (new_AGEMA_signal_15487), .Q (new_AGEMA_signal_15488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7667 ( .C (clk), .D (new_AGEMA_signal_15491), .Q (new_AGEMA_signal_15492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7671 ( .C (clk), .D (new_AGEMA_signal_15495), .Q (new_AGEMA_signal_15496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7675 ( .C (clk), .D (new_AGEMA_signal_15499), .Q (new_AGEMA_signal_15500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7679 ( .C (clk), .D (new_AGEMA_signal_15503), .Q (new_AGEMA_signal_15504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7683 ( .C (clk), .D (new_AGEMA_signal_15507), .Q (new_AGEMA_signal_15508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7687 ( .C (clk), .D (new_AGEMA_signal_15511), .Q (new_AGEMA_signal_15512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7691 ( .C (clk), .D (new_AGEMA_signal_15515), .Q (new_AGEMA_signal_15516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7695 ( .C (clk), .D (new_AGEMA_signal_15519), .Q (new_AGEMA_signal_15520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7699 ( .C (clk), .D (new_AGEMA_signal_15523), .Q (new_AGEMA_signal_15524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7703 ( .C (clk), .D (new_AGEMA_signal_15527), .Q (new_AGEMA_signal_15528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7707 ( .C (clk), .D (new_AGEMA_signal_15531), .Q (new_AGEMA_signal_15532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7711 ( .C (clk), .D (new_AGEMA_signal_15535), .Q (new_AGEMA_signal_15536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7715 ( .C (clk), .D (new_AGEMA_signal_15539), .Q (new_AGEMA_signal_15540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7719 ( .C (clk), .D (new_AGEMA_signal_15543), .Q (new_AGEMA_signal_15544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7723 ( .C (clk), .D (new_AGEMA_signal_15547), .Q (new_AGEMA_signal_15548) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7727 ( .C (clk), .D (new_AGEMA_signal_15551), .Q (new_AGEMA_signal_15552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7731 ( .C (clk), .D (new_AGEMA_signal_15555), .Q (new_AGEMA_signal_15556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7735 ( .C (clk), .D (new_AGEMA_signal_15559), .Q (new_AGEMA_signal_15560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7739 ( .C (clk), .D (new_AGEMA_signal_15563), .Q (new_AGEMA_signal_15564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7743 ( .C (clk), .D (new_AGEMA_signal_15567), .Q (new_AGEMA_signal_15568) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7747 ( .C (clk), .D (new_AGEMA_signal_15571), .Q (new_AGEMA_signal_15572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7751 ( .C (clk), .D (new_AGEMA_signal_15575), .Q (new_AGEMA_signal_15576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7755 ( .C (clk), .D (new_AGEMA_signal_15579), .Q (new_AGEMA_signal_15580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7759 ( .C (clk), .D (new_AGEMA_signal_15583), .Q (new_AGEMA_signal_15584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7763 ( .C (clk), .D (new_AGEMA_signal_15587), .Q (new_AGEMA_signal_15588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7767 ( .C (clk), .D (new_AGEMA_signal_15591), .Q (new_AGEMA_signal_15592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7771 ( .C (clk), .D (new_AGEMA_signal_15595), .Q (new_AGEMA_signal_15596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7775 ( .C (clk), .D (new_AGEMA_signal_15599), .Q (new_AGEMA_signal_15600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7779 ( .C (clk), .D (new_AGEMA_signal_15603), .Q (new_AGEMA_signal_15604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7783 ( .C (clk), .D (new_AGEMA_signal_15607), .Q (new_AGEMA_signal_15608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7787 ( .C (clk), .D (new_AGEMA_signal_15611), .Q (new_AGEMA_signal_15612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7791 ( .C (clk), .D (new_AGEMA_signal_15615), .Q (new_AGEMA_signal_15616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7795 ( .C (clk), .D (new_AGEMA_signal_15619), .Q (new_AGEMA_signal_15620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7799 ( .C (clk), .D (new_AGEMA_signal_15623), .Q (new_AGEMA_signal_15624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7803 ( .C (clk), .D (new_AGEMA_signal_15627), .Q (new_AGEMA_signal_15628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7807 ( .C (clk), .D (new_AGEMA_signal_15631), .Q (new_AGEMA_signal_15632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7811 ( .C (clk), .D (new_AGEMA_signal_15635), .Q (new_AGEMA_signal_15636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7815 ( .C (clk), .D (new_AGEMA_signal_15639), .Q (new_AGEMA_signal_15640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7819 ( .C (clk), .D (new_AGEMA_signal_15643), .Q (new_AGEMA_signal_15644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7823 ( .C (clk), .D (new_AGEMA_signal_15647), .Q (new_AGEMA_signal_15648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7827 ( .C (clk), .D (new_AGEMA_signal_15651), .Q (new_AGEMA_signal_15652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7831 ( .C (clk), .D (new_AGEMA_signal_15655), .Q (new_AGEMA_signal_15656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7835 ( .C (clk), .D (new_AGEMA_signal_15659), .Q (new_AGEMA_signal_15660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7839 ( .C (clk), .D (new_AGEMA_signal_15663), .Q (new_AGEMA_signal_15664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7843 ( .C (clk), .D (new_AGEMA_signal_15667), .Q (new_AGEMA_signal_15668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7847 ( .C (clk), .D (new_AGEMA_signal_15671), .Q (new_AGEMA_signal_15672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7851 ( .C (clk), .D (new_AGEMA_signal_15675), .Q (new_AGEMA_signal_15676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7855 ( .C (clk), .D (new_AGEMA_signal_15679), .Q (new_AGEMA_signal_15680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7859 ( .C (clk), .D (new_AGEMA_signal_15683), .Q (new_AGEMA_signal_15684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7863 ( .C (clk), .D (new_AGEMA_signal_15687), .Q (new_AGEMA_signal_15688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7867 ( .C (clk), .D (new_AGEMA_signal_15691), .Q (new_AGEMA_signal_15692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7871 ( .C (clk), .D (new_AGEMA_signal_15695), .Q (new_AGEMA_signal_15696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7875 ( .C (clk), .D (new_AGEMA_signal_15699), .Q (new_AGEMA_signal_15700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7879 ( .C (clk), .D (new_AGEMA_signal_15703), .Q (new_AGEMA_signal_15704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7883 ( .C (clk), .D (new_AGEMA_signal_15707), .Q (new_AGEMA_signal_15708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7887 ( .C (clk), .D (new_AGEMA_signal_15711), .Q (new_AGEMA_signal_15712) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7891 ( .C (clk), .D (new_AGEMA_signal_15715), .Q (new_AGEMA_signal_15716) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7895 ( .C (clk), .D (new_AGEMA_signal_15719), .Q (new_AGEMA_signal_15720) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7899 ( .C (clk), .D (new_AGEMA_signal_15723), .Q (new_AGEMA_signal_15724) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7903 ( .C (clk), .D (new_AGEMA_signal_15727), .Q (new_AGEMA_signal_15728) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7907 ( .C (clk), .D (new_AGEMA_signal_15731), .Q (new_AGEMA_signal_15732) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7911 ( .C (clk), .D (new_AGEMA_signal_15735), .Q (new_AGEMA_signal_15736) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7915 ( .C (clk), .D (new_AGEMA_signal_15739), .Q (new_AGEMA_signal_15740) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7919 ( .C (clk), .D (new_AGEMA_signal_15743), .Q (new_AGEMA_signal_15744) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7923 ( .C (clk), .D (new_AGEMA_signal_15747), .Q (new_AGEMA_signal_15748) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7927 ( .C (clk), .D (new_AGEMA_signal_15751), .Q (new_AGEMA_signal_15752) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7931 ( .C (clk), .D (new_AGEMA_signal_15755), .Q (new_AGEMA_signal_15756) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7935 ( .C (clk), .D (new_AGEMA_signal_15759), .Q (new_AGEMA_signal_15760) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7939 ( .C (clk), .D (new_AGEMA_signal_15763), .Q (new_AGEMA_signal_15764) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7943 ( .C (clk), .D (new_AGEMA_signal_15767), .Q (new_AGEMA_signal_15768) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7947 ( .C (clk), .D (new_AGEMA_signal_15771), .Q (new_AGEMA_signal_15772) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7951 ( .C (clk), .D (new_AGEMA_signal_15775), .Q (new_AGEMA_signal_15776) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7955 ( .C (clk), .D (new_AGEMA_signal_15779), .Q (new_AGEMA_signal_15780) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7959 ( .C (clk), .D (new_AGEMA_signal_15783), .Q (new_AGEMA_signal_15784) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7963 ( .C (clk), .D (new_AGEMA_signal_15787), .Q (new_AGEMA_signal_15788) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7967 ( .C (clk), .D (new_AGEMA_signal_15791), .Q (new_AGEMA_signal_15792) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7971 ( .C (clk), .D (new_AGEMA_signal_15795), .Q (new_AGEMA_signal_15796) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7975 ( .C (clk), .D (new_AGEMA_signal_15799), .Q (new_AGEMA_signal_15800) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7979 ( .C (clk), .D (new_AGEMA_signal_15803), .Q (new_AGEMA_signal_15804) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7983 ( .C (clk), .D (new_AGEMA_signal_15807), .Q (new_AGEMA_signal_15808) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7987 ( .C (clk), .D (new_AGEMA_signal_15811), .Q (new_AGEMA_signal_15812) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7991 ( .C (clk), .D (new_AGEMA_signal_15815), .Q (new_AGEMA_signal_15816) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7995 ( .C (clk), .D (new_AGEMA_signal_15819), .Q (new_AGEMA_signal_15820) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7999 ( .C (clk), .D (new_AGEMA_signal_15823), .Q (new_AGEMA_signal_15824) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8003 ( .C (clk), .D (new_AGEMA_signal_15827), .Q (new_AGEMA_signal_15828) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8007 ( .C (clk), .D (new_AGEMA_signal_15831), .Q (new_AGEMA_signal_15832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8011 ( .C (clk), .D (new_AGEMA_signal_15835), .Q (new_AGEMA_signal_15836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8015 ( .C (clk), .D (new_AGEMA_signal_15839), .Q (new_AGEMA_signal_15840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8019 ( .C (clk), .D (new_AGEMA_signal_15843), .Q (new_AGEMA_signal_15844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8023 ( .C (clk), .D (new_AGEMA_signal_15847), .Q (new_AGEMA_signal_15848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8027 ( .C (clk), .D (new_AGEMA_signal_15851), .Q (new_AGEMA_signal_15852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8031 ( .C (clk), .D (new_AGEMA_signal_15855), .Q (new_AGEMA_signal_15856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8035 ( .C (clk), .D (new_AGEMA_signal_15859), .Q (new_AGEMA_signal_15860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8039 ( .C (clk), .D (new_AGEMA_signal_15863), .Q (new_AGEMA_signal_15864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8043 ( .C (clk), .D (new_AGEMA_signal_15867), .Q (new_AGEMA_signal_15868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8047 ( .C (clk), .D (new_AGEMA_signal_15871), .Q (new_AGEMA_signal_15872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8051 ( .C (clk), .D (new_AGEMA_signal_15875), .Q (new_AGEMA_signal_15876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8055 ( .C (clk), .D (new_AGEMA_signal_15879), .Q (new_AGEMA_signal_15880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8059 ( .C (clk), .D (new_AGEMA_signal_15883), .Q (new_AGEMA_signal_15884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8063 ( .C (clk), .D (new_AGEMA_signal_15887), .Q (new_AGEMA_signal_15888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8067 ( .C (clk), .D (new_AGEMA_signal_15891), .Q (new_AGEMA_signal_15892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8071 ( .C (clk), .D (new_AGEMA_signal_15895), .Q (new_AGEMA_signal_15896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8075 ( .C (clk), .D (new_AGEMA_signal_15899), .Q (new_AGEMA_signal_15900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8079 ( .C (clk), .D (new_AGEMA_signal_15903), .Q (new_AGEMA_signal_15904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8083 ( .C (clk), .D (new_AGEMA_signal_15907), .Q (new_AGEMA_signal_15908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8087 ( .C (clk), .D (new_AGEMA_signal_15911), .Q (new_AGEMA_signal_15912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8091 ( .C (clk), .D (new_AGEMA_signal_15915), .Q (new_AGEMA_signal_15916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8095 ( .C (clk), .D (new_AGEMA_signal_15919), .Q (new_AGEMA_signal_15920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8099 ( .C (clk), .D (new_AGEMA_signal_15923), .Q (new_AGEMA_signal_15924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8103 ( .C (clk), .D (new_AGEMA_signal_15927), .Q (new_AGEMA_signal_15928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8107 ( .C (clk), .D (new_AGEMA_signal_15931), .Q (new_AGEMA_signal_15932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8111 ( .C (clk), .D (new_AGEMA_signal_15935), .Q (new_AGEMA_signal_15936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8115 ( .C (clk), .D (new_AGEMA_signal_15939), .Q (new_AGEMA_signal_15940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8119 ( .C (clk), .D (new_AGEMA_signal_15943), .Q (new_AGEMA_signal_15944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8123 ( .C (clk), .D (new_AGEMA_signal_15947), .Q (new_AGEMA_signal_15948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8127 ( .C (clk), .D (new_AGEMA_signal_15951), .Q (new_AGEMA_signal_15952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8131 ( .C (clk), .D (new_AGEMA_signal_15955), .Q (new_AGEMA_signal_15956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8135 ( .C (clk), .D (new_AGEMA_signal_15959), .Q (new_AGEMA_signal_15960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8139 ( .C (clk), .D (new_AGEMA_signal_15963), .Q (new_AGEMA_signal_15964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8143 ( .C (clk), .D (new_AGEMA_signal_15967), .Q (new_AGEMA_signal_15968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8147 ( .C (clk), .D (new_AGEMA_signal_15971), .Q (new_AGEMA_signal_15972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8151 ( .C (clk), .D (new_AGEMA_signal_15975), .Q (new_AGEMA_signal_15976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8155 ( .C (clk), .D (new_AGEMA_signal_15979), .Q (new_AGEMA_signal_15980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8159 ( .C (clk), .D (new_AGEMA_signal_15983), .Q (new_AGEMA_signal_15984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8163 ( .C (clk), .D (new_AGEMA_signal_15987), .Q (new_AGEMA_signal_15988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8167 ( .C (clk), .D (new_AGEMA_signal_15991), .Q (new_AGEMA_signal_15992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8171 ( .C (clk), .D (new_AGEMA_signal_15995), .Q (new_AGEMA_signal_15996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8175 ( .C (clk), .D (new_AGEMA_signal_15999), .Q (new_AGEMA_signal_16000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8179 ( .C (clk), .D (new_AGEMA_signal_16003), .Q (new_AGEMA_signal_16004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8183 ( .C (clk), .D (new_AGEMA_signal_16007), .Q (new_AGEMA_signal_16008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8187 ( .C (clk), .D (new_AGEMA_signal_16011), .Q (new_AGEMA_signal_16012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8191 ( .C (clk), .D (new_AGEMA_signal_16015), .Q (new_AGEMA_signal_16016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8195 ( .C (clk), .D (new_AGEMA_signal_16019), .Q (new_AGEMA_signal_16020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8199 ( .C (clk), .D (new_AGEMA_signal_16023), .Q (new_AGEMA_signal_16024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8203 ( .C (clk), .D (new_AGEMA_signal_16027), .Q (new_AGEMA_signal_16028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8207 ( .C (clk), .D (new_AGEMA_signal_16031), .Q (new_AGEMA_signal_16032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8211 ( .C (clk), .D (new_AGEMA_signal_16035), .Q (new_AGEMA_signal_16036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8215 ( .C (clk), .D (new_AGEMA_signal_16039), .Q (new_AGEMA_signal_16040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8219 ( .C (clk), .D (new_AGEMA_signal_16043), .Q (new_AGEMA_signal_16044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8223 ( .C (clk), .D (new_AGEMA_signal_16047), .Q (new_AGEMA_signal_16048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8227 ( .C (clk), .D (new_AGEMA_signal_16051), .Q (new_AGEMA_signal_16052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8231 ( .C (clk), .D (new_AGEMA_signal_16055), .Q (new_AGEMA_signal_16056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8235 ( .C (clk), .D (new_AGEMA_signal_16059), .Q (new_AGEMA_signal_16060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8239 ( .C (clk), .D (new_AGEMA_signal_16063), .Q (new_AGEMA_signal_16064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8243 ( .C (clk), .D (new_AGEMA_signal_16067), .Q (new_AGEMA_signal_16068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8247 ( .C (clk), .D (new_AGEMA_signal_16071), .Q (new_AGEMA_signal_16072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8251 ( .C (clk), .D (new_AGEMA_signal_16075), .Q (new_AGEMA_signal_16076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8255 ( .C (clk), .D (new_AGEMA_signal_16079), .Q (new_AGEMA_signal_16080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8259 ( .C (clk), .D (new_AGEMA_signal_16083), .Q (new_AGEMA_signal_16084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8263 ( .C (clk), .D (new_AGEMA_signal_16087), .Q (new_AGEMA_signal_16088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8267 ( .C (clk), .D (new_AGEMA_signal_16091), .Q (new_AGEMA_signal_16092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8271 ( .C (clk), .D (new_AGEMA_signal_16095), .Q (new_AGEMA_signal_16096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8275 ( .C (clk), .D (new_AGEMA_signal_16099), .Q (new_AGEMA_signal_16100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8279 ( .C (clk), .D (new_AGEMA_signal_16103), .Q (new_AGEMA_signal_16104) ) ;
    buf_clk new_AGEMA_reg_buffer_8283 ( .C (clk), .D (new_AGEMA_signal_16107), .Q (new_AGEMA_signal_16108) ) ;
    buf_clk new_AGEMA_reg_buffer_8287 ( .C (clk), .D (new_AGEMA_signal_16111), .Q (new_AGEMA_signal_16112) ) ;
    buf_clk new_AGEMA_reg_buffer_8291 ( .C (clk), .D (new_AGEMA_signal_16115), .Q (new_AGEMA_signal_16116) ) ;
    buf_clk new_AGEMA_reg_buffer_8295 ( .C (clk), .D (new_AGEMA_signal_16119), .Q (new_AGEMA_signal_16120) ) ;
    buf_clk new_AGEMA_reg_buffer_8299 ( .C (clk), .D (new_AGEMA_signal_16123), .Q (new_AGEMA_signal_16124) ) ;
    buf_clk new_AGEMA_reg_buffer_8303 ( .C (clk), .D (new_AGEMA_signal_16127), .Q (new_AGEMA_signal_16128) ) ;
    buf_clk new_AGEMA_reg_buffer_8307 ( .C (clk), .D (new_AGEMA_signal_16131), .Q (new_AGEMA_signal_16132) ) ;
    buf_clk new_AGEMA_reg_buffer_8311 ( .C (clk), .D (new_AGEMA_signal_16135), .Q (new_AGEMA_signal_16136) ) ;
    buf_clk new_AGEMA_reg_buffer_8315 ( .C (clk), .D (new_AGEMA_signal_16139), .Q (new_AGEMA_signal_16140) ) ;
    buf_clk new_AGEMA_reg_buffer_8319 ( .C (clk), .D (new_AGEMA_signal_16143), .Q (new_AGEMA_signal_16144) ) ;
    buf_clk new_AGEMA_reg_buffer_8323 ( .C (clk), .D (new_AGEMA_signal_16147), .Q (new_AGEMA_signal_16148) ) ;
    buf_clk new_AGEMA_reg_buffer_8327 ( .C (clk), .D (new_AGEMA_signal_16151), .Q (new_AGEMA_signal_16152) ) ;
    buf_clk new_AGEMA_reg_buffer_8331 ( .C (clk), .D (new_AGEMA_signal_16155), .Q (new_AGEMA_signal_16156) ) ;
    buf_clk new_AGEMA_reg_buffer_8335 ( .C (clk), .D (new_AGEMA_signal_16159), .Q (new_AGEMA_signal_16160) ) ;
    buf_clk new_AGEMA_reg_buffer_8339 ( .C (clk), .D (new_AGEMA_signal_16163), .Q (new_AGEMA_signal_16164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8343 ( .C (clk), .D (new_AGEMA_signal_16167), .Q (new_AGEMA_signal_16168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8347 ( .C (clk), .D (new_AGEMA_signal_16171), .Q (new_AGEMA_signal_16172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8351 ( .C (clk), .D (new_AGEMA_signal_16175), .Q (new_AGEMA_signal_16176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8355 ( .C (clk), .D (new_AGEMA_signal_16179), .Q (new_AGEMA_signal_16180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8359 ( .C (clk), .D (new_AGEMA_signal_16183), .Q (new_AGEMA_signal_16184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8363 ( .C (clk), .D (new_AGEMA_signal_16187), .Q (new_AGEMA_signal_16188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8367 ( .C (clk), .D (new_AGEMA_signal_16191), .Q (new_AGEMA_signal_16192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8371 ( .C (clk), .D (new_AGEMA_signal_16195), .Q (new_AGEMA_signal_16196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8375 ( .C (clk), .D (new_AGEMA_signal_16199), .Q (new_AGEMA_signal_16200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8379 ( .C (clk), .D (new_AGEMA_signal_16203), .Q (new_AGEMA_signal_16204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8383 ( .C (clk), .D (new_AGEMA_signal_16207), .Q (new_AGEMA_signal_16208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8387 ( .C (clk), .D (new_AGEMA_signal_16211), .Q (new_AGEMA_signal_16212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8391 ( .C (clk), .D (new_AGEMA_signal_16215), .Q (new_AGEMA_signal_16216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8395 ( .C (clk), .D (new_AGEMA_signal_16219), .Q (new_AGEMA_signal_16220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8399 ( .C (clk), .D (new_AGEMA_signal_16223), .Q (new_AGEMA_signal_16224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8403 ( .C (clk), .D (new_AGEMA_signal_16227), .Q (new_AGEMA_signal_16228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8407 ( .C (clk), .D (new_AGEMA_signal_16231), .Q (new_AGEMA_signal_16232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8411 ( .C (clk), .D (new_AGEMA_signal_16235), .Q (new_AGEMA_signal_16236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8415 ( .C (clk), .D (new_AGEMA_signal_16239), .Q (new_AGEMA_signal_16240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8419 ( .C (clk), .D (new_AGEMA_signal_16243), .Q (new_AGEMA_signal_16244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8423 ( .C (clk), .D (new_AGEMA_signal_16247), .Q (new_AGEMA_signal_16248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8427 ( .C (clk), .D (new_AGEMA_signal_16251), .Q (new_AGEMA_signal_16252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8431 ( .C (clk), .D (new_AGEMA_signal_16255), .Q (new_AGEMA_signal_16256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8435 ( .C (clk), .D (new_AGEMA_signal_16259), .Q (new_AGEMA_signal_16260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8439 ( .C (clk), .D (new_AGEMA_signal_16263), .Q (new_AGEMA_signal_16264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8443 ( .C (clk), .D (new_AGEMA_signal_16267), .Q (new_AGEMA_signal_16268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8447 ( .C (clk), .D (new_AGEMA_signal_16271), .Q (new_AGEMA_signal_16272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8451 ( .C (clk), .D (new_AGEMA_signal_16275), .Q (new_AGEMA_signal_16276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8455 ( .C (clk), .D (new_AGEMA_signal_16279), .Q (new_AGEMA_signal_16280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8459 ( .C (clk), .D (new_AGEMA_signal_16283), .Q (new_AGEMA_signal_16284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8463 ( .C (clk), .D (new_AGEMA_signal_16287), .Q (new_AGEMA_signal_16288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8467 ( .C (clk), .D (new_AGEMA_signal_16291), .Q (new_AGEMA_signal_16292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8471 ( .C (clk), .D (new_AGEMA_signal_16295), .Q (new_AGEMA_signal_16296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8475 ( .C (clk), .D (new_AGEMA_signal_16299), .Q (new_AGEMA_signal_16300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8479 ( .C (clk), .D (new_AGEMA_signal_16303), .Q (new_AGEMA_signal_16304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8483 ( .C (clk), .D (new_AGEMA_signal_16307), .Q (new_AGEMA_signal_16308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8487 ( .C (clk), .D (new_AGEMA_signal_16311), .Q (new_AGEMA_signal_16312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8491 ( .C (clk), .D (new_AGEMA_signal_16315), .Q (new_AGEMA_signal_16316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8495 ( .C (clk), .D (new_AGEMA_signal_16319), .Q (new_AGEMA_signal_16320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8499 ( .C (clk), .D (new_AGEMA_signal_16323), .Q (new_AGEMA_signal_16324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8503 ( .C (clk), .D (new_AGEMA_signal_16327), .Q (new_AGEMA_signal_16328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8507 ( .C (clk), .D (new_AGEMA_signal_16331), .Q (new_AGEMA_signal_16332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8511 ( .C (clk), .D (new_AGEMA_signal_16335), .Q (new_AGEMA_signal_16336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8515 ( .C (clk), .D (new_AGEMA_signal_16339), .Q (new_AGEMA_signal_16340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8519 ( .C (clk), .D (new_AGEMA_signal_16343), .Q (new_AGEMA_signal_16344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8523 ( .C (clk), .D (new_AGEMA_signal_16347), .Q (new_AGEMA_signal_16348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8527 ( .C (clk), .D (new_AGEMA_signal_16351), .Q (new_AGEMA_signal_16352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8531 ( .C (clk), .D (new_AGEMA_signal_16355), .Q (new_AGEMA_signal_16356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8535 ( .C (clk), .D (new_AGEMA_signal_16359), .Q (new_AGEMA_signal_16360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8539 ( .C (clk), .D (new_AGEMA_signal_16363), .Q (new_AGEMA_signal_16364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8543 ( .C (clk), .D (new_AGEMA_signal_16367), .Q (new_AGEMA_signal_16368) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8547 ( .C (clk), .D (new_AGEMA_signal_16371), .Q (new_AGEMA_signal_16372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8551 ( .C (clk), .D (new_AGEMA_signal_16375), .Q (new_AGEMA_signal_16376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8555 ( .C (clk), .D (new_AGEMA_signal_16379), .Q (new_AGEMA_signal_16380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8559 ( .C (clk), .D (new_AGEMA_signal_16383), .Q (new_AGEMA_signal_16384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8563 ( .C (clk), .D (new_AGEMA_signal_16387), .Q (new_AGEMA_signal_16388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8567 ( .C (clk), .D (new_AGEMA_signal_16391), .Q (new_AGEMA_signal_16392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8571 ( .C (clk), .D (new_AGEMA_signal_16395), .Q (new_AGEMA_signal_16396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8575 ( .C (clk), .D (new_AGEMA_signal_16399), .Q (new_AGEMA_signal_16400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8579 ( .C (clk), .D (new_AGEMA_signal_16403), .Q (new_AGEMA_signal_16404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8583 ( .C (clk), .D (new_AGEMA_signal_16407), .Q (new_AGEMA_signal_16408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8587 ( .C (clk), .D (new_AGEMA_signal_16411), .Q (new_AGEMA_signal_16412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8591 ( .C (clk), .D (new_AGEMA_signal_16415), .Q (new_AGEMA_signal_16416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8595 ( .C (clk), .D (new_AGEMA_signal_16419), .Q (new_AGEMA_signal_16420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8599 ( .C (clk), .D (new_AGEMA_signal_16423), .Q (new_AGEMA_signal_16424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8603 ( .C (clk), .D (new_AGEMA_signal_16427), .Q (new_AGEMA_signal_16428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8607 ( .C (clk), .D (new_AGEMA_signal_16431), .Q (new_AGEMA_signal_16432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8611 ( .C (clk), .D (new_AGEMA_signal_16435), .Q (new_AGEMA_signal_16436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8615 ( .C (clk), .D (new_AGEMA_signal_16439), .Q (new_AGEMA_signal_16440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8619 ( .C (clk), .D (new_AGEMA_signal_16443), .Q (new_AGEMA_signal_16444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8623 ( .C (clk), .D (new_AGEMA_signal_16447), .Q (new_AGEMA_signal_16448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8627 ( .C (clk), .D (new_AGEMA_signal_16451), .Q (new_AGEMA_signal_16452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8631 ( .C (clk), .D (new_AGEMA_signal_16455), .Q (new_AGEMA_signal_16456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8635 ( .C (clk), .D (new_AGEMA_signal_16459), .Q (new_AGEMA_signal_16460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8639 ( .C (clk), .D (new_AGEMA_signal_16463), .Q (new_AGEMA_signal_16464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8643 ( .C (clk), .D (new_AGEMA_signal_16467), .Q (new_AGEMA_signal_16468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8647 ( .C (clk), .D (new_AGEMA_signal_16471), .Q (new_AGEMA_signal_16472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8651 ( .C (clk), .D (new_AGEMA_signal_16475), .Q (new_AGEMA_signal_16476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8655 ( .C (clk), .D (new_AGEMA_signal_16479), .Q (new_AGEMA_signal_16480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8659 ( .C (clk), .D (new_AGEMA_signal_16483), .Q (new_AGEMA_signal_16484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8663 ( .C (clk), .D (new_AGEMA_signal_16487), .Q (new_AGEMA_signal_16488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8667 ( .C (clk), .D (new_AGEMA_signal_16491), .Q (new_AGEMA_signal_16492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8671 ( .C (clk), .D (new_AGEMA_signal_16495), .Q (new_AGEMA_signal_16496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8675 ( .C (clk), .D (new_AGEMA_signal_16499), .Q (new_AGEMA_signal_16500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8679 ( .C (clk), .D (new_AGEMA_signal_16503), .Q (new_AGEMA_signal_16504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8683 ( .C (clk), .D (new_AGEMA_signal_16507), .Q (new_AGEMA_signal_16508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8687 ( .C (clk), .D (new_AGEMA_signal_16511), .Q (new_AGEMA_signal_16512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8691 ( .C (clk), .D (new_AGEMA_signal_16515), .Q (new_AGEMA_signal_16516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8695 ( .C (clk), .D (new_AGEMA_signal_16519), .Q (new_AGEMA_signal_16520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8699 ( .C (clk), .D (new_AGEMA_signal_16523), .Q (new_AGEMA_signal_16524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8703 ( .C (clk), .D (new_AGEMA_signal_16527), .Q (new_AGEMA_signal_16528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8707 ( .C (clk), .D (new_AGEMA_signal_16531), .Q (new_AGEMA_signal_16532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8711 ( .C (clk), .D (new_AGEMA_signal_16535), .Q (new_AGEMA_signal_16536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8715 ( .C (clk), .D (new_AGEMA_signal_16539), .Q (new_AGEMA_signal_16540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8719 ( .C (clk), .D (new_AGEMA_signal_16543), .Q (new_AGEMA_signal_16544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8723 ( .C (clk), .D (new_AGEMA_signal_16547), .Q (new_AGEMA_signal_16548) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8727 ( .C (clk), .D (new_AGEMA_signal_16551), .Q (new_AGEMA_signal_16552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8731 ( .C (clk), .D (new_AGEMA_signal_16555), .Q (new_AGEMA_signal_16556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8735 ( .C (clk), .D (new_AGEMA_signal_16559), .Q (new_AGEMA_signal_16560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8739 ( .C (clk), .D (new_AGEMA_signal_16563), .Q (new_AGEMA_signal_16564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8743 ( .C (clk), .D (new_AGEMA_signal_16567), .Q (new_AGEMA_signal_16568) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8747 ( .C (clk), .D (new_AGEMA_signal_16571), .Q (new_AGEMA_signal_16572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8751 ( .C (clk), .D (new_AGEMA_signal_16575), .Q (new_AGEMA_signal_16576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8755 ( .C (clk), .D (new_AGEMA_signal_16579), .Q (new_AGEMA_signal_16580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8759 ( .C (clk), .D (new_AGEMA_signal_16583), .Q (new_AGEMA_signal_16584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8763 ( .C (clk), .D (new_AGEMA_signal_16587), .Q (new_AGEMA_signal_16588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8767 ( .C (clk), .D (new_AGEMA_signal_16591), .Q (new_AGEMA_signal_16592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8771 ( .C (clk), .D (new_AGEMA_signal_16595), .Q (new_AGEMA_signal_16596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8775 ( .C (clk), .D (new_AGEMA_signal_16599), .Q (new_AGEMA_signal_16600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8779 ( .C (clk), .D (new_AGEMA_signal_16603), .Q (new_AGEMA_signal_16604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8783 ( .C (clk), .D (new_AGEMA_signal_16607), .Q (new_AGEMA_signal_16608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8787 ( .C (clk), .D (new_AGEMA_signal_16611), .Q (new_AGEMA_signal_16612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8791 ( .C (clk), .D (new_AGEMA_signal_16615), .Q (new_AGEMA_signal_16616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8795 ( .C (clk), .D (new_AGEMA_signal_16619), .Q (new_AGEMA_signal_16620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8799 ( .C (clk), .D (new_AGEMA_signal_16623), .Q (new_AGEMA_signal_16624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8803 ( .C (clk), .D (new_AGEMA_signal_16627), .Q (new_AGEMA_signal_16628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8807 ( .C (clk), .D (new_AGEMA_signal_16631), .Q (new_AGEMA_signal_16632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8811 ( .C (clk), .D (new_AGEMA_signal_16635), .Q (new_AGEMA_signal_16636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8815 ( .C (clk), .D (new_AGEMA_signal_16639), .Q (new_AGEMA_signal_16640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8819 ( .C (clk), .D (new_AGEMA_signal_16643), .Q (new_AGEMA_signal_16644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8823 ( .C (clk), .D (new_AGEMA_signal_16647), .Q (new_AGEMA_signal_16648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8827 ( .C (clk), .D (new_AGEMA_signal_16651), .Q (new_AGEMA_signal_16652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8831 ( .C (clk), .D (new_AGEMA_signal_16655), .Q (new_AGEMA_signal_16656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8835 ( .C (clk), .D (new_AGEMA_signal_16659), .Q (new_AGEMA_signal_16660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8839 ( .C (clk), .D (new_AGEMA_signal_16663), .Q (new_AGEMA_signal_16664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8843 ( .C (clk), .D (new_AGEMA_signal_16667), .Q (new_AGEMA_signal_16668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8847 ( .C (clk), .D (new_AGEMA_signal_16671), .Q (new_AGEMA_signal_16672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8851 ( .C (clk), .D (new_AGEMA_signal_16675), .Q (new_AGEMA_signal_16676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8855 ( .C (clk), .D (new_AGEMA_signal_16679), .Q (new_AGEMA_signal_16680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8859 ( .C (clk), .D (new_AGEMA_signal_16683), .Q (new_AGEMA_signal_16684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8863 ( .C (clk), .D (new_AGEMA_signal_16687), .Q (new_AGEMA_signal_16688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8867 ( .C (clk), .D (new_AGEMA_signal_16691), .Q (new_AGEMA_signal_16692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8871 ( .C (clk), .D (new_AGEMA_signal_16695), .Q (new_AGEMA_signal_16696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8875 ( .C (clk), .D (new_AGEMA_signal_16699), .Q (new_AGEMA_signal_16700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8879 ( .C (clk), .D (new_AGEMA_signal_16703), .Q (new_AGEMA_signal_16704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8883 ( .C (clk), .D (new_AGEMA_signal_16707), .Q (new_AGEMA_signal_16708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8887 ( .C (clk), .D (new_AGEMA_signal_16711), .Q (new_AGEMA_signal_16712) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8891 ( .C (clk), .D (new_AGEMA_signal_16715), .Q (new_AGEMA_signal_16716) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8895 ( .C (clk), .D (new_AGEMA_signal_16719), .Q (new_AGEMA_signal_16720) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8899 ( .C (clk), .D (new_AGEMA_signal_16723), .Q (new_AGEMA_signal_16724) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8903 ( .C (clk), .D (new_AGEMA_signal_16727), .Q (new_AGEMA_signal_16728) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8907 ( .C (clk), .D (new_AGEMA_signal_16731), .Q (new_AGEMA_signal_16732) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8911 ( .C (clk), .D (new_AGEMA_signal_16735), .Q (new_AGEMA_signal_16736) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8915 ( .C (clk), .D (new_AGEMA_signal_16739), .Q (new_AGEMA_signal_16740) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8919 ( .C (clk), .D (new_AGEMA_signal_16743), .Q (new_AGEMA_signal_16744) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8923 ( .C (clk), .D (new_AGEMA_signal_16747), .Q (new_AGEMA_signal_16748) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8927 ( .C (clk), .D (new_AGEMA_signal_16751), .Q (new_AGEMA_signal_16752) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8931 ( .C (clk), .D (new_AGEMA_signal_16755), .Q (new_AGEMA_signal_16756) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8935 ( .C (clk), .D (new_AGEMA_signal_16759), .Q (new_AGEMA_signal_16760) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8939 ( .C (clk), .D (new_AGEMA_signal_16763), .Q (new_AGEMA_signal_16764) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8943 ( .C (clk), .D (new_AGEMA_signal_16767), .Q (new_AGEMA_signal_16768) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8947 ( .C (clk), .D (new_AGEMA_signal_16771), .Q (new_AGEMA_signal_16772) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8951 ( .C (clk), .D (new_AGEMA_signal_16775), .Q (new_AGEMA_signal_16776) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8955 ( .C (clk), .D (new_AGEMA_signal_16779), .Q (new_AGEMA_signal_16780) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8959 ( .C (clk), .D (new_AGEMA_signal_16783), .Q (new_AGEMA_signal_16784) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8963 ( .C (clk), .D (new_AGEMA_signal_16787), .Q (new_AGEMA_signal_16788) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8967 ( .C (clk), .D (new_AGEMA_signal_16791), .Q (new_AGEMA_signal_16792) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8971 ( .C (clk), .D (new_AGEMA_signal_16795), .Q (new_AGEMA_signal_16796) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8975 ( .C (clk), .D (new_AGEMA_signal_16799), .Q (new_AGEMA_signal_16800) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8979 ( .C (clk), .D (new_AGEMA_signal_16803), .Q (new_AGEMA_signal_16804) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8983 ( .C (clk), .D (new_AGEMA_signal_16807), .Q (new_AGEMA_signal_16808) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8987 ( .C (clk), .D (new_AGEMA_signal_16811), .Q (new_AGEMA_signal_16812) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8991 ( .C (clk), .D (new_AGEMA_signal_16815), .Q (new_AGEMA_signal_16816) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8995 ( .C (clk), .D (new_AGEMA_signal_16819), .Q (new_AGEMA_signal_16820) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8999 ( .C (clk), .D (new_AGEMA_signal_16823), .Q (new_AGEMA_signal_16824) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9003 ( .C (clk), .D (new_AGEMA_signal_16827), .Q (new_AGEMA_signal_16828) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9007 ( .C (clk), .D (new_AGEMA_signal_16831), .Q (new_AGEMA_signal_16832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9011 ( .C (clk), .D (new_AGEMA_signal_16835), .Q (new_AGEMA_signal_16836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9015 ( .C (clk), .D (new_AGEMA_signal_16839), .Q (new_AGEMA_signal_16840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9019 ( .C (clk), .D (new_AGEMA_signal_16843), .Q (new_AGEMA_signal_16844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9023 ( .C (clk), .D (new_AGEMA_signal_16847), .Q (new_AGEMA_signal_16848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9027 ( .C (clk), .D (new_AGEMA_signal_16851), .Q (new_AGEMA_signal_16852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9031 ( .C (clk), .D (new_AGEMA_signal_16855), .Q (new_AGEMA_signal_16856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9035 ( .C (clk), .D (new_AGEMA_signal_16859), .Q (new_AGEMA_signal_16860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9039 ( .C (clk), .D (new_AGEMA_signal_16863), .Q (new_AGEMA_signal_16864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9043 ( .C (clk), .D (new_AGEMA_signal_16867), .Q (new_AGEMA_signal_16868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9047 ( .C (clk), .D (new_AGEMA_signal_16871), .Q (new_AGEMA_signal_16872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9051 ( .C (clk), .D (new_AGEMA_signal_16875), .Q (new_AGEMA_signal_16876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9055 ( .C (clk), .D (new_AGEMA_signal_16879), .Q (new_AGEMA_signal_16880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9059 ( .C (clk), .D (new_AGEMA_signal_16883), .Q (new_AGEMA_signal_16884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9063 ( .C (clk), .D (new_AGEMA_signal_16887), .Q (new_AGEMA_signal_16888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9067 ( .C (clk), .D (new_AGEMA_signal_16891), .Q (new_AGEMA_signal_16892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9071 ( .C (clk), .D (new_AGEMA_signal_16895), .Q (new_AGEMA_signal_16896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9075 ( .C (clk), .D (new_AGEMA_signal_16899), .Q (new_AGEMA_signal_16900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9079 ( .C (clk), .D (new_AGEMA_signal_16903), .Q (new_AGEMA_signal_16904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9083 ( .C (clk), .D (new_AGEMA_signal_16907), .Q (new_AGEMA_signal_16908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9087 ( .C (clk), .D (new_AGEMA_signal_16911), .Q (new_AGEMA_signal_16912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9091 ( .C (clk), .D (new_AGEMA_signal_16915), .Q (new_AGEMA_signal_16916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9095 ( .C (clk), .D (new_AGEMA_signal_16919), .Q (new_AGEMA_signal_16920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9099 ( .C (clk), .D (new_AGEMA_signal_16923), .Q (new_AGEMA_signal_16924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9103 ( .C (clk), .D (new_AGEMA_signal_16927), .Q (new_AGEMA_signal_16928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9107 ( .C (clk), .D (new_AGEMA_signal_16931), .Q (new_AGEMA_signal_16932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9111 ( .C (clk), .D (new_AGEMA_signal_16935), .Q (new_AGEMA_signal_16936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9115 ( .C (clk), .D (new_AGEMA_signal_16939), .Q (new_AGEMA_signal_16940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9119 ( .C (clk), .D (new_AGEMA_signal_16943), .Q (new_AGEMA_signal_16944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9123 ( .C (clk), .D (new_AGEMA_signal_16947), .Q (new_AGEMA_signal_16948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9127 ( .C (clk), .D (new_AGEMA_signal_16951), .Q (new_AGEMA_signal_16952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9131 ( .C (clk), .D (new_AGEMA_signal_16955), .Q (new_AGEMA_signal_16956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9135 ( .C (clk), .D (new_AGEMA_signal_16959), .Q (new_AGEMA_signal_16960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9139 ( .C (clk), .D (new_AGEMA_signal_16963), .Q (new_AGEMA_signal_16964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9143 ( .C (clk), .D (new_AGEMA_signal_16967), .Q (new_AGEMA_signal_16968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9147 ( .C (clk), .D (new_AGEMA_signal_16971), .Q (new_AGEMA_signal_16972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9151 ( .C (clk), .D (new_AGEMA_signal_16975), .Q (new_AGEMA_signal_16976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9155 ( .C (clk), .D (new_AGEMA_signal_16979), .Q (new_AGEMA_signal_16980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9159 ( .C (clk), .D (new_AGEMA_signal_16983), .Q (new_AGEMA_signal_16984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9163 ( .C (clk), .D (new_AGEMA_signal_16987), .Q (new_AGEMA_signal_16988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9167 ( .C (clk), .D (new_AGEMA_signal_16991), .Q (new_AGEMA_signal_16992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9171 ( .C (clk), .D (new_AGEMA_signal_16995), .Q (new_AGEMA_signal_16996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9175 ( .C (clk), .D (new_AGEMA_signal_16999), .Q (new_AGEMA_signal_17000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9179 ( .C (clk), .D (new_AGEMA_signal_17003), .Q (new_AGEMA_signal_17004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9183 ( .C (clk), .D (new_AGEMA_signal_17007), .Q (new_AGEMA_signal_17008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9187 ( .C (clk), .D (new_AGEMA_signal_17011), .Q (new_AGEMA_signal_17012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9191 ( .C (clk), .D (new_AGEMA_signal_17015), .Q (new_AGEMA_signal_17016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9195 ( .C (clk), .D (new_AGEMA_signal_17019), .Q (new_AGEMA_signal_17020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9199 ( .C (clk), .D (new_AGEMA_signal_17023), .Q (new_AGEMA_signal_17024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9203 ( .C (clk), .D (new_AGEMA_signal_17027), .Q (new_AGEMA_signal_17028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9207 ( .C (clk), .D (new_AGEMA_signal_17031), .Q (new_AGEMA_signal_17032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9211 ( .C (clk), .D (new_AGEMA_signal_17035), .Q (new_AGEMA_signal_17036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9215 ( .C (clk), .D (new_AGEMA_signal_17039), .Q (new_AGEMA_signal_17040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9219 ( .C (clk), .D (new_AGEMA_signal_17043), .Q (new_AGEMA_signal_17044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9223 ( .C (clk), .D (new_AGEMA_signal_17047), .Q (new_AGEMA_signal_17048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9227 ( .C (clk), .D (new_AGEMA_signal_17051), .Q (new_AGEMA_signal_17052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9231 ( .C (clk), .D (new_AGEMA_signal_17055), .Q (new_AGEMA_signal_17056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9235 ( .C (clk), .D (new_AGEMA_signal_17059), .Q (new_AGEMA_signal_17060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9239 ( .C (clk), .D (new_AGEMA_signal_17063), .Q (new_AGEMA_signal_17064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9243 ( .C (clk), .D (new_AGEMA_signal_17067), .Q (new_AGEMA_signal_17068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9247 ( .C (clk), .D (new_AGEMA_signal_17071), .Q (new_AGEMA_signal_17072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9251 ( .C (clk), .D (new_AGEMA_signal_17075), .Q (new_AGEMA_signal_17076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9255 ( .C (clk), .D (new_AGEMA_signal_17079), .Q (new_AGEMA_signal_17080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9259 ( .C (clk), .D (new_AGEMA_signal_17083), .Q (new_AGEMA_signal_17084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9263 ( .C (clk), .D (new_AGEMA_signal_17087), .Q (new_AGEMA_signal_17088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9267 ( .C (clk), .D (new_AGEMA_signal_17091), .Q (new_AGEMA_signal_17092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9271 ( .C (clk), .D (new_AGEMA_signal_17095), .Q (new_AGEMA_signal_17096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9275 ( .C (clk), .D (new_AGEMA_signal_17099), .Q (new_AGEMA_signal_17100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9279 ( .C (clk), .D (new_AGEMA_signal_17103), .Q (new_AGEMA_signal_17104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9283 ( .C (clk), .D (new_AGEMA_signal_17107), .Q (new_AGEMA_signal_17108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9287 ( .C (clk), .D (new_AGEMA_signal_17111), .Q (new_AGEMA_signal_17112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9291 ( .C (clk), .D (new_AGEMA_signal_17115), .Q (new_AGEMA_signal_17116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9295 ( .C (clk), .D (new_AGEMA_signal_17119), .Q (new_AGEMA_signal_17120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9299 ( .C (clk), .D (new_AGEMA_signal_17123), .Q (new_AGEMA_signal_17124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9303 ( .C (clk), .D (new_AGEMA_signal_17127), .Q (new_AGEMA_signal_17128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9307 ( .C (clk), .D (new_AGEMA_signal_17131), .Q (new_AGEMA_signal_17132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9311 ( .C (clk), .D (new_AGEMA_signal_17135), .Q (new_AGEMA_signal_17136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9315 ( .C (clk), .D (new_AGEMA_signal_17139), .Q (new_AGEMA_signal_17140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9319 ( .C (clk), .D (new_AGEMA_signal_17143), .Q (new_AGEMA_signal_17144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9323 ( .C (clk), .D (new_AGEMA_signal_17147), .Q (new_AGEMA_signal_17148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9327 ( .C (clk), .D (new_AGEMA_signal_17151), .Q (new_AGEMA_signal_17152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9331 ( .C (clk), .D (new_AGEMA_signal_17155), .Q (new_AGEMA_signal_17156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9335 ( .C (clk), .D (new_AGEMA_signal_17159), .Q (new_AGEMA_signal_17160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9339 ( .C (clk), .D (new_AGEMA_signal_17163), .Q (new_AGEMA_signal_17164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9343 ( .C (clk), .D (new_AGEMA_signal_17167), .Q (new_AGEMA_signal_17168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9347 ( .C (clk), .D (new_AGEMA_signal_17171), .Q (new_AGEMA_signal_17172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9351 ( .C (clk), .D (new_AGEMA_signal_17175), .Q (new_AGEMA_signal_17176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9355 ( .C (clk), .D (new_AGEMA_signal_17179), .Q (new_AGEMA_signal_17180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9359 ( .C (clk), .D (new_AGEMA_signal_17183), .Q (new_AGEMA_signal_17184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9363 ( .C (clk), .D (new_AGEMA_signal_17187), .Q (new_AGEMA_signal_17188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9367 ( .C (clk), .D (new_AGEMA_signal_17191), .Q (new_AGEMA_signal_17192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9371 ( .C (clk), .D (new_AGEMA_signal_17195), .Q (new_AGEMA_signal_17196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9375 ( .C (clk), .D (new_AGEMA_signal_17199), .Q (new_AGEMA_signal_17200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9379 ( .C (clk), .D (new_AGEMA_signal_17203), .Q (new_AGEMA_signal_17204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9383 ( .C (clk), .D (new_AGEMA_signal_17207), .Q (new_AGEMA_signal_17208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9387 ( .C (clk), .D (new_AGEMA_signal_17211), .Q (new_AGEMA_signal_17212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9391 ( .C (clk), .D (new_AGEMA_signal_17215), .Q (new_AGEMA_signal_17216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9395 ( .C (clk), .D (new_AGEMA_signal_17219), .Q (new_AGEMA_signal_17220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9399 ( .C (clk), .D (new_AGEMA_signal_17223), .Q (new_AGEMA_signal_17224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9403 ( .C (clk), .D (new_AGEMA_signal_17227), .Q (new_AGEMA_signal_17228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9407 ( .C (clk), .D (new_AGEMA_signal_17231), .Q (new_AGEMA_signal_17232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9411 ( .C (clk), .D (new_AGEMA_signal_17235), .Q (new_AGEMA_signal_17236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9415 ( .C (clk), .D (new_AGEMA_signal_17239), .Q (new_AGEMA_signal_17240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9419 ( .C (clk), .D (new_AGEMA_signal_17243), .Q (new_AGEMA_signal_17244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9423 ( .C (clk), .D (new_AGEMA_signal_17247), .Q (new_AGEMA_signal_17248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9427 ( .C (clk), .D (new_AGEMA_signal_17251), .Q (new_AGEMA_signal_17252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9431 ( .C (clk), .D (new_AGEMA_signal_17255), .Q (new_AGEMA_signal_17256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9435 ( .C (clk), .D (new_AGEMA_signal_17259), .Q (new_AGEMA_signal_17260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9439 ( .C (clk), .D (new_AGEMA_signal_17263), .Q (new_AGEMA_signal_17264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9443 ( .C (clk), .D (new_AGEMA_signal_17267), .Q (new_AGEMA_signal_17268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9447 ( .C (clk), .D (new_AGEMA_signal_17271), .Q (new_AGEMA_signal_17272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9451 ( .C (clk), .D (new_AGEMA_signal_17275), .Q (new_AGEMA_signal_17276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9455 ( .C (clk), .D (new_AGEMA_signal_17279), .Q (new_AGEMA_signal_17280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9459 ( .C (clk), .D (new_AGEMA_signal_17283), .Q (new_AGEMA_signal_17284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9463 ( .C (clk), .D (new_AGEMA_signal_17287), .Q (new_AGEMA_signal_17288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9467 ( .C (clk), .D (new_AGEMA_signal_17291), .Q (new_AGEMA_signal_17292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9471 ( .C (clk), .D (new_AGEMA_signal_17295), .Q (new_AGEMA_signal_17296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9475 ( .C (clk), .D (new_AGEMA_signal_17299), .Q (new_AGEMA_signal_17300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9479 ( .C (clk), .D (new_AGEMA_signal_17303), .Q (new_AGEMA_signal_17304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9483 ( .C (clk), .D (new_AGEMA_signal_17307), .Q (new_AGEMA_signal_17308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9487 ( .C (clk), .D (new_AGEMA_signal_17311), .Q (new_AGEMA_signal_17312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9491 ( .C (clk), .D (new_AGEMA_signal_17315), .Q (new_AGEMA_signal_17316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9495 ( .C (clk), .D (new_AGEMA_signal_17319), .Q (new_AGEMA_signal_17320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9499 ( .C (clk), .D (new_AGEMA_signal_17323), .Q (new_AGEMA_signal_17324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9503 ( .C (clk), .D (new_AGEMA_signal_17327), .Q (new_AGEMA_signal_17328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9507 ( .C (clk), .D (new_AGEMA_signal_17331), .Q (new_AGEMA_signal_17332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9511 ( .C (clk), .D (new_AGEMA_signal_17335), .Q (new_AGEMA_signal_17336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9515 ( .C (clk), .D (new_AGEMA_signal_17339), .Q (new_AGEMA_signal_17340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9519 ( .C (clk), .D (new_AGEMA_signal_17343), .Q (new_AGEMA_signal_17344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9523 ( .C (clk), .D (new_AGEMA_signal_17347), .Q (new_AGEMA_signal_17348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9527 ( .C (clk), .D (new_AGEMA_signal_17351), .Q (new_AGEMA_signal_17352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9531 ( .C (clk), .D (new_AGEMA_signal_17355), .Q (new_AGEMA_signal_17356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9535 ( .C (clk), .D (new_AGEMA_signal_17359), .Q (new_AGEMA_signal_17360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9539 ( .C (clk), .D (new_AGEMA_signal_17363), .Q (new_AGEMA_signal_17364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9543 ( .C (clk), .D (new_AGEMA_signal_17367), .Q (new_AGEMA_signal_17368) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9547 ( .C (clk), .D (new_AGEMA_signal_17371), .Q (new_AGEMA_signal_17372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9551 ( .C (clk), .D (new_AGEMA_signal_17375), .Q (new_AGEMA_signal_17376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9555 ( .C (clk), .D (new_AGEMA_signal_17379), .Q (new_AGEMA_signal_17380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9559 ( .C (clk), .D (new_AGEMA_signal_17383), .Q (new_AGEMA_signal_17384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9563 ( .C (clk), .D (new_AGEMA_signal_17387), .Q (new_AGEMA_signal_17388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9567 ( .C (clk), .D (new_AGEMA_signal_17391), .Q (new_AGEMA_signal_17392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9571 ( .C (clk), .D (new_AGEMA_signal_17395), .Q (new_AGEMA_signal_17396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9575 ( .C (clk), .D (new_AGEMA_signal_17399), .Q (new_AGEMA_signal_17400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9579 ( .C (clk), .D (new_AGEMA_signal_17403), .Q (new_AGEMA_signal_17404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9583 ( .C (clk), .D (new_AGEMA_signal_17407), .Q (new_AGEMA_signal_17408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9587 ( .C (clk), .D (new_AGEMA_signal_17411), .Q (new_AGEMA_signal_17412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9591 ( .C (clk), .D (new_AGEMA_signal_17415), .Q (new_AGEMA_signal_17416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9595 ( .C (clk), .D (new_AGEMA_signal_17419), .Q (new_AGEMA_signal_17420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9599 ( .C (clk), .D (new_AGEMA_signal_17423), .Q (new_AGEMA_signal_17424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9603 ( .C (clk), .D (new_AGEMA_signal_17427), .Q (new_AGEMA_signal_17428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9607 ( .C (clk), .D (new_AGEMA_signal_17431), .Q (new_AGEMA_signal_17432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9611 ( .C (clk), .D (new_AGEMA_signal_17435), .Q (new_AGEMA_signal_17436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9615 ( .C (clk), .D (new_AGEMA_signal_17439), .Q (new_AGEMA_signal_17440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9619 ( .C (clk), .D (new_AGEMA_signal_17443), .Q (new_AGEMA_signal_17444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9623 ( .C (clk), .D (new_AGEMA_signal_17447), .Q (new_AGEMA_signal_17448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9627 ( .C (clk), .D (new_AGEMA_signal_17451), .Q (new_AGEMA_signal_17452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9631 ( .C (clk), .D (new_AGEMA_signal_17455), .Q (new_AGEMA_signal_17456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9635 ( .C (clk), .D (new_AGEMA_signal_17459), .Q (new_AGEMA_signal_17460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9639 ( .C (clk), .D (new_AGEMA_signal_17463), .Q (new_AGEMA_signal_17464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9643 ( .C (clk), .D (new_AGEMA_signal_17467), .Q (new_AGEMA_signal_17468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9647 ( .C (clk), .D (new_AGEMA_signal_17471), .Q (new_AGEMA_signal_17472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9651 ( .C (clk), .D (new_AGEMA_signal_17475), .Q (new_AGEMA_signal_17476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9655 ( .C (clk), .D (new_AGEMA_signal_17479), .Q (new_AGEMA_signal_17480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9659 ( .C (clk), .D (new_AGEMA_signal_17483), .Q (new_AGEMA_signal_17484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9663 ( .C (clk), .D (new_AGEMA_signal_17487), .Q (new_AGEMA_signal_17488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9667 ( .C (clk), .D (new_AGEMA_signal_17491), .Q (new_AGEMA_signal_17492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9671 ( .C (clk), .D (new_AGEMA_signal_17495), .Q (new_AGEMA_signal_17496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9675 ( .C (clk), .D (new_AGEMA_signal_17499), .Q (new_AGEMA_signal_17500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9679 ( .C (clk), .D (new_AGEMA_signal_17503), .Q (new_AGEMA_signal_17504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9683 ( .C (clk), .D (new_AGEMA_signal_17507), .Q (new_AGEMA_signal_17508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9687 ( .C (clk), .D (new_AGEMA_signal_17511), .Q (new_AGEMA_signal_17512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9691 ( .C (clk), .D (new_AGEMA_signal_17515), .Q (new_AGEMA_signal_17516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9695 ( .C (clk), .D (new_AGEMA_signal_17519), .Q (new_AGEMA_signal_17520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9699 ( .C (clk), .D (new_AGEMA_signal_17523), .Q (new_AGEMA_signal_17524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9703 ( .C (clk), .D (new_AGEMA_signal_17527), .Q (new_AGEMA_signal_17528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9707 ( .C (clk), .D (new_AGEMA_signal_17531), .Q (new_AGEMA_signal_17532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9711 ( .C (clk), .D (new_AGEMA_signal_17535), .Q (new_AGEMA_signal_17536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9715 ( .C (clk), .D (new_AGEMA_signal_17539), .Q (new_AGEMA_signal_17540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9719 ( .C (clk), .D (new_AGEMA_signal_17543), .Q (new_AGEMA_signal_17544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9723 ( .C (clk), .D (new_AGEMA_signal_17547), .Q (new_AGEMA_signal_17548) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9727 ( .C (clk), .D (new_AGEMA_signal_17551), .Q (new_AGEMA_signal_17552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9731 ( .C (clk), .D (new_AGEMA_signal_17555), .Q (new_AGEMA_signal_17556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9735 ( .C (clk), .D (new_AGEMA_signal_17559), .Q (new_AGEMA_signal_17560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9739 ( .C (clk), .D (new_AGEMA_signal_17563), .Q (new_AGEMA_signal_17564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9743 ( .C (clk), .D (new_AGEMA_signal_17567), .Q (new_AGEMA_signal_17568) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9747 ( .C (clk), .D (new_AGEMA_signal_17571), .Q (new_AGEMA_signal_17572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9751 ( .C (clk), .D (new_AGEMA_signal_17575), .Q (new_AGEMA_signal_17576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9755 ( .C (clk), .D (new_AGEMA_signal_17579), .Q (new_AGEMA_signal_17580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9759 ( .C (clk), .D (new_AGEMA_signal_17583), .Q (new_AGEMA_signal_17584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9763 ( .C (clk), .D (new_AGEMA_signal_17587), .Q (new_AGEMA_signal_17588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9767 ( .C (clk), .D (new_AGEMA_signal_17591), .Q (new_AGEMA_signal_17592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9771 ( .C (clk), .D (new_AGEMA_signal_17595), .Q (new_AGEMA_signal_17596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9775 ( .C (clk), .D (new_AGEMA_signal_17599), .Q (new_AGEMA_signal_17600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9779 ( .C (clk), .D (new_AGEMA_signal_17603), .Q (new_AGEMA_signal_17604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9783 ( .C (clk), .D (new_AGEMA_signal_17607), .Q (new_AGEMA_signal_17608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9787 ( .C (clk), .D (new_AGEMA_signal_17611), .Q (new_AGEMA_signal_17612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9791 ( .C (clk), .D (new_AGEMA_signal_17615), .Q (new_AGEMA_signal_17616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9795 ( .C (clk), .D (new_AGEMA_signal_17619), .Q (new_AGEMA_signal_17620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9799 ( .C (clk), .D (new_AGEMA_signal_17623), .Q (new_AGEMA_signal_17624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9803 ( .C (clk), .D (new_AGEMA_signal_17627), .Q (new_AGEMA_signal_17628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9807 ( .C (clk), .D (new_AGEMA_signal_17631), .Q (new_AGEMA_signal_17632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9811 ( .C (clk), .D (new_AGEMA_signal_17635), .Q (new_AGEMA_signal_17636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9815 ( .C (clk), .D (new_AGEMA_signal_17639), .Q (new_AGEMA_signal_17640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9819 ( .C (clk), .D (new_AGEMA_signal_17643), .Q (new_AGEMA_signal_17644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9823 ( .C (clk), .D (new_AGEMA_signal_17647), .Q (new_AGEMA_signal_17648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9827 ( .C (clk), .D (new_AGEMA_signal_17651), .Q (new_AGEMA_signal_17652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9831 ( .C (clk), .D (new_AGEMA_signal_17655), .Q (new_AGEMA_signal_17656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9835 ( .C (clk), .D (new_AGEMA_signal_17659), .Q (new_AGEMA_signal_17660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9839 ( .C (clk), .D (new_AGEMA_signal_17663), .Q (new_AGEMA_signal_17664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9843 ( .C (clk), .D (new_AGEMA_signal_17667), .Q (new_AGEMA_signal_17668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9847 ( .C (clk), .D (new_AGEMA_signal_17671), .Q (new_AGEMA_signal_17672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9851 ( .C (clk), .D (new_AGEMA_signal_17675), .Q (new_AGEMA_signal_17676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9855 ( .C (clk), .D (new_AGEMA_signal_17679), .Q (new_AGEMA_signal_17680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9859 ( .C (clk), .D (new_AGEMA_signal_17683), .Q (new_AGEMA_signal_17684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9863 ( .C (clk), .D (new_AGEMA_signal_17687), .Q (new_AGEMA_signal_17688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9867 ( .C (clk), .D (new_AGEMA_signal_17691), .Q (new_AGEMA_signal_17692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9871 ( .C (clk), .D (new_AGEMA_signal_17695), .Q (new_AGEMA_signal_17696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9875 ( .C (clk), .D (new_AGEMA_signal_17699), .Q (new_AGEMA_signal_17700) ) ;
    buf_clk new_AGEMA_reg_buffer_9879 ( .C (clk), .D (new_AGEMA_signal_17703), .Q (new_AGEMA_signal_17704) ) ;
    buf_clk new_AGEMA_reg_buffer_9883 ( .C (clk), .D (new_AGEMA_signal_17707), .Q (new_AGEMA_signal_17708) ) ;
    buf_clk new_AGEMA_reg_buffer_9887 ( .C (clk), .D (new_AGEMA_signal_17711), .Q (new_AGEMA_signal_17712) ) ;
    buf_clk new_AGEMA_reg_buffer_9891 ( .C (clk), .D (new_AGEMA_signal_17715), .Q (new_AGEMA_signal_17716) ) ;
    buf_clk new_AGEMA_reg_buffer_9895 ( .C (clk), .D (new_AGEMA_signal_17719), .Q (new_AGEMA_signal_17720) ) ;
    buf_clk new_AGEMA_reg_buffer_9899 ( .C (clk), .D (new_AGEMA_signal_17723), .Q (new_AGEMA_signal_17724) ) ;
    buf_clk new_AGEMA_reg_buffer_9903 ( .C (clk), .D (new_AGEMA_signal_17727), .Q (new_AGEMA_signal_17728) ) ;

    /* cells in depth 4 */
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7431, new_AGEMA_signal_7430, new_AGEMA_signal_7429, RoundOutput[0]}), .a ({new_AGEMA_signal_10097, new_AGEMA_signal_10093, new_AGEMA_signal_10089, new_AGEMA_signal_10085}), .c ({new_AGEMA_signal_7794, new_AGEMA_signal_7793, new_AGEMA_signal_7792, RoundReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7911, new_AGEMA_signal_7910, new_AGEMA_signal_7909, RoundOutput[1]}), .a ({new_AGEMA_signal_10113, new_AGEMA_signal_10109, new_AGEMA_signal_10105, new_AGEMA_signal_10101}), .c ({new_AGEMA_signal_8145, new_AGEMA_signal_8144, new_AGEMA_signal_8143, RoundReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7434, new_AGEMA_signal_7433, new_AGEMA_signal_7432, RoundOutput[2]}), .a ({new_AGEMA_signal_10129, new_AGEMA_signal_10125, new_AGEMA_signal_10121, new_AGEMA_signal_10117}), .c ({new_AGEMA_signal_7800, new_AGEMA_signal_7799, new_AGEMA_signal_7798, RoundReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7914, new_AGEMA_signal_7913, new_AGEMA_signal_7912, RoundOutput[3]}), .a ({new_AGEMA_signal_10145, new_AGEMA_signal_10141, new_AGEMA_signal_10137, new_AGEMA_signal_10133}), .c ({new_AGEMA_signal_8151, new_AGEMA_signal_8150, new_AGEMA_signal_8149, RoundReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7917, new_AGEMA_signal_7916, new_AGEMA_signal_7915, RoundOutput[4]}), .a ({new_AGEMA_signal_10161, new_AGEMA_signal_10157, new_AGEMA_signal_10153, new_AGEMA_signal_10149}), .c ({new_AGEMA_signal_8157, new_AGEMA_signal_8156, new_AGEMA_signal_8155, RoundReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7437, new_AGEMA_signal_7436, new_AGEMA_signal_7435, RoundOutput[5]}), .a ({new_AGEMA_signal_10177, new_AGEMA_signal_10173, new_AGEMA_signal_10169, new_AGEMA_signal_10165}), .c ({new_AGEMA_signal_7806, new_AGEMA_signal_7805, new_AGEMA_signal_7804, RoundReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7440, new_AGEMA_signal_7439, new_AGEMA_signal_7438, RoundOutput[6]}), .a ({new_AGEMA_signal_10193, new_AGEMA_signal_10189, new_AGEMA_signal_10185, new_AGEMA_signal_10181}), .c ({new_AGEMA_signal_7812, new_AGEMA_signal_7811, new_AGEMA_signal_7810, RoundReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7443, new_AGEMA_signal_7442, new_AGEMA_signal_7441, RoundOutput[7]}), .a ({new_AGEMA_signal_10209, new_AGEMA_signal_10205, new_AGEMA_signal_10201, new_AGEMA_signal_10197}), .c ({new_AGEMA_signal_7818, new_AGEMA_signal_7817, new_AGEMA_signal_7816, RoundReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7446, new_AGEMA_signal_7445, new_AGEMA_signal_7444, RoundOutput[8]}), .a ({new_AGEMA_signal_10225, new_AGEMA_signal_10221, new_AGEMA_signal_10217, new_AGEMA_signal_10213}), .c ({new_AGEMA_signal_7824, new_AGEMA_signal_7823, new_AGEMA_signal_7822, RoundReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7920, new_AGEMA_signal_7919, new_AGEMA_signal_7918, RoundOutput[9]}), .a ({new_AGEMA_signal_10241, new_AGEMA_signal_10237, new_AGEMA_signal_10233, new_AGEMA_signal_10229}), .c ({new_AGEMA_signal_8163, new_AGEMA_signal_8162, new_AGEMA_signal_8161, RoundReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7449, new_AGEMA_signal_7448, new_AGEMA_signal_7447, RoundOutput[10]}), .a ({new_AGEMA_signal_10257, new_AGEMA_signal_10253, new_AGEMA_signal_10249, new_AGEMA_signal_10245}), .c ({new_AGEMA_signal_7830, new_AGEMA_signal_7829, new_AGEMA_signal_7828, RoundReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7923, new_AGEMA_signal_7922, new_AGEMA_signal_7921, RoundOutput[11]}), .a ({new_AGEMA_signal_10273, new_AGEMA_signal_10269, new_AGEMA_signal_10265, new_AGEMA_signal_10261}), .c ({new_AGEMA_signal_8169, new_AGEMA_signal_8168, new_AGEMA_signal_8167, RoundReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7926, new_AGEMA_signal_7925, new_AGEMA_signal_7924, RoundOutput[12]}), .a ({new_AGEMA_signal_10289, new_AGEMA_signal_10285, new_AGEMA_signal_10281, new_AGEMA_signal_10277}), .c ({new_AGEMA_signal_8175, new_AGEMA_signal_8174, new_AGEMA_signal_8173, RoundReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7452, new_AGEMA_signal_7451, new_AGEMA_signal_7450, RoundOutput[13]}), .a ({new_AGEMA_signal_10305, new_AGEMA_signal_10301, new_AGEMA_signal_10297, new_AGEMA_signal_10293}), .c ({new_AGEMA_signal_7836, new_AGEMA_signal_7835, new_AGEMA_signal_7834, RoundReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7455, new_AGEMA_signal_7454, new_AGEMA_signal_7453, RoundOutput[14]}), .a ({new_AGEMA_signal_10321, new_AGEMA_signal_10317, new_AGEMA_signal_10313, new_AGEMA_signal_10309}), .c ({new_AGEMA_signal_7842, new_AGEMA_signal_7841, new_AGEMA_signal_7840, RoundReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7458, new_AGEMA_signal_7457, new_AGEMA_signal_7456, RoundOutput[15]}), .a ({new_AGEMA_signal_10337, new_AGEMA_signal_10333, new_AGEMA_signal_10329, new_AGEMA_signal_10325}), .c ({new_AGEMA_signal_7848, new_AGEMA_signal_7847, new_AGEMA_signal_7846, RoundReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7461, new_AGEMA_signal_7460, new_AGEMA_signal_7459, RoundOutput[16]}), .a ({new_AGEMA_signal_10353, new_AGEMA_signal_10349, new_AGEMA_signal_10345, new_AGEMA_signal_10341}), .c ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, new_AGEMA_signal_7852, RoundReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7929, new_AGEMA_signal_7928, new_AGEMA_signal_7927, RoundOutput[17]}), .a ({new_AGEMA_signal_10369, new_AGEMA_signal_10365, new_AGEMA_signal_10361, new_AGEMA_signal_10357}), .c ({new_AGEMA_signal_8181, new_AGEMA_signal_8180, new_AGEMA_signal_8179, RoundReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7464, new_AGEMA_signal_7463, new_AGEMA_signal_7462, RoundOutput[18]}), .a ({new_AGEMA_signal_10385, new_AGEMA_signal_10381, new_AGEMA_signal_10377, new_AGEMA_signal_10373}), .c ({new_AGEMA_signal_7860, new_AGEMA_signal_7859, new_AGEMA_signal_7858, RoundReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7932, new_AGEMA_signal_7931, new_AGEMA_signal_7930, RoundOutput[19]}), .a ({new_AGEMA_signal_10401, new_AGEMA_signal_10397, new_AGEMA_signal_10393, new_AGEMA_signal_10389}), .c ({new_AGEMA_signal_8187, new_AGEMA_signal_8186, new_AGEMA_signal_8185, RoundReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7935, new_AGEMA_signal_7934, new_AGEMA_signal_7933, RoundOutput[20]}), .a ({new_AGEMA_signal_10417, new_AGEMA_signal_10413, new_AGEMA_signal_10409, new_AGEMA_signal_10405}), .c ({new_AGEMA_signal_8193, new_AGEMA_signal_8192, new_AGEMA_signal_8191, RoundReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7467, new_AGEMA_signal_7466, new_AGEMA_signal_7465, RoundOutput[21]}), .a ({new_AGEMA_signal_10433, new_AGEMA_signal_10429, new_AGEMA_signal_10425, new_AGEMA_signal_10421}), .c ({new_AGEMA_signal_7866, new_AGEMA_signal_7865, new_AGEMA_signal_7864, RoundReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7470, new_AGEMA_signal_7469, new_AGEMA_signal_7468, RoundOutput[22]}), .a ({new_AGEMA_signal_10449, new_AGEMA_signal_10445, new_AGEMA_signal_10441, new_AGEMA_signal_10437}), .c ({new_AGEMA_signal_7872, new_AGEMA_signal_7871, new_AGEMA_signal_7870, RoundReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7473, new_AGEMA_signal_7472, new_AGEMA_signal_7471, RoundOutput[23]}), .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10461, new_AGEMA_signal_10457, new_AGEMA_signal_10453}), .c ({new_AGEMA_signal_7878, new_AGEMA_signal_7877, new_AGEMA_signal_7876, RoundReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7476, new_AGEMA_signal_7475, new_AGEMA_signal_7474, RoundOutput[24]}), .a ({new_AGEMA_signal_10481, new_AGEMA_signal_10477, new_AGEMA_signal_10473, new_AGEMA_signal_10469}), .c ({new_AGEMA_signal_7884, new_AGEMA_signal_7883, new_AGEMA_signal_7882, RoundReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7938, new_AGEMA_signal_7937, new_AGEMA_signal_7936, RoundOutput[25]}), .a ({new_AGEMA_signal_10497, new_AGEMA_signal_10493, new_AGEMA_signal_10489, new_AGEMA_signal_10485}), .c ({new_AGEMA_signal_8199, new_AGEMA_signal_8198, new_AGEMA_signal_8197, RoundReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7479, new_AGEMA_signal_7478, new_AGEMA_signal_7477, RoundOutput[26]}), .a ({new_AGEMA_signal_10513, new_AGEMA_signal_10509, new_AGEMA_signal_10505, new_AGEMA_signal_10501}), .c ({new_AGEMA_signal_7890, new_AGEMA_signal_7889, new_AGEMA_signal_7888, RoundReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7941, new_AGEMA_signal_7940, new_AGEMA_signal_7939, RoundOutput[27]}), .a ({new_AGEMA_signal_10529, new_AGEMA_signal_10525, new_AGEMA_signal_10521, new_AGEMA_signal_10517}), .c ({new_AGEMA_signal_8205, new_AGEMA_signal_8204, new_AGEMA_signal_8203, RoundReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7944, new_AGEMA_signal_7943, new_AGEMA_signal_7942, RoundOutput[28]}), .a ({new_AGEMA_signal_10545, new_AGEMA_signal_10541, new_AGEMA_signal_10537, new_AGEMA_signal_10533}), .c ({new_AGEMA_signal_8211, new_AGEMA_signal_8210, new_AGEMA_signal_8209, RoundReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7482, new_AGEMA_signal_7481, new_AGEMA_signal_7480, RoundOutput[29]}), .a ({new_AGEMA_signal_10561, new_AGEMA_signal_10557, new_AGEMA_signal_10553, new_AGEMA_signal_10549}), .c ({new_AGEMA_signal_7896, new_AGEMA_signal_7895, new_AGEMA_signal_7894, RoundReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, new_AGEMA_signal_7483, RoundOutput[30]}), .a ({new_AGEMA_signal_10577, new_AGEMA_signal_10573, new_AGEMA_signal_10569, new_AGEMA_signal_10565}), .c ({new_AGEMA_signal_7902, new_AGEMA_signal_7901, new_AGEMA_signal_7900, RoundReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7488, new_AGEMA_signal_7487, new_AGEMA_signal_7486, RoundOutput[31]}), .a ({new_AGEMA_signal_10593, new_AGEMA_signal_10589, new_AGEMA_signal_10585, new_AGEMA_signal_10581}), .c ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, new_AGEMA_signal_7906, RoundReg_Inst_ff_SDE_31_next_state}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_5265, new_AGEMA_signal_5264, new_AGEMA_signal_5263, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_10605, new_AGEMA_signal_10602, new_AGEMA_signal_10599, new_AGEMA_signal_10596}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_5403, new_AGEMA_signal_5402, new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_0_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_5217, new_AGEMA_signal_5216, new_AGEMA_signal_5215, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_10617, new_AGEMA_signal_10614, new_AGEMA_signal_10611, new_AGEMA_signal_10608}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_5268, new_AGEMA_signal_5267, new_AGEMA_signal_5266, SubBytesIns_Inst_Sbox_0_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_5214, new_AGEMA_signal_5213, new_AGEMA_signal_5212, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_10629, new_AGEMA_signal_10626, new_AGEMA_signal_10623, new_AGEMA_signal_10620}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_5271, new_AGEMA_signal_5270, new_AGEMA_signal_5269, SubBytesIns_Inst_Sbox_0_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_5262, new_AGEMA_signal_5261, new_AGEMA_signal_5260, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_10641, new_AGEMA_signal_10638, new_AGEMA_signal_10635, new_AGEMA_signal_10632}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810], Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_5406, new_AGEMA_signal_5405, new_AGEMA_signal_5404, SubBytesIns_Inst_Sbox_0_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_5211, new_AGEMA_signal_5210, new_AGEMA_signal_5209, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_10653, new_AGEMA_signal_10650, new_AGEMA_signal_10647, new_AGEMA_signal_10644}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_5274, new_AGEMA_signal_5273, new_AGEMA_signal_5272, SubBytesIns_Inst_Sbox_0_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_5208, new_AGEMA_signal_5207, new_AGEMA_signal_5206, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_10665, new_AGEMA_signal_10662, new_AGEMA_signal_10659, new_AGEMA_signal_10656}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_5277, new_AGEMA_signal_5276, new_AGEMA_signal_5275, SubBytesIns_Inst_Sbox_0_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_5259, new_AGEMA_signal_5258, new_AGEMA_signal_5257, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_10677, new_AGEMA_signal_10674, new_AGEMA_signal_10671, new_AGEMA_signal_10668}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_5409, new_AGEMA_signal_5408, new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_0_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, new_AGEMA_signal_5398, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_10689, new_AGEMA_signal_10686, new_AGEMA_signal_10683, new_AGEMA_signal_10680}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_5544, new_AGEMA_signal_5543, new_AGEMA_signal_5542, SubBytesIns_Inst_Sbox_0_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_5256, new_AGEMA_signal_5255, new_AGEMA_signal_5254, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_10701, new_AGEMA_signal_10698, new_AGEMA_signal_10695, new_AGEMA_signal_10692}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870], Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_5412, new_AGEMA_signal_5411, new_AGEMA_signal_5410, SubBytesIns_Inst_Sbox_0_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_5265, new_AGEMA_signal_5264, new_AGEMA_signal_5263, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_10713, new_AGEMA_signal_10710, new_AGEMA_signal_10707, new_AGEMA_signal_10704}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_5415, new_AGEMA_signal_5414, new_AGEMA_signal_5413, SubBytesIns_Inst_Sbox_0_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_5217, new_AGEMA_signal_5216, new_AGEMA_signal_5215, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_10725, new_AGEMA_signal_10722, new_AGEMA_signal_10719, new_AGEMA_signal_10716}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_5280, new_AGEMA_signal_5279, new_AGEMA_signal_5278, SubBytesIns_Inst_Sbox_0_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_5214, new_AGEMA_signal_5213, new_AGEMA_signal_5212, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_10737, new_AGEMA_signal_10734, new_AGEMA_signal_10731, new_AGEMA_signal_10728}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_5283, new_AGEMA_signal_5282, new_AGEMA_signal_5281, SubBytesIns_Inst_Sbox_0_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_5262, new_AGEMA_signal_5261, new_AGEMA_signal_5260, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_10749, new_AGEMA_signal_10746, new_AGEMA_signal_10743, new_AGEMA_signal_10740}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, new_AGEMA_signal_5416, SubBytesIns_Inst_Sbox_0_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_5211, new_AGEMA_signal_5210, new_AGEMA_signal_5209, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_10761, new_AGEMA_signal_10758, new_AGEMA_signal_10755, new_AGEMA_signal_10752}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930], Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_5286, new_AGEMA_signal_5285, new_AGEMA_signal_5284, SubBytesIns_Inst_Sbox_0_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_5208, new_AGEMA_signal_5207, new_AGEMA_signal_5206, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_10773, new_AGEMA_signal_10770, new_AGEMA_signal_10767, new_AGEMA_signal_10764}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942], Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_5289, new_AGEMA_signal_5288, new_AGEMA_signal_5287, SubBytesIns_Inst_Sbox_0_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_5259, new_AGEMA_signal_5258, new_AGEMA_signal_5257, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_10785, new_AGEMA_signal_10782, new_AGEMA_signal_10779, new_AGEMA_signal_10776}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_5421, new_AGEMA_signal_5420, new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_0_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, new_AGEMA_signal_5398, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_10797, new_AGEMA_signal_10794, new_AGEMA_signal_10791, new_AGEMA_signal_10788}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_5547, new_AGEMA_signal_5546, new_AGEMA_signal_5545, SubBytesIns_Inst_Sbox_0_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_5256, new_AGEMA_signal_5255, new_AGEMA_signal_5254, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_10809, new_AGEMA_signal_10806, new_AGEMA_signal_10803, new_AGEMA_signal_10800}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978], Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_5424, new_AGEMA_signal_5423, new_AGEMA_signal_5422, SubBytesIns_Inst_Sbox_0_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_5421, new_AGEMA_signal_5420, new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_5547, new_AGEMA_signal_5546, new_AGEMA_signal_5545, SubBytesIns_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_5664, new_AGEMA_signal_5663, new_AGEMA_signal_5662, SubBytesIns_Inst_Sbox_0_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_5274, new_AGEMA_signal_5273, new_AGEMA_signal_5272, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_5280, new_AGEMA_signal_5279, new_AGEMA_signal_5278, SubBytesIns_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_5427, new_AGEMA_signal_5426, new_AGEMA_signal_5425, SubBytesIns_Inst_Sbox_0_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_5403, new_AGEMA_signal_5402, new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_5271, new_AGEMA_signal_5270, new_AGEMA_signal_5269, SubBytesIns_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_5550, new_AGEMA_signal_5549, new_AGEMA_signal_5548, SubBytesIns_Inst_Sbox_0_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_5268, new_AGEMA_signal_5267, new_AGEMA_signal_5266, SubBytesIns_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_5415, new_AGEMA_signal_5414, new_AGEMA_signal_5413, SubBytesIns_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_5553, new_AGEMA_signal_5552, new_AGEMA_signal_5551, SubBytesIns_Inst_Sbox_0_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_5412, new_AGEMA_signal_5411, new_AGEMA_signal_5410, SubBytesIns_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, new_AGEMA_signal_5416, SubBytesIns_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_5556, new_AGEMA_signal_5555, new_AGEMA_signal_5554, SubBytesIns_Inst_Sbox_0_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_5406, new_AGEMA_signal_5405, new_AGEMA_signal_5404, SubBytesIns_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_5421, new_AGEMA_signal_5420, new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_5559, new_AGEMA_signal_5558, new_AGEMA_signal_5557, SubBytesIns_Inst_Sbox_0_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_5547, new_AGEMA_signal_5546, new_AGEMA_signal_5545, SubBytesIns_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_5559, new_AGEMA_signal_5558, new_AGEMA_signal_5557, SubBytesIns_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_5667, new_AGEMA_signal_5666, new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_0_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_5403, new_AGEMA_signal_5402, new_AGEMA_signal_5401, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_5553, new_AGEMA_signal_5552, new_AGEMA_signal_5551, SubBytesIns_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_5670, new_AGEMA_signal_5669, new_AGEMA_signal_5668, SubBytesIns_Inst_Sbox_0_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_5277, new_AGEMA_signal_5276, new_AGEMA_signal_5275, SubBytesIns_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_5286, new_AGEMA_signal_5285, new_AGEMA_signal_5284, SubBytesIns_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_5430, new_AGEMA_signal_5429, new_AGEMA_signal_5428, SubBytesIns_Inst_Sbox_0_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_5409, new_AGEMA_signal_5408, new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_5544, new_AGEMA_signal_5543, new_AGEMA_signal_5542, SubBytesIns_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_5673, new_AGEMA_signal_5672, new_AGEMA_signal_5671, SubBytesIns_Inst_Sbox_0_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_5544, new_AGEMA_signal_5543, new_AGEMA_signal_5542, SubBytesIns_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_5556, new_AGEMA_signal_5555, new_AGEMA_signal_5554, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_5676, new_AGEMA_signal_5675, new_AGEMA_signal_5674, SubBytesIns_Inst_Sbox_0_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_5289, new_AGEMA_signal_5288, new_AGEMA_signal_5287, SubBytesIns_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_5550, new_AGEMA_signal_5549, new_AGEMA_signal_5548, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_5679, new_AGEMA_signal_5678, new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_0_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_5271, new_AGEMA_signal_5270, new_AGEMA_signal_5269, SubBytesIns_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_5277, new_AGEMA_signal_5276, new_AGEMA_signal_5275, SubBytesIns_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_5433, new_AGEMA_signal_5432, new_AGEMA_signal_5431, SubBytesIns_Inst_Sbox_0_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_5274, new_AGEMA_signal_5273, new_AGEMA_signal_5272, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_5664, new_AGEMA_signal_5663, new_AGEMA_signal_5662, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_5772, new_AGEMA_signal_5771, new_AGEMA_signal_5770, SubBytesIns_Inst_Sbox_0_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_5409, new_AGEMA_signal_5408, new_AGEMA_signal_5407, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_5421, new_AGEMA_signal_5420, new_AGEMA_signal_5419, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_5562, new_AGEMA_signal_5561, new_AGEMA_signal_5560, SubBytesIns_Inst_Sbox_0_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_5415, new_AGEMA_signal_5414, new_AGEMA_signal_5413, SubBytesIns_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_5427, new_AGEMA_signal_5426, new_AGEMA_signal_5425, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_5565, new_AGEMA_signal_5564, new_AGEMA_signal_5563, SubBytesIns_Inst_Sbox_0_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_5280, new_AGEMA_signal_5279, new_AGEMA_signal_5278, SubBytesIns_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_5664, new_AGEMA_signal_5663, new_AGEMA_signal_5662, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_5775, new_AGEMA_signal_5774, new_AGEMA_signal_5773, SubBytesIns_Inst_Sbox_0_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_5283, new_AGEMA_signal_5282, new_AGEMA_signal_5281, SubBytesIns_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_5427, new_AGEMA_signal_5426, new_AGEMA_signal_5425, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, new_AGEMA_signal_5566, SubBytesIns_Inst_Sbox_0_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, new_AGEMA_signal_5416, SubBytesIns_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_5430, new_AGEMA_signal_5429, new_AGEMA_signal_5428, SubBytesIns_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_5571, new_AGEMA_signal_5570, new_AGEMA_signal_5569, SubBytesIns_Inst_Sbox_0_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_5424, new_AGEMA_signal_5423, new_AGEMA_signal_5422, SubBytesIns_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_5556, new_AGEMA_signal_5555, new_AGEMA_signal_5554, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_5682, new_AGEMA_signal_5681, new_AGEMA_signal_5680, SubBytesIns_Inst_Sbox_0_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_5664, new_AGEMA_signal_5663, new_AGEMA_signal_5662, SubBytesIns_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_5427, new_AGEMA_signal_5426, new_AGEMA_signal_5425, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, new_AGEMA_signal_5776, SubBytesIns_Inst_Sbox_0_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_5427, new_AGEMA_signal_5426, new_AGEMA_signal_5425, SubBytesIns_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_5670, new_AGEMA_signal_5669, new_AGEMA_signal_5668, SubBytesIns_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_5781, new_AGEMA_signal_5780, new_AGEMA_signal_5779, SubBytesIns_Inst_Sbox_0_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_5553, new_AGEMA_signal_5552, new_AGEMA_signal_5551, SubBytesIns_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_5433, new_AGEMA_signal_5432, new_AGEMA_signal_5431, SubBytesIns_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_5685, new_AGEMA_signal_5684, new_AGEMA_signal_5683, SubBytesIns_Inst_Sbox_0_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_5571, new_AGEMA_signal_5570, new_AGEMA_signal_5569, SubBytesIns_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_5550, new_AGEMA_signal_5549, new_AGEMA_signal_5548, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, new_AGEMA_signal_5686, SubBytesIns_Inst_Sbox_0_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_5565, new_AGEMA_signal_5564, new_AGEMA_signal_5563, SubBytesIns_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_5673, new_AGEMA_signal_5672, new_AGEMA_signal_5671, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, new_AGEMA_signal_5782, SubBytesIns_Inst_Sbox_0_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_5667, new_AGEMA_signal_5666, new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_5676, new_AGEMA_signal_5675, new_AGEMA_signal_5674, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_5787, new_AGEMA_signal_5786, new_AGEMA_signal_5785, SubBytesIns_Inst_Sbox_0_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_5670, new_AGEMA_signal_5669, new_AGEMA_signal_5668, SubBytesIns_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_5673, new_AGEMA_signal_5672, new_AGEMA_signal_5671, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_5790, new_AGEMA_signal_5789, new_AGEMA_signal_5788, SubBytesIns_Inst_Sbox_0_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_5430, new_AGEMA_signal_5429, new_AGEMA_signal_5428, SubBytesIns_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_5676, new_AGEMA_signal_5675, new_AGEMA_signal_5674, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_5793, new_AGEMA_signal_5792, new_AGEMA_signal_5791, SubBytesIns_Inst_Sbox_0_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_5679, new_AGEMA_signal_5678, new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_5562, new_AGEMA_signal_5561, new_AGEMA_signal_5560, SubBytesIns_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_5796, new_AGEMA_signal_5795, new_AGEMA_signal_5794, SubBytesIns_Inst_Sbox_0_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_5679, new_AGEMA_signal_5678, new_AGEMA_signal_5677, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, new_AGEMA_signal_5566, SubBytesIns_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_5799, new_AGEMA_signal_5798, new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_0_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_5667, new_AGEMA_signal_5666, new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, new_AGEMA_signal_5782, SubBytesIns_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, new_AGEMA_signal_5902, MixColumnsIns_DoubleBytes[0]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_5775, new_AGEMA_signal_5774, new_AGEMA_signal_5773, SubBytesIns_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_5790, new_AGEMA_signal_5789, new_AGEMA_signal_5788, SubBytesIns_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_5907, new_AGEMA_signal_5906, new_AGEMA_signal_5905, MixColumnsIns_DoubleBytes[7]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_5682, new_AGEMA_signal_5681, new_AGEMA_signal_5680, SubBytesIns_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_5796, new_AGEMA_signal_5795, new_AGEMA_signal_5794, SubBytesIns_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, new_AGEMA_signal_5908, MixColumnsIns_DoubleBytes[6]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_5667, new_AGEMA_signal_5666, new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_5781, new_AGEMA_signal_5780, new_AGEMA_signal_5779, SubBytesIns_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, MixColumnsIns_DoubleBytes[5]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, new_AGEMA_signal_5776, SubBytesIns_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_5685, new_AGEMA_signal_5684, new_AGEMA_signal_5683, SubBytesIns_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, new_AGEMA_signal_5914, SubBytesOutput[3]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_5787, new_AGEMA_signal_5786, new_AGEMA_signal_5785, SubBytesIns_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_5799, new_AGEMA_signal_5798, new_AGEMA_signal_5797, SubBytesIns_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesOutput[2]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_5772, new_AGEMA_signal_5771, new_AGEMA_signal_5770, SubBytesIns_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_5793, new_AGEMA_signal_5792, new_AGEMA_signal_5791, SubBytesIns_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, new_AGEMA_signal_5920, MixColumnsIns_DoubleBytes[2]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_5667, new_AGEMA_signal_5666, new_AGEMA_signal_5665, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, new_AGEMA_signal_5686, SubBytesIns_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, new_AGEMA_signal_5800, SubBytesOutput[0]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, new_AGEMA_signal_5299, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_10821, new_AGEMA_signal_10818, new_AGEMA_signal_10815, new_AGEMA_signal_10812}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990], Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_5439, new_AGEMA_signal_5438, new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_1_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_5229, new_AGEMA_signal_5228, new_AGEMA_signal_5227, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_10833, new_AGEMA_signal_10830, new_AGEMA_signal_10827, new_AGEMA_signal_10824}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_5304, new_AGEMA_signal_5303, new_AGEMA_signal_5302, SubBytesIns_Inst_Sbox_1_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_5226, new_AGEMA_signal_5225, new_AGEMA_signal_5224, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_10845, new_AGEMA_signal_10842, new_AGEMA_signal_10839, new_AGEMA_signal_10836}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_5307, new_AGEMA_signal_5306, new_AGEMA_signal_5305, SubBytesIns_Inst_Sbox_1_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_5298, new_AGEMA_signal_5297, new_AGEMA_signal_5296, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_10857, new_AGEMA_signal_10854, new_AGEMA_signal_10851, new_AGEMA_signal_10848}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026], Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_5442, new_AGEMA_signal_5441, new_AGEMA_signal_5440, SubBytesIns_Inst_Sbox_1_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_5223, new_AGEMA_signal_5222, new_AGEMA_signal_5221, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_10869, new_AGEMA_signal_10866, new_AGEMA_signal_10863, new_AGEMA_signal_10860}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038], Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_5310, new_AGEMA_signal_5309, new_AGEMA_signal_5308, SubBytesIns_Inst_Sbox_1_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_5220, new_AGEMA_signal_5219, new_AGEMA_signal_5218, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_10881, new_AGEMA_signal_10878, new_AGEMA_signal_10875, new_AGEMA_signal_10872}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050], Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_5313, new_AGEMA_signal_5312, new_AGEMA_signal_5311, SubBytesIns_Inst_Sbox_1_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_5295, new_AGEMA_signal_5294, new_AGEMA_signal_5293, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_10893, new_AGEMA_signal_10890, new_AGEMA_signal_10887, new_AGEMA_signal_10884}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062], Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_5445, new_AGEMA_signal_5444, new_AGEMA_signal_5443, SubBytesIns_Inst_Sbox_1_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_5436, new_AGEMA_signal_5435, new_AGEMA_signal_5434, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_10905, new_AGEMA_signal_10902, new_AGEMA_signal_10899, new_AGEMA_signal_10896}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074], Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_5574, new_AGEMA_signal_5573, new_AGEMA_signal_5572, SubBytesIns_Inst_Sbox_1_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_5292, new_AGEMA_signal_5291, new_AGEMA_signal_5290, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_10917, new_AGEMA_signal_10914, new_AGEMA_signal_10911, new_AGEMA_signal_10908}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086], Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_5448, new_AGEMA_signal_5447, new_AGEMA_signal_5446, SubBytesIns_Inst_Sbox_1_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, new_AGEMA_signal_5299, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_10929, new_AGEMA_signal_10926, new_AGEMA_signal_10923, new_AGEMA_signal_10920}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098], Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_5451, new_AGEMA_signal_5450, new_AGEMA_signal_5449, SubBytesIns_Inst_Sbox_1_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_5229, new_AGEMA_signal_5228, new_AGEMA_signal_5227, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_10941, new_AGEMA_signal_10938, new_AGEMA_signal_10935, new_AGEMA_signal_10932}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110], Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_5316, new_AGEMA_signal_5315, new_AGEMA_signal_5314, SubBytesIns_Inst_Sbox_1_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_5226, new_AGEMA_signal_5225, new_AGEMA_signal_5224, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_10953, new_AGEMA_signal_10950, new_AGEMA_signal_10947, new_AGEMA_signal_10944}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122], Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_5319, new_AGEMA_signal_5318, new_AGEMA_signal_5317, SubBytesIns_Inst_Sbox_1_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_5298, new_AGEMA_signal_5297, new_AGEMA_signal_5296, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_10965, new_AGEMA_signal_10962, new_AGEMA_signal_10959, new_AGEMA_signal_10956}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134], Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_5454, new_AGEMA_signal_5453, new_AGEMA_signal_5452, SubBytesIns_Inst_Sbox_1_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_5223, new_AGEMA_signal_5222, new_AGEMA_signal_5221, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_10977, new_AGEMA_signal_10974, new_AGEMA_signal_10971, new_AGEMA_signal_10968}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146], Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_5322, new_AGEMA_signal_5321, new_AGEMA_signal_5320, SubBytesIns_Inst_Sbox_1_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_5220, new_AGEMA_signal_5219, new_AGEMA_signal_5218, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_10989, new_AGEMA_signal_10986, new_AGEMA_signal_10983, new_AGEMA_signal_10980}), .clk (clk), .r ({Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158], Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({new_AGEMA_signal_5325, new_AGEMA_signal_5324, new_AGEMA_signal_5323, SubBytesIns_Inst_Sbox_1_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_5295, new_AGEMA_signal_5294, new_AGEMA_signal_5293, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_11001, new_AGEMA_signal_10998, new_AGEMA_signal_10995, new_AGEMA_signal_10992}), .clk (clk), .r ({Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170], Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({new_AGEMA_signal_5457, new_AGEMA_signal_5456, new_AGEMA_signal_5455, SubBytesIns_Inst_Sbox_1_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_5436, new_AGEMA_signal_5435, new_AGEMA_signal_5434, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_11013, new_AGEMA_signal_11010, new_AGEMA_signal_11007, new_AGEMA_signal_11004}), .clk (clk), .r ({Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182], Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({new_AGEMA_signal_5577, new_AGEMA_signal_5576, new_AGEMA_signal_5575, SubBytesIns_Inst_Sbox_1_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_5292, new_AGEMA_signal_5291, new_AGEMA_signal_5290, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_11025, new_AGEMA_signal_11022, new_AGEMA_signal_11019, new_AGEMA_signal_11016}), .clk (clk), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194], Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({new_AGEMA_signal_5460, new_AGEMA_signal_5459, new_AGEMA_signal_5458, SubBytesIns_Inst_Sbox_1_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_5457, new_AGEMA_signal_5456, new_AGEMA_signal_5455, SubBytesIns_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_5577, new_AGEMA_signal_5576, new_AGEMA_signal_5575, SubBytesIns_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_5691, new_AGEMA_signal_5690, new_AGEMA_signal_5689, SubBytesIns_Inst_Sbox_1_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_5310, new_AGEMA_signal_5309, new_AGEMA_signal_5308, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_5316, new_AGEMA_signal_5315, new_AGEMA_signal_5314, SubBytesIns_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_5463, new_AGEMA_signal_5462, new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_1_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_5439, new_AGEMA_signal_5438, new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_5307, new_AGEMA_signal_5306, new_AGEMA_signal_5305, SubBytesIns_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, new_AGEMA_signal_5578, SubBytesIns_Inst_Sbox_1_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_5304, new_AGEMA_signal_5303, new_AGEMA_signal_5302, SubBytesIns_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_5451, new_AGEMA_signal_5450, new_AGEMA_signal_5449, SubBytesIns_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_5583, new_AGEMA_signal_5582, new_AGEMA_signal_5581, SubBytesIns_Inst_Sbox_1_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_5448, new_AGEMA_signal_5447, new_AGEMA_signal_5446, SubBytesIns_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_5454, new_AGEMA_signal_5453, new_AGEMA_signal_5452, SubBytesIns_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, new_AGEMA_signal_5584, SubBytesIns_Inst_Sbox_1_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_5442, new_AGEMA_signal_5441, new_AGEMA_signal_5440, SubBytesIns_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_5457, new_AGEMA_signal_5456, new_AGEMA_signal_5455, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_5589, new_AGEMA_signal_5588, new_AGEMA_signal_5587, SubBytesIns_Inst_Sbox_1_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_5577, new_AGEMA_signal_5576, new_AGEMA_signal_5575, SubBytesIns_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_5589, new_AGEMA_signal_5588, new_AGEMA_signal_5587, SubBytesIns_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_5694, new_AGEMA_signal_5693, new_AGEMA_signal_5692, SubBytesIns_Inst_Sbox_1_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_5439, new_AGEMA_signal_5438, new_AGEMA_signal_5437, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_5583, new_AGEMA_signal_5582, new_AGEMA_signal_5581, SubBytesIns_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, new_AGEMA_signal_5695, SubBytesIns_Inst_Sbox_1_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_5313, new_AGEMA_signal_5312, new_AGEMA_signal_5311, SubBytesIns_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_5322, new_AGEMA_signal_5321, new_AGEMA_signal_5320, SubBytesIns_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_5466, new_AGEMA_signal_5465, new_AGEMA_signal_5464, SubBytesIns_Inst_Sbox_1_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_5445, new_AGEMA_signal_5444, new_AGEMA_signal_5443, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_5574, new_AGEMA_signal_5573, new_AGEMA_signal_5572, SubBytesIns_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_5700, new_AGEMA_signal_5699, new_AGEMA_signal_5698, SubBytesIns_Inst_Sbox_1_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_5574, new_AGEMA_signal_5573, new_AGEMA_signal_5572, SubBytesIns_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, new_AGEMA_signal_5584, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, new_AGEMA_signal_5701, SubBytesIns_Inst_Sbox_1_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_5325, new_AGEMA_signal_5324, new_AGEMA_signal_5323, SubBytesIns_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, new_AGEMA_signal_5578, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, new_AGEMA_signal_5704, SubBytesIns_Inst_Sbox_1_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_5307, new_AGEMA_signal_5306, new_AGEMA_signal_5305, SubBytesIns_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_5313, new_AGEMA_signal_5312, new_AGEMA_signal_5311, SubBytesIns_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_5469, new_AGEMA_signal_5468, new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_1_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_5310, new_AGEMA_signal_5309, new_AGEMA_signal_5308, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_5691, new_AGEMA_signal_5690, new_AGEMA_signal_5689, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_5805, new_AGEMA_signal_5804, new_AGEMA_signal_5803, SubBytesIns_Inst_Sbox_1_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_5445, new_AGEMA_signal_5444, new_AGEMA_signal_5443, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_5457, new_AGEMA_signal_5456, new_AGEMA_signal_5455, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_5592, new_AGEMA_signal_5591, new_AGEMA_signal_5590, SubBytesIns_Inst_Sbox_1_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_5451, new_AGEMA_signal_5450, new_AGEMA_signal_5449, SubBytesIns_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_5463, new_AGEMA_signal_5462, new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_5595, new_AGEMA_signal_5594, new_AGEMA_signal_5593, SubBytesIns_Inst_Sbox_1_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_5316, new_AGEMA_signal_5315, new_AGEMA_signal_5314, SubBytesIns_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_5691, new_AGEMA_signal_5690, new_AGEMA_signal_5689, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, new_AGEMA_signal_5806, SubBytesIns_Inst_Sbox_1_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_5319, new_AGEMA_signal_5318, new_AGEMA_signal_5317, SubBytesIns_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_5463, new_AGEMA_signal_5462, new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, SubBytesIns_Inst_Sbox_1_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_5454, new_AGEMA_signal_5453, new_AGEMA_signal_5452, SubBytesIns_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_5466, new_AGEMA_signal_5465, new_AGEMA_signal_5464, SubBytesIns_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_5601, new_AGEMA_signal_5600, new_AGEMA_signal_5599, SubBytesIns_Inst_Sbox_1_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_5460, new_AGEMA_signal_5459, new_AGEMA_signal_5458, SubBytesIns_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, new_AGEMA_signal_5584, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_5709, new_AGEMA_signal_5708, new_AGEMA_signal_5707, SubBytesIns_Inst_Sbox_1_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_5691, new_AGEMA_signal_5690, new_AGEMA_signal_5689, SubBytesIns_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_5463, new_AGEMA_signal_5462, new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_5811, new_AGEMA_signal_5810, new_AGEMA_signal_5809, SubBytesIns_Inst_Sbox_1_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_5463, new_AGEMA_signal_5462, new_AGEMA_signal_5461, SubBytesIns_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, new_AGEMA_signal_5695, SubBytesIns_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, new_AGEMA_signal_5812, SubBytesIns_Inst_Sbox_1_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_5583, new_AGEMA_signal_5582, new_AGEMA_signal_5581, SubBytesIns_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_5469, new_AGEMA_signal_5468, new_AGEMA_signal_5467, SubBytesIns_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_5712, new_AGEMA_signal_5711, new_AGEMA_signal_5710, SubBytesIns_Inst_Sbox_1_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_5601, new_AGEMA_signal_5600, new_AGEMA_signal_5599, SubBytesIns_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, new_AGEMA_signal_5578, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_5715, new_AGEMA_signal_5714, new_AGEMA_signal_5713, SubBytesIns_Inst_Sbox_1_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_5595, new_AGEMA_signal_5594, new_AGEMA_signal_5593, SubBytesIns_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_5700, new_AGEMA_signal_5699, new_AGEMA_signal_5698, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_5817, new_AGEMA_signal_5816, new_AGEMA_signal_5815, SubBytesIns_Inst_Sbox_1_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_5694, new_AGEMA_signal_5693, new_AGEMA_signal_5692, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, new_AGEMA_signal_5701, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_5820, new_AGEMA_signal_5819, new_AGEMA_signal_5818, SubBytesIns_Inst_Sbox_1_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, new_AGEMA_signal_5695, SubBytesIns_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_5700, new_AGEMA_signal_5699, new_AGEMA_signal_5698, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_1_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_5466, new_AGEMA_signal_5465, new_AGEMA_signal_5464, SubBytesIns_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, new_AGEMA_signal_5701, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_1_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, new_AGEMA_signal_5704, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_5592, new_AGEMA_signal_5591, new_AGEMA_signal_5590, SubBytesIns_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_5829, new_AGEMA_signal_5828, new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_1_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, new_AGEMA_signal_5704, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, SubBytesIns_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_5832, new_AGEMA_signal_5831, new_AGEMA_signal_5830, SubBytesIns_Inst_Sbox_1_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_5694, new_AGEMA_signal_5693, new_AGEMA_signal_5692, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_5817, new_AGEMA_signal_5816, new_AGEMA_signal_5815, SubBytesIns_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, KeyExpansionIns_tmp[23]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, new_AGEMA_signal_5806, SubBytesIns_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, new_AGEMA_signal_5926, KeyExpansionIns_tmp[22]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_5709, new_AGEMA_signal_5708, new_AGEMA_signal_5707, SubBytesIns_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_5829, new_AGEMA_signal_5828, new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_5931, new_AGEMA_signal_5930, new_AGEMA_signal_5929, KeyExpansionIns_tmp[21]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_5694, new_AGEMA_signal_5693, new_AGEMA_signal_5692, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, new_AGEMA_signal_5812, SubBytesIns_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, new_AGEMA_signal_5932, KeyExpansionIns_tmp[20]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_5811, new_AGEMA_signal_5810, new_AGEMA_signal_5809, SubBytesIns_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_5712, new_AGEMA_signal_5711, new_AGEMA_signal_5710, SubBytesIns_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_5937, new_AGEMA_signal_5936, new_AGEMA_signal_5935, KeyExpansionIns_tmp[19]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_5820, new_AGEMA_signal_5819, new_AGEMA_signal_5818, SubBytesIns_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_5832, new_AGEMA_signal_5831, new_AGEMA_signal_5830, SubBytesIns_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, new_AGEMA_signal_5938, KeyExpansionIns_tmp[18]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_5805, new_AGEMA_signal_5804, new_AGEMA_signal_5803, SubBytesIns_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, KeyExpansionIns_tmp[17]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_5694, new_AGEMA_signal_5693, new_AGEMA_signal_5692, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_5715, new_AGEMA_signal_5714, new_AGEMA_signal_5713, SubBytesIns_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, new_AGEMA_signal_5833, KeyExpansionIns_tmp[16]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_5337, new_AGEMA_signal_5336, new_AGEMA_signal_5335, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_11037, new_AGEMA_signal_11034, new_AGEMA_signal_11031, new_AGEMA_signal_11028}), .clk (clk), .r ({Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206], Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({new_AGEMA_signal_5475, new_AGEMA_signal_5474, new_AGEMA_signal_5473, SubBytesIns_Inst_Sbox_2_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_5241, new_AGEMA_signal_5240, new_AGEMA_signal_5239, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_11049, new_AGEMA_signal_11046, new_AGEMA_signal_11043, new_AGEMA_signal_11040}), .clk (clk), .r ({Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218], Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({new_AGEMA_signal_5340, new_AGEMA_signal_5339, new_AGEMA_signal_5338, SubBytesIns_Inst_Sbox_2_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_5238, new_AGEMA_signal_5237, new_AGEMA_signal_5236, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_11061, new_AGEMA_signal_11058, new_AGEMA_signal_11055, new_AGEMA_signal_11052}), .clk (clk), .r ({Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230], Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({new_AGEMA_signal_5343, new_AGEMA_signal_5342, new_AGEMA_signal_5341, SubBytesIns_Inst_Sbox_2_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_5334, new_AGEMA_signal_5333, new_AGEMA_signal_5332, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_11073, new_AGEMA_signal_11070, new_AGEMA_signal_11067, new_AGEMA_signal_11064}), .clk (clk), .r ({Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242], Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, new_AGEMA_signal_5476, SubBytesIns_Inst_Sbox_2_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_5235, new_AGEMA_signal_5234, new_AGEMA_signal_5233, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_11085, new_AGEMA_signal_11082, new_AGEMA_signal_11079, new_AGEMA_signal_11076}), .clk (clk), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254], Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, new_AGEMA_signal_5344, SubBytesIns_Inst_Sbox_2_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_5232, new_AGEMA_signal_5231, new_AGEMA_signal_5230, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_11097, new_AGEMA_signal_11094, new_AGEMA_signal_11091, new_AGEMA_signal_11088}), .clk (clk), .r ({Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266], Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({new_AGEMA_signal_5349, new_AGEMA_signal_5348, new_AGEMA_signal_5347, SubBytesIns_Inst_Sbox_2_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_5331, new_AGEMA_signal_5330, new_AGEMA_signal_5329, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_11109, new_AGEMA_signal_11106, new_AGEMA_signal_11103, new_AGEMA_signal_11100}), .clk (clk), .r ({Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278], Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({new_AGEMA_signal_5481, new_AGEMA_signal_5480, new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_2_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_5472, new_AGEMA_signal_5471, new_AGEMA_signal_5470, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_11121, new_AGEMA_signal_11118, new_AGEMA_signal_11115, new_AGEMA_signal_11112}), .clk (clk), .r ({Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290], Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({new_AGEMA_signal_5604, new_AGEMA_signal_5603, new_AGEMA_signal_5602, SubBytesIns_Inst_Sbox_2_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, new_AGEMA_signal_5326, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_11133, new_AGEMA_signal_11130, new_AGEMA_signal_11127, new_AGEMA_signal_11124}), .clk (clk), .r ({Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302], Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({new_AGEMA_signal_5484, new_AGEMA_signal_5483, new_AGEMA_signal_5482, SubBytesIns_Inst_Sbox_2_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_5337, new_AGEMA_signal_5336, new_AGEMA_signal_5335, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_11145, new_AGEMA_signal_11142, new_AGEMA_signal_11139, new_AGEMA_signal_11136}), .clk (clk), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314], Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({new_AGEMA_signal_5487, new_AGEMA_signal_5486, new_AGEMA_signal_5485, SubBytesIns_Inst_Sbox_2_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_5241, new_AGEMA_signal_5240, new_AGEMA_signal_5239, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_11157, new_AGEMA_signal_11154, new_AGEMA_signal_11151, new_AGEMA_signal_11148}), .clk (clk), .r ({Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326], Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({new_AGEMA_signal_5352, new_AGEMA_signal_5351, new_AGEMA_signal_5350, SubBytesIns_Inst_Sbox_2_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_5238, new_AGEMA_signal_5237, new_AGEMA_signal_5236, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_11169, new_AGEMA_signal_11166, new_AGEMA_signal_11163, new_AGEMA_signal_11160}), .clk (clk), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338], Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({new_AGEMA_signal_5355, new_AGEMA_signal_5354, new_AGEMA_signal_5353, SubBytesIns_Inst_Sbox_2_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_5334, new_AGEMA_signal_5333, new_AGEMA_signal_5332, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_11181, new_AGEMA_signal_11178, new_AGEMA_signal_11175, new_AGEMA_signal_11172}), .clk (clk), .r ({Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350], Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({new_AGEMA_signal_5490, new_AGEMA_signal_5489, new_AGEMA_signal_5488, SubBytesIns_Inst_Sbox_2_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_5235, new_AGEMA_signal_5234, new_AGEMA_signal_5233, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_11193, new_AGEMA_signal_11190, new_AGEMA_signal_11187, new_AGEMA_signal_11184}), .clk (clk), .r ({Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362], Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({new_AGEMA_signal_5358, new_AGEMA_signal_5357, new_AGEMA_signal_5356, SubBytesIns_Inst_Sbox_2_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_5232, new_AGEMA_signal_5231, new_AGEMA_signal_5230, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_11205, new_AGEMA_signal_11202, new_AGEMA_signal_11199, new_AGEMA_signal_11196}), .clk (clk), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374], Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({new_AGEMA_signal_5361, new_AGEMA_signal_5360, new_AGEMA_signal_5359, SubBytesIns_Inst_Sbox_2_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_5331, new_AGEMA_signal_5330, new_AGEMA_signal_5329, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_11217, new_AGEMA_signal_11214, new_AGEMA_signal_11211, new_AGEMA_signal_11208}), .clk (clk), .r ({Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386], Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({new_AGEMA_signal_5493, new_AGEMA_signal_5492, new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_2_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_5472, new_AGEMA_signal_5471, new_AGEMA_signal_5470, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_11229, new_AGEMA_signal_11226, new_AGEMA_signal_11223, new_AGEMA_signal_11220}), .clk (clk), .r ({Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398], Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({new_AGEMA_signal_5607, new_AGEMA_signal_5606, new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_2_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, new_AGEMA_signal_5326, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_11241, new_AGEMA_signal_11238, new_AGEMA_signal_11235, new_AGEMA_signal_11232}), .clk (clk), .r ({Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410], Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({new_AGEMA_signal_5496, new_AGEMA_signal_5495, new_AGEMA_signal_5494, SubBytesIns_Inst_Sbox_2_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_5493, new_AGEMA_signal_5492, new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_5607, new_AGEMA_signal_5606, new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, new_AGEMA_signal_5716, SubBytesIns_Inst_Sbox_2_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, new_AGEMA_signal_5344, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_5352, new_AGEMA_signal_5351, new_AGEMA_signal_5350, SubBytesIns_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_5499, new_AGEMA_signal_5498, new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_2_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_5475, new_AGEMA_signal_5474, new_AGEMA_signal_5473, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_5343, new_AGEMA_signal_5342, new_AGEMA_signal_5341, SubBytesIns_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_5610, new_AGEMA_signal_5609, new_AGEMA_signal_5608, SubBytesIns_Inst_Sbox_2_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_5340, new_AGEMA_signal_5339, new_AGEMA_signal_5338, SubBytesIns_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_5487, new_AGEMA_signal_5486, new_AGEMA_signal_5485, SubBytesIns_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_5613, new_AGEMA_signal_5612, new_AGEMA_signal_5611, SubBytesIns_Inst_Sbox_2_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_5484, new_AGEMA_signal_5483, new_AGEMA_signal_5482, SubBytesIns_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_5490, new_AGEMA_signal_5489, new_AGEMA_signal_5488, SubBytesIns_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_5616, new_AGEMA_signal_5615, new_AGEMA_signal_5614, SubBytesIns_Inst_Sbox_2_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, new_AGEMA_signal_5476, SubBytesIns_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_5493, new_AGEMA_signal_5492, new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_5619, new_AGEMA_signal_5618, new_AGEMA_signal_5617, SubBytesIns_Inst_Sbox_2_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_5607, new_AGEMA_signal_5606, new_AGEMA_signal_5605, SubBytesIns_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_5619, new_AGEMA_signal_5618, new_AGEMA_signal_5617, SubBytesIns_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_5721, new_AGEMA_signal_5720, new_AGEMA_signal_5719, SubBytesIns_Inst_Sbox_2_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_5475, new_AGEMA_signal_5474, new_AGEMA_signal_5473, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_5613, new_AGEMA_signal_5612, new_AGEMA_signal_5611, SubBytesIns_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_5724, new_AGEMA_signal_5723, new_AGEMA_signal_5722, SubBytesIns_Inst_Sbox_2_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_5349, new_AGEMA_signal_5348, new_AGEMA_signal_5347, SubBytesIns_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_5358, new_AGEMA_signal_5357, new_AGEMA_signal_5356, SubBytesIns_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_5502, new_AGEMA_signal_5501, new_AGEMA_signal_5500, SubBytesIns_Inst_Sbox_2_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_5481, new_AGEMA_signal_5480, new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_5604, new_AGEMA_signal_5603, new_AGEMA_signal_5602, SubBytesIns_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_5727, new_AGEMA_signal_5726, new_AGEMA_signal_5725, SubBytesIns_Inst_Sbox_2_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_5604, new_AGEMA_signal_5603, new_AGEMA_signal_5602, SubBytesIns_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_5616, new_AGEMA_signal_5615, new_AGEMA_signal_5614, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_5730, new_AGEMA_signal_5729, new_AGEMA_signal_5728, SubBytesIns_Inst_Sbox_2_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_5361, new_AGEMA_signal_5360, new_AGEMA_signal_5359, SubBytesIns_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_5610, new_AGEMA_signal_5609, new_AGEMA_signal_5608, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, new_AGEMA_signal_5731, SubBytesIns_Inst_Sbox_2_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_5343, new_AGEMA_signal_5342, new_AGEMA_signal_5341, SubBytesIns_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_5349, new_AGEMA_signal_5348, new_AGEMA_signal_5347, SubBytesIns_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_5505, new_AGEMA_signal_5504, new_AGEMA_signal_5503, SubBytesIns_Inst_Sbox_2_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, new_AGEMA_signal_5344, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, new_AGEMA_signal_5716, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, new_AGEMA_signal_5836, SubBytesIns_Inst_Sbox_2_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_5481, new_AGEMA_signal_5480, new_AGEMA_signal_5479, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_5493, new_AGEMA_signal_5492, new_AGEMA_signal_5491, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, new_AGEMA_signal_5620, SubBytesIns_Inst_Sbox_2_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_5487, new_AGEMA_signal_5486, new_AGEMA_signal_5485, SubBytesIns_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_5499, new_AGEMA_signal_5498, new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_5625, new_AGEMA_signal_5624, new_AGEMA_signal_5623, SubBytesIns_Inst_Sbox_2_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_5352, new_AGEMA_signal_5351, new_AGEMA_signal_5350, SubBytesIns_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, new_AGEMA_signal_5716, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_5841, new_AGEMA_signal_5840, new_AGEMA_signal_5839, SubBytesIns_Inst_Sbox_2_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_5355, new_AGEMA_signal_5354, new_AGEMA_signal_5353, SubBytesIns_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_5499, new_AGEMA_signal_5498, new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_5628, new_AGEMA_signal_5627, new_AGEMA_signal_5626, SubBytesIns_Inst_Sbox_2_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_5490, new_AGEMA_signal_5489, new_AGEMA_signal_5488, SubBytesIns_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_5502, new_AGEMA_signal_5501, new_AGEMA_signal_5500, SubBytesIns_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_5631, new_AGEMA_signal_5630, new_AGEMA_signal_5629, SubBytesIns_Inst_Sbox_2_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_5496, new_AGEMA_signal_5495, new_AGEMA_signal_5494, SubBytesIns_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_5616, new_AGEMA_signal_5615, new_AGEMA_signal_5614, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, new_AGEMA_signal_5734, SubBytesIns_Inst_Sbox_2_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, new_AGEMA_signal_5716, SubBytesIns_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_5499, new_AGEMA_signal_5498, new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_5844, new_AGEMA_signal_5843, new_AGEMA_signal_5842, SubBytesIns_Inst_Sbox_2_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_5499, new_AGEMA_signal_5498, new_AGEMA_signal_5497, SubBytesIns_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_5724, new_AGEMA_signal_5723, new_AGEMA_signal_5722, SubBytesIns_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_5847, new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_2_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_5613, new_AGEMA_signal_5612, new_AGEMA_signal_5611, SubBytesIns_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_5505, new_AGEMA_signal_5504, new_AGEMA_signal_5503, SubBytesIns_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_5739, new_AGEMA_signal_5738, new_AGEMA_signal_5737, SubBytesIns_Inst_Sbox_2_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_5631, new_AGEMA_signal_5630, new_AGEMA_signal_5629, SubBytesIns_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_5610, new_AGEMA_signal_5609, new_AGEMA_signal_5608, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, new_AGEMA_signal_5740, SubBytesIns_Inst_Sbox_2_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_5625, new_AGEMA_signal_5624, new_AGEMA_signal_5623, SubBytesIns_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_5727, new_AGEMA_signal_5726, new_AGEMA_signal_5725, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_5850, new_AGEMA_signal_5849, new_AGEMA_signal_5848, SubBytesIns_Inst_Sbox_2_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_5721, new_AGEMA_signal_5720, new_AGEMA_signal_5719, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_5730, new_AGEMA_signal_5729, new_AGEMA_signal_5728, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_5853, new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_2_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_5724, new_AGEMA_signal_5723, new_AGEMA_signal_5722, SubBytesIns_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_5727, new_AGEMA_signal_5726, new_AGEMA_signal_5725, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_2_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_5502, new_AGEMA_signal_5501, new_AGEMA_signal_5500, SubBytesIns_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_5730, new_AGEMA_signal_5729, new_AGEMA_signal_5728, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_5859, new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_2_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, new_AGEMA_signal_5731, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, new_AGEMA_signal_5620, SubBytesIns_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_2_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, new_AGEMA_signal_5731, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_5628, new_AGEMA_signal_5627, new_AGEMA_signal_5626, SubBytesIns_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_5865, new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_2_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_5721, new_AGEMA_signal_5720, new_AGEMA_signal_5719, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_5850, new_AGEMA_signal_5849, new_AGEMA_signal_5848, SubBytesIns_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, KeyExpansionIns_tmp[15]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_5841, new_AGEMA_signal_5840, new_AGEMA_signal_5839, SubBytesIns_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, new_AGEMA_signal_5947, KeyExpansionIns_tmp[14]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, new_AGEMA_signal_5734, SubBytesIns_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, new_AGEMA_signal_5950, KeyExpansionIns_tmp[13]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_5721, new_AGEMA_signal_5720, new_AGEMA_signal_5719, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_5847, new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, new_AGEMA_signal_5953, KeyExpansionIns_tmp[12]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_5844, new_AGEMA_signal_5843, new_AGEMA_signal_5842, SubBytesIns_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_5739, new_AGEMA_signal_5738, new_AGEMA_signal_5737, SubBytesIns_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, new_AGEMA_signal_5956, KeyExpansionIns_tmp[11]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_5853, new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_5865, new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_5961, new_AGEMA_signal_5960, new_AGEMA_signal_5959, KeyExpansionIns_tmp[10]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, new_AGEMA_signal_5836, SubBytesIns_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_5859, new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, new_AGEMA_signal_5962, KeyExpansionIns_tmp[9]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_5721, new_AGEMA_signal_5720, new_AGEMA_signal_5719, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, new_AGEMA_signal_5740, SubBytesIns_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, new_AGEMA_signal_5866, KeyExpansionIns_tmp[8]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_5373, new_AGEMA_signal_5372, new_AGEMA_signal_5371, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_11253, new_AGEMA_signal_11250, new_AGEMA_signal_11247, new_AGEMA_signal_11244}), .clk (clk), .r ({Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422], Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({new_AGEMA_signal_5511, new_AGEMA_signal_5510, new_AGEMA_signal_5509, SubBytesIns_Inst_Sbox_3_M46}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_5253, new_AGEMA_signal_5252, new_AGEMA_signal_5251, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_11265, new_AGEMA_signal_11262, new_AGEMA_signal_11259, new_AGEMA_signal_11256}), .clk (clk), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434], Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({new_AGEMA_signal_5376, new_AGEMA_signal_5375, new_AGEMA_signal_5374, SubBytesIns_Inst_Sbox_3_M47}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_5250, new_AGEMA_signal_5249, new_AGEMA_signal_5248, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_11277, new_AGEMA_signal_11274, new_AGEMA_signal_11271, new_AGEMA_signal_11268}), .clk (clk), .r ({Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446], Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({new_AGEMA_signal_5379, new_AGEMA_signal_5378, new_AGEMA_signal_5377, SubBytesIns_Inst_Sbox_3_M48}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_5370, new_AGEMA_signal_5369, new_AGEMA_signal_5368, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_11289, new_AGEMA_signal_11286, new_AGEMA_signal_11283, new_AGEMA_signal_11280}), .clk (clk), .r ({Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458], Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({new_AGEMA_signal_5514, new_AGEMA_signal_5513, new_AGEMA_signal_5512, SubBytesIns_Inst_Sbox_3_M49}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_5247, new_AGEMA_signal_5246, new_AGEMA_signal_5245, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_11301, new_AGEMA_signal_11298, new_AGEMA_signal_11295, new_AGEMA_signal_11292}), .clk (clk), .r ({Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470], Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, new_AGEMA_signal_5380, SubBytesIns_Inst_Sbox_3_M50}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_5244, new_AGEMA_signal_5243, new_AGEMA_signal_5242, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_11313, new_AGEMA_signal_11310, new_AGEMA_signal_11307, new_AGEMA_signal_11304}), .clk (clk), .r ({Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482], Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({new_AGEMA_signal_5385, new_AGEMA_signal_5384, new_AGEMA_signal_5383, SubBytesIns_Inst_Sbox_3_M51}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_5367, new_AGEMA_signal_5366, new_AGEMA_signal_5365, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_11325, new_AGEMA_signal_11322, new_AGEMA_signal_11319, new_AGEMA_signal_11316}), .clk (clk), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494], Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({new_AGEMA_signal_5517, new_AGEMA_signal_5516, new_AGEMA_signal_5515, SubBytesIns_Inst_Sbox_3_M52}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, new_AGEMA_signal_5506, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_11337, new_AGEMA_signal_11334, new_AGEMA_signal_11331, new_AGEMA_signal_11328}), .clk (clk), .r ({Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506], Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({new_AGEMA_signal_5634, new_AGEMA_signal_5633, new_AGEMA_signal_5632, SubBytesIns_Inst_Sbox_3_M53}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, new_AGEMA_signal_5362, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_11349, new_AGEMA_signal_11346, new_AGEMA_signal_11343, new_AGEMA_signal_11340}), .clk (clk), .r ({Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518], Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({new_AGEMA_signal_5520, new_AGEMA_signal_5519, new_AGEMA_signal_5518, SubBytesIns_Inst_Sbox_3_M54}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_5373, new_AGEMA_signal_5372, new_AGEMA_signal_5371, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_11361, new_AGEMA_signal_11358, new_AGEMA_signal_11355, new_AGEMA_signal_11352}), .clk (clk), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530], Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({new_AGEMA_signal_5523, new_AGEMA_signal_5522, new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_3_M55}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_5253, new_AGEMA_signal_5252, new_AGEMA_signal_5251, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_11373, new_AGEMA_signal_11370, new_AGEMA_signal_11367, new_AGEMA_signal_11364}), .clk (clk), .r ({Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542], Fresh[1541], Fresh[1540], Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536]}), .c ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, new_AGEMA_signal_5386, SubBytesIns_Inst_Sbox_3_M56}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_5250, new_AGEMA_signal_5249, new_AGEMA_signal_5248, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_11385, new_AGEMA_signal_11382, new_AGEMA_signal_11379, new_AGEMA_signal_11376}), .clk (clk), .r ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554], Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550], Fresh[1549], Fresh[1548]}), .c ({new_AGEMA_signal_5391, new_AGEMA_signal_5390, new_AGEMA_signal_5389, SubBytesIns_Inst_Sbox_3_M57}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_5370, new_AGEMA_signal_5369, new_AGEMA_signal_5368, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_11397, new_AGEMA_signal_11394, new_AGEMA_signal_11391, new_AGEMA_signal_11388}), .clk (clk), .r ({Fresh[1571], Fresh[1570], Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566], Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, new_AGEMA_signal_5524, SubBytesIns_Inst_Sbox_3_M58}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_5247, new_AGEMA_signal_5246, new_AGEMA_signal_5245, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_11409, new_AGEMA_signal_11406, new_AGEMA_signal_11403, new_AGEMA_signal_11400}), .clk (clk), .r ({Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580], Fresh[1579], Fresh[1578], Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572]}), .c ({new_AGEMA_signal_5394, new_AGEMA_signal_5393, new_AGEMA_signal_5392, SubBytesIns_Inst_Sbox_3_M59}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_5244, new_AGEMA_signal_5243, new_AGEMA_signal_5242, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_11421, new_AGEMA_signal_11418, new_AGEMA_signal_11415, new_AGEMA_signal_11412}), .clk (clk), .r ({Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590], Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584]}), .c ({new_AGEMA_signal_5397, new_AGEMA_signal_5396, new_AGEMA_signal_5395, SubBytesIns_Inst_Sbox_3_M60}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_5367, new_AGEMA_signal_5366, new_AGEMA_signal_5365, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_11433, new_AGEMA_signal_11430, new_AGEMA_signal_11427, new_AGEMA_signal_11424}), .clk (clk), .r ({Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602], Fresh[1601], Fresh[1600], Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596]}), .c ({new_AGEMA_signal_5529, new_AGEMA_signal_5528, new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_3_M61}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, new_AGEMA_signal_5506, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_11445, new_AGEMA_signal_11442, new_AGEMA_signal_11439, new_AGEMA_signal_11436}), .clk (clk), .r ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614], Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610], Fresh[1609], Fresh[1608]}), .c ({new_AGEMA_signal_5637, new_AGEMA_signal_5636, new_AGEMA_signal_5635, SubBytesIns_Inst_Sbox_3_M62}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, new_AGEMA_signal_5362, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_11457, new_AGEMA_signal_11454, new_AGEMA_signal_11451, new_AGEMA_signal_11448}), .clk (clk), .r ({Fresh[1631], Fresh[1630], Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626], Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({new_AGEMA_signal_5532, new_AGEMA_signal_5531, new_AGEMA_signal_5530, SubBytesIns_Inst_Sbox_3_M63}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_5529, new_AGEMA_signal_5528, new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_5637, new_AGEMA_signal_5636, new_AGEMA_signal_5635, SubBytesIns_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_5745, new_AGEMA_signal_5744, new_AGEMA_signal_5743, SubBytesIns_Inst_Sbox_3_L0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, new_AGEMA_signal_5380, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, new_AGEMA_signal_5386, SubBytesIns_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_5535, new_AGEMA_signal_5534, new_AGEMA_signal_5533, SubBytesIns_Inst_Sbox_3_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_5511, new_AGEMA_signal_5510, new_AGEMA_signal_5509, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_5379, new_AGEMA_signal_5378, new_AGEMA_signal_5377, SubBytesIns_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_5640, new_AGEMA_signal_5639, new_AGEMA_signal_5638, SubBytesIns_Inst_Sbox_3_L2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_5376, new_AGEMA_signal_5375, new_AGEMA_signal_5374, SubBytesIns_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_5523, new_AGEMA_signal_5522, new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_5643, new_AGEMA_signal_5642, new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_3_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_5520, new_AGEMA_signal_5519, new_AGEMA_signal_5518, SubBytesIns_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, new_AGEMA_signal_5524, SubBytesIns_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_5646, new_AGEMA_signal_5645, new_AGEMA_signal_5644, SubBytesIns_Inst_Sbox_3_L4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_5514, new_AGEMA_signal_5513, new_AGEMA_signal_5512, SubBytesIns_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_5529, new_AGEMA_signal_5528, new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_5649, new_AGEMA_signal_5648, new_AGEMA_signal_5647, SubBytesIns_Inst_Sbox_3_L5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_5637, new_AGEMA_signal_5636, new_AGEMA_signal_5635, SubBytesIns_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_5649, new_AGEMA_signal_5648, new_AGEMA_signal_5647, SubBytesIns_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, new_AGEMA_signal_5746, SubBytesIns_Inst_Sbox_3_L6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_5511, new_AGEMA_signal_5510, new_AGEMA_signal_5509, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_5643, new_AGEMA_signal_5642, new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_5751, new_AGEMA_signal_5750, new_AGEMA_signal_5749, SubBytesIns_Inst_Sbox_3_L7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_5385, new_AGEMA_signal_5384, new_AGEMA_signal_5383, SubBytesIns_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_5394, new_AGEMA_signal_5393, new_AGEMA_signal_5392, SubBytesIns_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_5538, new_AGEMA_signal_5537, new_AGEMA_signal_5536, SubBytesIns_Inst_Sbox_3_L8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_5517, new_AGEMA_signal_5516, new_AGEMA_signal_5515, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_5634, new_AGEMA_signal_5633, new_AGEMA_signal_5632, SubBytesIns_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_5754, new_AGEMA_signal_5753, new_AGEMA_signal_5752, SubBytesIns_Inst_Sbox_3_L9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_5634, new_AGEMA_signal_5633, new_AGEMA_signal_5632, SubBytesIns_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_5646, new_AGEMA_signal_5645, new_AGEMA_signal_5644, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_5757, new_AGEMA_signal_5756, new_AGEMA_signal_5755, SubBytesIns_Inst_Sbox_3_L10}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_5397, new_AGEMA_signal_5396, new_AGEMA_signal_5395, SubBytesIns_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_5640, new_AGEMA_signal_5639, new_AGEMA_signal_5638, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_5760, new_AGEMA_signal_5759, new_AGEMA_signal_5758, SubBytesIns_Inst_Sbox_3_L11}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_5379, new_AGEMA_signal_5378, new_AGEMA_signal_5377, SubBytesIns_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_5385, new_AGEMA_signal_5384, new_AGEMA_signal_5383, SubBytesIns_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_5541, new_AGEMA_signal_5540, new_AGEMA_signal_5539, SubBytesIns_Inst_Sbox_3_L12}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, new_AGEMA_signal_5380, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_5745, new_AGEMA_signal_5744, new_AGEMA_signal_5743, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_5871, new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_3_L13}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_5517, new_AGEMA_signal_5516, new_AGEMA_signal_5515, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_5529, new_AGEMA_signal_5528, new_AGEMA_signal_5527, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_5652, new_AGEMA_signal_5651, new_AGEMA_signal_5650, SubBytesIns_Inst_Sbox_3_L14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_5523, new_AGEMA_signal_5522, new_AGEMA_signal_5521, SubBytesIns_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_5535, new_AGEMA_signal_5534, new_AGEMA_signal_5533, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_5655, new_AGEMA_signal_5654, new_AGEMA_signal_5653, SubBytesIns_Inst_Sbox_3_L15}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, new_AGEMA_signal_5386, SubBytesIns_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_5745, new_AGEMA_signal_5744, new_AGEMA_signal_5743, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_5874, new_AGEMA_signal_5873, new_AGEMA_signal_5872, SubBytesIns_Inst_Sbox_3_L16}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_5391, new_AGEMA_signal_5390, new_AGEMA_signal_5389, SubBytesIns_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_5535, new_AGEMA_signal_5534, new_AGEMA_signal_5533, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, new_AGEMA_signal_5656, SubBytesIns_Inst_Sbox_3_L17}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, new_AGEMA_signal_5524, SubBytesIns_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_5538, new_AGEMA_signal_5537, new_AGEMA_signal_5536, SubBytesIns_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_5661, new_AGEMA_signal_5660, new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_3_L18}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_5532, new_AGEMA_signal_5531, new_AGEMA_signal_5530, SubBytesIns_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_5646, new_AGEMA_signal_5645, new_AGEMA_signal_5644, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, new_AGEMA_signal_5761, SubBytesIns_Inst_Sbox_3_L19}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_5745, new_AGEMA_signal_5744, new_AGEMA_signal_5743, SubBytesIns_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_5535, new_AGEMA_signal_5534, new_AGEMA_signal_5533, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_5877, new_AGEMA_signal_5876, new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_3_L20}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_5535, new_AGEMA_signal_5534, new_AGEMA_signal_5533, SubBytesIns_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_5751, new_AGEMA_signal_5750, new_AGEMA_signal_5749, SubBytesIns_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_5880, new_AGEMA_signal_5879, new_AGEMA_signal_5878, SubBytesIns_Inst_Sbox_3_L21}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_5643, new_AGEMA_signal_5642, new_AGEMA_signal_5641, SubBytesIns_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_5541, new_AGEMA_signal_5540, new_AGEMA_signal_5539, SubBytesIns_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, new_AGEMA_signal_5764, SubBytesIns_Inst_Sbox_3_L22}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_5661, new_AGEMA_signal_5660, new_AGEMA_signal_5659, SubBytesIns_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_5640, new_AGEMA_signal_5639, new_AGEMA_signal_5638, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_5769, new_AGEMA_signal_5768, new_AGEMA_signal_5767, SubBytesIns_Inst_Sbox_3_L23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_5655, new_AGEMA_signal_5654, new_AGEMA_signal_5653, SubBytesIns_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_5754, new_AGEMA_signal_5753, new_AGEMA_signal_5752, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_3_L24}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, new_AGEMA_signal_5746, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_5757, new_AGEMA_signal_5756, new_AGEMA_signal_5755, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_3_L25}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_5751, new_AGEMA_signal_5750, new_AGEMA_signal_5749, SubBytesIns_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_5754, new_AGEMA_signal_5753, new_AGEMA_signal_5752, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_5889, new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_3_L26}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_5538, new_AGEMA_signal_5537, new_AGEMA_signal_5536, SubBytesIns_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_5757, new_AGEMA_signal_5756, new_AGEMA_signal_5755, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_5892, new_AGEMA_signal_5891, new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_3_L27}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_5760, new_AGEMA_signal_5759, new_AGEMA_signal_5758, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_5652, new_AGEMA_signal_5651, new_AGEMA_signal_5650, SubBytesIns_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_5895, new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_3_L28}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_5760, new_AGEMA_signal_5759, new_AGEMA_signal_5758, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, new_AGEMA_signal_5656, SubBytesIns_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_3_L29}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, new_AGEMA_signal_5746, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, new_AGEMA_signal_5965, KeyExpansionIns_tmp[7]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_5874, new_AGEMA_signal_5873, new_AGEMA_signal_5872, SubBytesIns_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_5889, new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, new_AGEMA_signal_5968, KeyExpansionIns_tmp[6]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, new_AGEMA_signal_5761, SubBytesIns_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_5895, new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, KeyExpansionIns_tmp[5]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, new_AGEMA_signal_5746, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_5880, new_AGEMA_signal_5879, new_AGEMA_signal_5878, SubBytesIns_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, new_AGEMA_signal_5974, KeyExpansionIns_tmp[4]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_5877, new_AGEMA_signal_5876, new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, new_AGEMA_signal_5764, SubBytesIns_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, new_AGEMA_signal_5977, KeyExpansionIns_tmp[3]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, new_AGEMA_signal_5980, KeyExpansionIns_tmp[2]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_5871, new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_5892, new_AGEMA_signal_5891, new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_5985, new_AGEMA_signal_5984, new_AGEMA_signal_5983, KeyExpansionIns_tmp[1]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, new_AGEMA_signal_5746, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_5769, new_AGEMA_signal_5768, new_AGEMA_signal_5767, SubBytesIns_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_5901, new_AGEMA_signal_5900, new_AGEMA_signal_5899, KeyExpansionIns_tmp[0]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U96 ( .a ({new_AGEMA_signal_6486, new_AGEMA_signal_6485, new_AGEMA_signal_6484, MixColumnsIns_n64}), .b ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, new_AGEMA_signal_5962, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_6924, new_AGEMA_signal_6923, new_AGEMA_signal_6922, MixColumnsOutput[9]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U95 ( .a ({new_AGEMA_signal_6264, new_AGEMA_signal_6263, new_AGEMA_signal_6262, MixColumnsIns_n63}), .b ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, new_AGEMA_signal_6250, MixColumnsIns_n62}), .c ({new_AGEMA_signal_6486, new_AGEMA_signal_6485, new_AGEMA_signal_6484, MixColumnsIns_n64}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U94 ( .a ({new_AGEMA_signal_6201, new_AGEMA_signal_6200, new_AGEMA_signal_6199, MixColumnsIns_n61}), .b ({new_AGEMA_signal_6027, new_AGEMA_signal_6026, new_AGEMA_signal_6025, MixColumnsIns_n60}), .c ({new_AGEMA_signal_6489, new_AGEMA_signal_6488, new_AGEMA_signal_6487, MixColumnsOutput[8]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U93 ( .a ({new_AGEMA_signal_6057, new_AGEMA_signal_6056, new_AGEMA_signal_6055, MixColumnsIns_n59}), .b ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, new_AGEMA_signal_5866, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_6201, new_AGEMA_signal_6200, new_AGEMA_signal_6199, MixColumnsIns_n61}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U92 ( .a ({new_AGEMA_signal_6204, new_AGEMA_signal_6203, new_AGEMA_signal_6202, MixColumnsIns_n58}), .b ({new_AGEMA_signal_6000, new_AGEMA_signal_5999, new_AGEMA_signal_5998, MixColumnsIns_n57}), .c ({new_AGEMA_signal_6492, new_AGEMA_signal_6491, new_AGEMA_signal_6490, MixColumnsOutput[7]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U91 ( .a ({new_AGEMA_signal_6033, new_AGEMA_signal_6032, new_AGEMA_signal_6031, MixColumnsIns_n56}), .b ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_6204, new_AGEMA_signal_6203, new_AGEMA_signal_6202, MixColumnsIns_n58}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U90 ( .a ({new_AGEMA_signal_6207, new_AGEMA_signal_6206, new_AGEMA_signal_6205, MixColumnsIns_n55}), .b ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, new_AGEMA_signal_6001, MixColumnsIns_n54}), .c ({new_AGEMA_signal_6495, new_AGEMA_signal_6494, new_AGEMA_signal_6493, MixColumnsOutput[6]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U89 ( .a ({new_AGEMA_signal_6039, new_AGEMA_signal_6038, new_AGEMA_signal_6037, MixColumnsIns_n53}), .b ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, new_AGEMA_signal_5926, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_6207, new_AGEMA_signal_6206, new_AGEMA_signal_6205, MixColumnsIns_n55}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U88 ( .a ({new_AGEMA_signal_6210, new_AGEMA_signal_6209, new_AGEMA_signal_6208, MixColumnsIns_n52}), .b ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, new_AGEMA_signal_6004, MixColumnsIns_n51}), .c ({new_AGEMA_signal_6498, new_AGEMA_signal_6497, new_AGEMA_signal_6496, MixColumnsOutput[5]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U87 ( .a ({new_AGEMA_signal_6045, new_AGEMA_signal_6044, new_AGEMA_signal_6043, MixColumnsIns_n50}), .b ({new_AGEMA_signal_5931, new_AGEMA_signal_5930, new_AGEMA_signal_5929, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_6210, new_AGEMA_signal_6209, new_AGEMA_signal_6208, MixColumnsIns_n52}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U86 ( .a ({new_AGEMA_signal_6501, new_AGEMA_signal_6500, new_AGEMA_signal_6499, MixColumnsIns_n49}), .b ({new_AGEMA_signal_6225, new_AGEMA_signal_6224, new_AGEMA_signal_6223, MixColumnsIns_n48}), .c ({new_AGEMA_signal_6927, new_AGEMA_signal_6926, new_AGEMA_signal_6925, MixColumnsOutput[4]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U85 ( .a ({new_AGEMA_signal_6282, new_AGEMA_signal_6281, new_AGEMA_signal_6280, MixColumnsIns_n47}), .b ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, new_AGEMA_signal_5932, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_6501, new_AGEMA_signal_6500, new_AGEMA_signal_6499, MixColumnsIns_n49}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U84 ( .a ({new_AGEMA_signal_6504, new_AGEMA_signal_6503, new_AGEMA_signal_6502, MixColumnsIns_n46}), .b ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, new_AGEMA_signal_6226, MixColumnsIns_n45}), .c ({new_AGEMA_signal_6930, new_AGEMA_signal_6929, new_AGEMA_signal_6928, MixColumnsOutput[3]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U83 ( .a ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, new_AGEMA_signal_6286, MixColumnsIns_n44}), .b ({new_AGEMA_signal_5937, new_AGEMA_signal_5936, new_AGEMA_signal_5935, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_6504, new_AGEMA_signal_6503, new_AGEMA_signal_6502, MixColumnsIns_n46}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U82 ( .a ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, new_AGEMA_signal_6211, MixColumnsIns_n43}), .b ({new_AGEMA_signal_6000, new_AGEMA_signal_5999, new_AGEMA_signal_5998, MixColumnsIns_n57}), .c ({new_AGEMA_signal_6507, new_AGEMA_signal_6506, new_AGEMA_signal_6505, MixColumnsOutput[31]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U81 ( .a ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, new_AGEMA_signal_5968, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_6000, new_AGEMA_signal_5999, new_AGEMA_signal_5998, MixColumnsIns_n57}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U80 ( .a ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, new_AGEMA_signal_5902, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_6012, new_AGEMA_signal_6011, new_AGEMA_signal_6010, MixColumnsIns_n42}), .c ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, new_AGEMA_signal_6211, MixColumnsIns_n43}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U79 ( .a ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, new_AGEMA_signal_6214, MixColumnsIns_n41}), .b ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, new_AGEMA_signal_6001, MixColumnsIns_n54}), .c ({new_AGEMA_signal_6510, new_AGEMA_signal_6509, new_AGEMA_signal_6508, MixColumnsOutput[30]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U78 ( .a ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, new_AGEMA_signal_5947, KeyExpansionIns_tmp[14]}), .b ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, new_AGEMA_signal_6001, MixColumnsIns_n54}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U77 ( .a ({new_AGEMA_signal_5907, new_AGEMA_signal_5906, new_AGEMA_signal_5905, MixColumnsIns_DoubleBytes[7]}), .b ({new_AGEMA_signal_6015, new_AGEMA_signal_6014, new_AGEMA_signal_6013, MixColumnsIns_n40}), .c ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, new_AGEMA_signal_6214, MixColumnsIns_n41}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U76 ( .a ({new_AGEMA_signal_6219, new_AGEMA_signal_6218, new_AGEMA_signal_6217, MixColumnsIns_n39}), .b ({new_AGEMA_signal_6009, new_AGEMA_signal_6008, new_AGEMA_signal_6007, MixColumnsIns_n38}), .c ({new_AGEMA_signal_6513, new_AGEMA_signal_6512, new_AGEMA_signal_6511, MixColumnsOutput[2]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U75 ( .a ({new_AGEMA_signal_6051, new_AGEMA_signal_6050, new_AGEMA_signal_6049, MixColumnsIns_n37}), .b ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, new_AGEMA_signal_5938, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_6219, new_AGEMA_signal_6218, new_AGEMA_signal_6217, MixColumnsIns_n39}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U74 ( .a ({new_AGEMA_signal_6222, new_AGEMA_signal_6221, new_AGEMA_signal_6220, MixColumnsIns_n36}), .b ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, new_AGEMA_signal_6004, MixColumnsIns_n51}), .c ({new_AGEMA_signal_6516, new_AGEMA_signal_6515, new_AGEMA_signal_6514, MixColumnsOutput[29]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U73 ( .a ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, new_AGEMA_signal_5950, KeyExpansionIns_tmp[13]}), .b ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, new_AGEMA_signal_5974, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, new_AGEMA_signal_6004, MixColumnsIns_n51}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U72 ( .a ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, new_AGEMA_signal_5908, MixColumnsIns_DoubleBytes[6]}), .b ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, new_AGEMA_signal_6016, MixColumnsIns_n35}), .c ({new_AGEMA_signal_6222, new_AGEMA_signal_6221, new_AGEMA_signal_6220, MixColumnsIns_n36}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U71 ( .a ({new_AGEMA_signal_6519, new_AGEMA_signal_6518, new_AGEMA_signal_6517, MixColumnsIns_n34}), .b ({new_AGEMA_signal_6225, new_AGEMA_signal_6224, new_AGEMA_signal_6223, MixColumnsIns_n48}), .c ({new_AGEMA_signal_6933, new_AGEMA_signal_6932, new_AGEMA_signal_6931, MixColumnsOutput[28]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U70 ( .a ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, new_AGEMA_signal_5953, KeyExpansionIns_tmp[12]}), .b ({new_AGEMA_signal_6060, new_AGEMA_signal_6059, new_AGEMA_signal_6058, MixColumnsIns_DoubleBytes[28]}), .c ({new_AGEMA_signal_6225, new_AGEMA_signal_6224, new_AGEMA_signal_6223, MixColumnsIns_n48}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U69 ( .a ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, MixColumnsIns_DoubleBytes[5]}), .b ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, new_AGEMA_signal_6244, MixColumnsIns_n33}), .c ({new_AGEMA_signal_6519, new_AGEMA_signal_6518, new_AGEMA_signal_6517, MixColumnsIns_n34}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U68 ( .a ({new_AGEMA_signal_6522, new_AGEMA_signal_6521, new_AGEMA_signal_6520, MixColumnsIns_n32}), .b ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, new_AGEMA_signal_6226, MixColumnsIns_n45}), .c ({new_AGEMA_signal_6936, new_AGEMA_signal_6935, new_AGEMA_signal_6934, MixColumnsOutput[27]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U67 ( .a ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, new_AGEMA_signal_5956, KeyExpansionIns_tmp[11]}), .b ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, new_AGEMA_signal_6061, MixColumnsIns_DoubleBytes[27]}), .c ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, new_AGEMA_signal_6226, MixColumnsIns_n45}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U66 ( .a ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, new_AGEMA_signal_5914, SubBytesOutput[3]}), .b ({new_AGEMA_signal_6255, new_AGEMA_signal_6254, new_AGEMA_signal_6253, MixColumnsIns_n31}), .c ({new_AGEMA_signal_6522, new_AGEMA_signal_6521, new_AGEMA_signal_6520, MixColumnsIns_n32}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U65 ( .a ({new_AGEMA_signal_6231, new_AGEMA_signal_6230, new_AGEMA_signal_6229, MixColumnsIns_n30}), .b ({new_AGEMA_signal_6009, new_AGEMA_signal_6008, new_AGEMA_signal_6007, MixColumnsIns_n38}), .c ({new_AGEMA_signal_6525, new_AGEMA_signal_6524, new_AGEMA_signal_6523, MixColumnsOutput[26]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U64 ( .a ({new_AGEMA_signal_5961, new_AGEMA_signal_5960, new_AGEMA_signal_5959, KeyExpansionIns_tmp[10]}), .b ({new_AGEMA_signal_5985, new_AGEMA_signal_5984, new_AGEMA_signal_5983, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_6009, new_AGEMA_signal_6008, new_AGEMA_signal_6007, MixColumnsIns_n38}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U63 ( .a ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesOutput[2]}), .b ({new_AGEMA_signal_6021, new_AGEMA_signal_6020, new_AGEMA_signal_6019, MixColumnsIns_n29}), .c ({new_AGEMA_signal_6231, new_AGEMA_signal_6230, new_AGEMA_signal_6229, MixColumnsIns_n30}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U62 ( .a ({new_AGEMA_signal_6528, new_AGEMA_signal_6527, new_AGEMA_signal_6526, MixColumnsIns_n28}), .b ({new_AGEMA_signal_6249, new_AGEMA_signal_6248, new_AGEMA_signal_6247, MixColumnsIns_n27}), .c ({new_AGEMA_signal_6939, new_AGEMA_signal_6938, new_AGEMA_signal_6937, MixColumnsOutput[25]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U61 ( .a ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, new_AGEMA_signal_5920, MixColumnsIns_DoubleBytes[2]}), .b ({new_AGEMA_signal_6261, new_AGEMA_signal_6260, new_AGEMA_signal_6259, MixColumnsIns_n26}), .c ({new_AGEMA_signal_6528, new_AGEMA_signal_6527, new_AGEMA_signal_6526, MixColumnsIns_n28}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U60 ( .a ({new_AGEMA_signal_6234, new_AGEMA_signal_6233, new_AGEMA_signal_6232, MixColumnsIns_n25}), .b ({new_AGEMA_signal_6024, new_AGEMA_signal_6023, new_AGEMA_signal_6022, MixColumnsIns_n24}), .c ({new_AGEMA_signal_6531, new_AGEMA_signal_6530, new_AGEMA_signal_6529, MixColumnsOutput[24]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U59 ( .a ({new_AGEMA_signal_6054, new_AGEMA_signal_6053, new_AGEMA_signal_6052, MixColumnsIns_n23}), .b ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, new_AGEMA_signal_5800, SubBytesOutput[0]}), .c ({new_AGEMA_signal_6234, new_AGEMA_signal_6233, new_AGEMA_signal_6232, MixColumnsIns_n25}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U58 ( .a ({new_AGEMA_signal_6237, new_AGEMA_signal_6236, new_AGEMA_signal_6235, MixColumnsIns_n22}), .b ({new_AGEMA_signal_6012, new_AGEMA_signal_6011, new_AGEMA_signal_6010, MixColumnsIns_n42}), .c ({new_AGEMA_signal_6534, new_AGEMA_signal_6533, new_AGEMA_signal_6532, MixColumnsOutput[23]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U57 ( .a ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, new_AGEMA_signal_5947, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_6012, new_AGEMA_signal_6011, new_AGEMA_signal_6010, MixColumnsIns_n42}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U56 ( .a ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, new_AGEMA_signal_5965, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_6030, new_AGEMA_signal_6029, new_AGEMA_signal_6028, MixColumnsIns_n21}), .c ({new_AGEMA_signal_6237, new_AGEMA_signal_6236, new_AGEMA_signal_6235, MixColumnsIns_n22}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U55 ( .a ({new_AGEMA_signal_6240, new_AGEMA_signal_6239, new_AGEMA_signal_6238, MixColumnsIns_n20}), .b ({new_AGEMA_signal_6015, new_AGEMA_signal_6014, new_AGEMA_signal_6013, MixColumnsIns_n40}), .c ({new_AGEMA_signal_6537, new_AGEMA_signal_6536, new_AGEMA_signal_6535, MixColumnsOutput[22]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U54 ( .a ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, new_AGEMA_signal_5926, KeyExpansionIns_tmp[22]}), .b ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, new_AGEMA_signal_5950, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_6015, new_AGEMA_signal_6014, new_AGEMA_signal_6013, MixColumnsIns_n40}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U53 ( .a ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, new_AGEMA_signal_5968, KeyExpansionIns_tmp[6]}), .b ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, new_AGEMA_signal_6034, MixColumnsIns_n19}), .c ({new_AGEMA_signal_6240, new_AGEMA_signal_6239, new_AGEMA_signal_6238, MixColumnsIns_n20}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U52 ( .a ({new_AGEMA_signal_6243, new_AGEMA_signal_6242, new_AGEMA_signal_6241, MixColumnsIns_n18}), .b ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, new_AGEMA_signal_6016, MixColumnsIns_n35}), .c ({new_AGEMA_signal_6540, new_AGEMA_signal_6539, new_AGEMA_signal_6538, MixColumnsOutput[21]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U51 ( .a ({new_AGEMA_signal_5931, new_AGEMA_signal_5930, new_AGEMA_signal_5929, KeyExpansionIns_tmp[21]}), .b ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, new_AGEMA_signal_5953, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, new_AGEMA_signal_6016, MixColumnsIns_n35}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U50 ( .a ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, KeyExpansionIns_tmp[5]}), .b ({new_AGEMA_signal_6042, new_AGEMA_signal_6041, new_AGEMA_signal_6040, MixColumnsIns_n17}), .c ({new_AGEMA_signal_6243, new_AGEMA_signal_6242, new_AGEMA_signal_6241, MixColumnsIns_n18}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U49 ( .a ({new_AGEMA_signal_6543, new_AGEMA_signal_6542, new_AGEMA_signal_6541, MixColumnsIns_n16}), .b ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, new_AGEMA_signal_6244, MixColumnsIns_n33}), .c ({new_AGEMA_signal_6942, new_AGEMA_signal_6941, new_AGEMA_signal_6940, MixColumnsOutput[20]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U48 ( .a ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, new_AGEMA_signal_5932, KeyExpansionIns_tmp[20]}), .b ({new_AGEMA_signal_6069, new_AGEMA_signal_6068, new_AGEMA_signal_6067, MixColumnsIns_DoubleBytes[20]}), .c ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, new_AGEMA_signal_6244, MixColumnsIns_n33}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U47 ( .a ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, new_AGEMA_signal_5974, KeyExpansionIns_tmp[4]}), .b ({new_AGEMA_signal_6279, new_AGEMA_signal_6278, new_AGEMA_signal_6277, MixColumnsIns_n15}), .c ({new_AGEMA_signal_6543, new_AGEMA_signal_6542, new_AGEMA_signal_6541, MixColumnsIns_n16}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U46 ( .a ({new_AGEMA_signal_6546, new_AGEMA_signal_6545, new_AGEMA_signal_6544, MixColumnsIns_n14}), .b ({new_AGEMA_signal_6249, new_AGEMA_signal_6248, new_AGEMA_signal_6247, MixColumnsIns_n27}), .c ({new_AGEMA_signal_6945, new_AGEMA_signal_6944, new_AGEMA_signal_6943, MixColumnsOutput[1]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U45 ( .a ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, new_AGEMA_signal_5962, KeyExpansionIns_tmp[9]}), .b ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, new_AGEMA_signal_6064, MixColumnsIns_DoubleBytes[25]}), .c ({new_AGEMA_signal_6249, new_AGEMA_signal_6248, new_AGEMA_signal_6247, MixColumnsIns_n27}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U44 ( .a ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, KeyExpansionIns_tmp[17]}), .b ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, new_AGEMA_signal_6250, MixColumnsIns_n62}), .c ({new_AGEMA_signal_6546, new_AGEMA_signal_6545, new_AGEMA_signal_6544, MixColumnsIns_n14}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U43 ( .a ({new_AGEMA_signal_5985, new_AGEMA_signal_5984, new_AGEMA_signal_5983, KeyExpansionIns_tmp[1]}), .b ({new_AGEMA_signal_6093, new_AGEMA_signal_6092, new_AGEMA_signal_6091, MixColumnsIns_DoubleBytes[1]}), .c ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, new_AGEMA_signal_6250, MixColumnsIns_n62}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U42 ( .a ({new_AGEMA_signal_6549, new_AGEMA_signal_6548, new_AGEMA_signal_6547, MixColumnsIns_n13}), .b ({new_AGEMA_signal_6255, new_AGEMA_signal_6254, new_AGEMA_signal_6253, MixColumnsIns_n31}), .c ({new_AGEMA_signal_6948, new_AGEMA_signal_6947, new_AGEMA_signal_6946, MixColumnsOutput[19]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U41 ( .a ({new_AGEMA_signal_5937, new_AGEMA_signal_5936, new_AGEMA_signal_5935, KeyExpansionIns_tmp[19]}), .b ({new_AGEMA_signal_6072, new_AGEMA_signal_6071, new_AGEMA_signal_6070, MixColumnsIns_DoubleBytes[19]}), .c ({new_AGEMA_signal_6255, new_AGEMA_signal_6254, new_AGEMA_signal_6253, MixColumnsIns_n31}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U40 ( .a ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, new_AGEMA_signal_5977, KeyExpansionIns_tmp[3]}), .b ({new_AGEMA_signal_6285, new_AGEMA_signal_6284, new_AGEMA_signal_6283, MixColumnsIns_n12}), .c ({new_AGEMA_signal_6549, new_AGEMA_signal_6548, new_AGEMA_signal_6547, MixColumnsIns_n13}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U39 ( .a ({new_AGEMA_signal_6258, new_AGEMA_signal_6257, new_AGEMA_signal_6256, MixColumnsIns_n11}), .b ({new_AGEMA_signal_6021, new_AGEMA_signal_6020, new_AGEMA_signal_6019, MixColumnsIns_n29}), .c ({new_AGEMA_signal_6552, new_AGEMA_signal_6551, new_AGEMA_signal_6550, MixColumnsOutput[18]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U38 ( .a ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, new_AGEMA_signal_5938, KeyExpansionIns_tmp[18]}), .b ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, new_AGEMA_signal_5962, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_6021, new_AGEMA_signal_6020, new_AGEMA_signal_6019, MixColumnsIns_n29}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U37 ( .a ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, new_AGEMA_signal_5980, KeyExpansionIns_tmp[2]}), .b ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, new_AGEMA_signal_6046, MixColumnsIns_n10}), .c ({new_AGEMA_signal_6258, new_AGEMA_signal_6257, new_AGEMA_signal_6256, MixColumnsIns_n11}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U36 ( .a ({new_AGEMA_signal_6555, new_AGEMA_signal_6554, new_AGEMA_signal_6553, MixColumnsIns_n9}), .b ({new_AGEMA_signal_6261, new_AGEMA_signal_6260, new_AGEMA_signal_6259, MixColumnsIns_n26}), .c ({new_AGEMA_signal_6951, new_AGEMA_signal_6950, new_AGEMA_signal_6949, MixColumnsOutput[17]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U35 ( .a ({new_AGEMA_signal_6075, new_AGEMA_signal_6074, new_AGEMA_signal_6073, MixColumnsIns_DoubleBytes[17]}), .b ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_6261, new_AGEMA_signal_6260, new_AGEMA_signal_6259, MixColumnsIns_n26}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U34 ( .a ({new_AGEMA_signal_6264, new_AGEMA_signal_6263, new_AGEMA_signal_6262, MixColumnsIns_n63}), .b ({new_AGEMA_signal_5985, new_AGEMA_signal_5984, new_AGEMA_signal_5983, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_6555, new_AGEMA_signal_6554, new_AGEMA_signal_6553, MixColumnsIns_n9}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U33 ( .a ({new_AGEMA_signal_6084, new_AGEMA_signal_6083, new_AGEMA_signal_6082, MixColumnsIns_DoubleBytes[9]}), .b ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, new_AGEMA_signal_5920, MixColumnsIns_DoubleBytes[2]}), .c ({new_AGEMA_signal_6264, new_AGEMA_signal_6263, new_AGEMA_signal_6262, MixColumnsIns_n63}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U32 ( .a ({new_AGEMA_signal_6267, new_AGEMA_signal_6266, new_AGEMA_signal_6265, MixColumnsIns_n8}), .b ({new_AGEMA_signal_6024, new_AGEMA_signal_6023, new_AGEMA_signal_6022, MixColumnsIns_n24}), .c ({new_AGEMA_signal_6558, new_AGEMA_signal_6557, new_AGEMA_signal_6556, MixColumnsOutput[16]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U31 ( .a ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, new_AGEMA_signal_5833, KeyExpansionIns_tmp[16]}), .b ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_6024, new_AGEMA_signal_6023, new_AGEMA_signal_6022, MixColumnsIns_n24}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U30 ( .a ({new_AGEMA_signal_5901, new_AGEMA_signal_5900, new_AGEMA_signal_5899, KeyExpansionIns_tmp[0]}), .b ({new_AGEMA_signal_6027, new_AGEMA_signal_6026, new_AGEMA_signal_6025, MixColumnsIns_n60}), .c ({new_AGEMA_signal_6267, new_AGEMA_signal_6266, new_AGEMA_signal_6265, MixColumnsIns_n8}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U29 ( .a ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, new_AGEMA_signal_5800, SubBytesOutput[0]}), .c ({new_AGEMA_signal_6027, new_AGEMA_signal_6026, new_AGEMA_signal_6025, MixColumnsIns_n60}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U28 ( .a ({new_AGEMA_signal_6270, new_AGEMA_signal_6269, new_AGEMA_signal_6268, MixColumnsIns_n7}), .b ({new_AGEMA_signal_6030, new_AGEMA_signal_6029, new_AGEMA_signal_6028, MixColumnsIns_n21}), .c ({new_AGEMA_signal_6561, new_AGEMA_signal_6560, new_AGEMA_signal_6559, MixColumnsOutput[15]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U27 ( .a ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, new_AGEMA_signal_5902, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, new_AGEMA_signal_5926, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_6030, new_AGEMA_signal_6029, new_AGEMA_signal_6028, MixColumnsIns_n21}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U26 ( .a ({new_AGEMA_signal_6033, new_AGEMA_signal_6032, new_AGEMA_signal_6031, MixColumnsIns_n56}), .b ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_6270, new_AGEMA_signal_6269, new_AGEMA_signal_6268, MixColumnsIns_n7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U25 ( .a ({new_AGEMA_signal_5907, new_AGEMA_signal_5906, new_AGEMA_signal_5905, MixColumnsIns_DoubleBytes[7]}), .b ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, new_AGEMA_signal_5965, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_6033, new_AGEMA_signal_6032, new_AGEMA_signal_6031, MixColumnsIns_n56}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U24 ( .a ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, new_AGEMA_signal_6271, MixColumnsIns_n6}), .b ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, new_AGEMA_signal_6034, MixColumnsIns_n19}), .c ({new_AGEMA_signal_6564, new_AGEMA_signal_6563, new_AGEMA_signal_6562, MixColumnsOutput[14]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U23 ( .a ({new_AGEMA_signal_5907, new_AGEMA_signal_5906, new_AGEMA_signal_5905, MixColumnsIns_DoubleBytes[7]}), .b ({new_AGEMA_signal_5931, new_AGEMA_signal_5930, new_AGEMA_signal_5929, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, new_AGEMA_signal_6034, MixColumnsIns_n19}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U22 ( .a ({new_AGEMA_signal_6039, new_AGEMA_signal_6038, new_AGEMA_signal_6037, MixColumnsIns_n53}), .b ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, new_AGEMA_signal_5947, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, new_AGEMA_signal_6271, MixColumnsIns_n6}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U21 ( .a ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, new_AGEMA_signal_5908, MixColumnsIns_DoubleBytes[6]}), .b ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, new_AGEMA_signal_5968, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_6039, new_AGEMA_signal_6038, new_AGEMA_signal_6037, MixColumnsIns_n53}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U20 ( .a ({new_AGEMA_signal_6276, new_AGEMA_signal_6275, new_AGEMA_signal_6274, MixColumnsIns_n5}), .b ({new_AGEMA_signal_6042, new_AGEMA_signal_6041, new_AGEMA_signal_6040, MixColumnsIns_n17}), .c ({new_AGEMA_signal_6567, new_AGEMA_signal_6566, new_AGEMA_signal_6565, MixColumnsOutput[13]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U19 ( .a ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, new_AGEMA_signal_5908, MixColumnsIns_DoubleBytes[6]}), .b ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, new_AGEMA_signal_5932, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_6042, new_AGEMA_signal_6041, new_AGEMA_signal_6040, MixColumnsIns_n17}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U18 ( .a ({new_AGEMA_signal_6045, new_AGEMA_signal_6044, new_AGEMA_signal_6043, MixColumnsIns_n50}), .b ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, new_AGEMA_signal_5950, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_6276, new_AGEMA_signal_6275, new_AGEMA_signal_6274, MixColumnsIns_n5}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U17 ( .a ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, MixColumnsIns_DoubleBytes[5]}), .b ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_6045, new_AGEMA_signal_6044, new_AGEMA_signal_6043, MixColumnsIns_n50}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U16 ( .a ({new_AGEMA_signal_6570, new_AGEMA_signal_6569, new_AGEMA_signal_6568, MixColumnsIns_n4}), .b ({new_AGEMA_signal_6279, new_AGEMA_signal_6278, new_AGEMA_signal_6277, MixColumnsIns_n15}), .c ({new_AGEMA_signal_6954, new_AGEMA_signal_6953, new_AGEMA_signal_6952, MixColumnsOutput[12]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U15 ( .a ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, MixColumnsIns_DoubleBytes[5]}), .b ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, new_AGEMA_signal_6076, MixColumnsIns_DoubleBytes[12]}), .c ({new_AGEMA_signal_6279, new_AGEMA_signal_6278, new_AGEMA_signal_6277, MixColumnsIns_n15}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U14 ( .a ({new_AGEMA_signal_6282, new_AGEMA_signal_6281, new_AGEMA_signal_6280, MixColumnsIns_n47}), .b ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, new_AGEMA_signal_5953, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_6570, new_AGEMA_signal_6569, new_AGEMA_signal_6568, MixColumnsIns_n4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U13 ( .a ({new_AGEMA_signal_6087, new_AGEMA_signal_6086, new_AGEMA_signal_6085, MixColumnsIns_DoubleBytes[4]}), .b ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, new_AGEMA_signal_5974, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_6282, new_AGEMA_signal_6281, new_AGEMA_signal_6280, MixColumnsIns_n47}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U12 ( .a ({new_AGEMA_signal_6573, new_AGEMA_signal_6572, new_AGEMA_signal_6571, MixColumnsIns_n3}), .b ({new_AGEMA_signal_6285, new_AGEMA_signal_6284, new_AGEMA_signal_6283, MixColumnsIns_n12}), .c ({new_AGEMA_signal_6957, new_AGEMA_signal_6956, new_AGEMA_signal_6955, MixColumnsOutput[11]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U11 ( .a ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, new_AGEMA_signal_5914, SubBytesOutput[3]}), .b ({new_AGEMA_signal_6081, new_AGEMA_signal_6080, new_AGEMA_signal_6079, MixColumnsIns_DoubleBytes[11]}), .c ({new_AGEMA_signal_6285, new_AGEMA_signal_6284, new_AGEMA_signal_6283, MixColumnsIns_n12}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U10 ( .a ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, new_AGEMA_signal_6286, MixColumnsIns_n44}), .b ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, new_AGEMA_signal_5956, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_6573, new_AGEMA_signal_6572, new_AGEMA_signal_6571, MixColumnsIns_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U9 ( .a ({new_AGEMA_signal_6090, new_AGEMA_signal_6089, new_AGEMA_signal_6088, MixColumnsIns_DoubleBytes[3]}), .b ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, new_AGEMA_signal_5977, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, new_AGEMA_signal_6286, MixColumnsIns_n44}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U8 ( .a ({new_AGEMA_signal_6291, new_AGEMA_signal_6290, new_AGEMA_signal_6289, MixColumnsIns_n2}), .b ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, new_AGEMA_signal_6046, MixColumnsIns_n10}), .c ({new_AGEMA_signal_6576, new_AGEMA_signal_6575, new_AGEMA_signal_6574, MixColumnsOutput[10]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U7 ( .a ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesOutput[2]}), .b ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, new_AGEMA_signal_6046, MixColumnsIns_n10}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U6 ( .a ({new_AGEMA_signal_6051, new_AGEMA_signal_6050, new_AGEMA_signal_6049, MixColumnsIns_n37}), .b ({new_AGEMA_signal_5961, new_AGEMA_signal_5960, new_AGEMA_signal_5959, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_6291, new_AGEMA_signal_6290, new_AGEMA_signal_6289, MixColumnsIns_n2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U5 ( .a ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, new_AGEMA_signal_5920, MixColumnsIns_DoubleBytes[2]}), .b ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, new_AGEMA_signal_5980, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_6051, new_AGEMA_signal_6050, new_AGEMA_signal_6049, MixColumnsIns_n37}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U4 ( .a ({new_AGEMA_signal_6294, new_AGEMA_signal_6293, new_AGEMA_signal_6292, MixColumnsIns_n1}), .b ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, new_AGEMA_signal_5833, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_6579, new_AGEMA_signal_6578, new_AGEMA_signal_6577, MixColumnsOutput[0]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U3 ( .a ({new_AGEMA_signal_6057, new_AGEMA_signal_6056, new_AGEMA_signal_6055, MixColumnsIns_n59}), .b ({new_AGEMA_signal_6054, new_AGEMA_signal_6053, new_AGEMA_signal_6052, MixColumnsIns_n23}), .c ({new_AGEMA_signal_6294, new_AGEMA_signal_6293, new_AGEMA_signal_6292, MixColumnsIns_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U2 ( .a ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, new_AGEMA_signal_5866, KeyExpansionIns_tmp[8]}), .b ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, new_AGEMA_signal_5965, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_6054, new_AGEMA_signal_6053, new_AGEMA_signal_6052, MixColumnsIns_n23}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_U1 ( .a ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, new_AGEMA_signal_5902, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_5901, new_AGEMA_signal_5900, new_AGEMA_signal_5899, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_6057, new_AGEMA_signal_6056, new_AGEMA_signal_6055, MixColumnsIns_n59}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, new_AGEMA_signal_5965, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, new_AGEMA_signal_5977, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_6060, new_AGEMA_signal_6059, new_AGEMA_signal_6058, MixColumnsIns_DoubleBytes[28]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, new_AGEMA_signal_5965, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, new_AGEMA_signal_5980, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, new_AGEMA_signal_6061, MixColumnsIns_DoubleBytes[27]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, new_AGEMA_signal_5965, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_5901, new_AGEMA_signal_5900, new_AGEMA_signal_5899, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, new_AGEMA_signal_6064, MixColumnsIns_DoubleBytes[25]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, new_AGEMA_signal_5956, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_6069, new_AGEMA_signal_6068, new_AGEMA_signal_6067, MixColumnsIns_DoubleBytes[20]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_5961, new_AGEMA_signal_5960, new_AGEMA_signal_5959, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_6072, new_AGEMA_signal_6071, new_AGEMA_signal_6070, MixColumnsIns_DoubleBytes[19]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, new_AGEMA_signal_5866, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_6075, new_AGEMA_signal_6074, new_AGEMA_signal_6073, MixColumnsIns_DoubleBytes[17]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_5937, new_AGEMA_signal_5936, new_AGEMA_signal_5935, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, new_AGEMA_signal_6076, MixColumnsIns_DoubleBytes[12]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, new_AGEMA_signal_5938, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_6081, new_AGEMA_signal_6080, new_AGEMA_signal_6079, MixColumnsIns_DoubleBytes[11]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, new_AGEMA_signal_5833, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_6084, new_AGEMA_signal_6083, new_AGEMA_signal_6082, MixColumnsIns_DoubleBytes[9]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, new_AGEMA_signal_5902, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, new_AGEMA_signal_5914, SubBytesOutput[3]}), .c ({new_AGEMA_signal_6087, new_AGEMA_signal_6086, new_AGEMA_signal_6085, MixColumnsIns_DoubleBytes[4]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, new_AGEMA_signal_5902, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesOutput[2]}), .c ({new_AGEMA_signal_6090, new_AGEMA_signal_6089, new_AGEMA_signal_6088, MixColumnsIns_DoubleBytes[3]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) MixColumnsIns_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, new_AGEMA_signal_5902, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, new_AGEMA_signal_5800, SubBytesOutput[0]}), .c ({new_AGEMA_signal_6093, new_AGEMA_signal_6092, new_AGEMA_signal_6091, MixColumnsIns_DoubleBytes[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_0_U1 ( .s (new_AGEMA_signal_11461), .b ({new_AGEMA_signal_6579, new_AGEMA_signal_6578, new_AGEMA_signal_6577, MixColumnsOutput[0]}), .a ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, new_AGEMA_signal_5800, SubBytesOutput[0]}), .c ({new_AGEMA_signal_6960, new_AGEMA_signal_6959, new_AGEMA_signal_6958, ColumnOutput[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_1_U1 ( .s (new_AGEMA_signal_11465), .b ({new_AGEMA_signal_6945, new_AGEMA_signal_6944, new_AGEMA_signal_6943, MixColumnsOutput[1]}), .a ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, new_AGEMA_signal_5920, MixColumnsIns_DoubleBytes[2]}), .c ({new_AGEMA_signal_7395, new_AGEMA_signal_7394, new_AGEMA_signal_7393, ColumnOutput[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_2_U1 ( .s (new_AGEMA_signal_11465), .b ({new_AGEMA_signal_6513, new_AGEMA_signal_6512, new_AGEMA_signal_6511, MixColumnsOutput[2]}), .a ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesOutput[2]}), .c ({new_AGEMA_signal_6963, new_AGEMA_signal_6962, new_AGEMA_signal_6961, ColumnOutput[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_3_U1 ( .s (new_AGEMA_signal_11465), .b ({new_AGEMA_signal_6930, new_AGEMA_signal_6929, new_AGEMA_signal_6928, MixColumnsOutput[3]}), .a ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, new_AGEMA_signal_5914, SubBytesOutput[3]}), .c ({new_AGEMA_signal_7398, new_AGEMA_signal_7397, new_AGEMA_signal_7396, ColumnOutput[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_4_U1 ( .s (new_AGEMA_signal_11465), .b ({new_AGEMA_signal_6927, new_AGEMA_signal_6926, new_AGEMA_signal_6925, MixColumnsOutput[4]}), .a ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, MixColumnsIns_DoubleBytes[5]}), .c ({new_AGEMA_signal_7401, new_AGEMA_signal_7400, new_AGEMA_signal_7399, ColumnOutput[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_5_U1 ( .s (new_AGEMA_signal_11465), .b ({new_AGEMA_signal_6498, new_AGEMA_signal_6497, new_AGEMA_signal_6496, MixColumnsOutput[5]}), .a ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, new_AGEMA_signal_5908, MixColumnsIns_DoubleBytes[6]}), .c ({new_AGEMA_signal_6966, new_AGEMA_signal_6965, new_AGEMA_signal_6964, ColumnOutput[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_6_U1 ( .s (new_AGEMA_signal_11465), .b ({new_AGEMA_signal_6495, new_AGEMA_signal_6494, new_AGEMA_signal_6493, MixColumnsOutput[6]}), .a ({new_AGEMA_signal_5907, new_AGEMA_signal_5906, new_AGEMA_signal_5905, MixColumnsIns_DoubleBytes[7]}), .c ({new_AGEMA_signal_6969, new_AGEMA_signal_6968, new_AGEMA_signal_6967, ColumnOutput[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_7_U1 ( .s (new_AGEMA_signal_11469), .b ({new_AGEMA_signal_6492, new_AGEMA_signal_6491, new_AGEMA_signal_6490, MixColumnsOutput[7]}), .a ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, new_AGEMA_signal_5902, MixColumnsIns_DoubleBytes[0]}), .c ({new_AGEMA_signal_6972, new_AGEMA_signal_6971, new_AGEMA_signal_6970, ColumnOutput[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_8_U1 ( .s (new_AGEMA_signal_11461), .b ({new_AGEMA_signal_6489, new_AGEMA_signal_6488, new_AGEMA_signal_6487, MixColumnsOutput[8]}), .a ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, new_AGEMA_signal_5833, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_6975, new_AGEMA_signal_6974, new_AGEMA_signal_6973, ColumnOutput[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_9_U1 ( .s (new_AGEMA_signal_11461), .b ({new_AGEMA_signal_6924, new_AGEMA_signal_6923, new_AGEMA_signal_6922, MixColumnsOutput[9]}), .a ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_7404, new_AGEMA_signal_7403, new_AGEMA_signal_7402, ColumnOutput[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_10_U1 ( .s (new_AGEMA_signal_11461), .b ({new_AGEMA_signal_6576, new_AGEMA_signal_6575, new_AGEMA_signal_6574, MixColumnsOutput[10]}), .a ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, new_AGEMA_signal_5938, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_6978, new_AGEMA_signal_6977, new_AGEMA_signal_6976, ColumnOutput[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_11_U1 ( .s (new_AGEMA_signal_11461), .b ({new_AGEMA_signal_6957, new_AGEMA_signal_6956, new_AGEMA_signal_6955, MixColumnsOutput[11]}), .a ({new_AGEMA_signal_5937, new_AGEMA_signal_5936, new_AGEMA_signal_5935, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_7407, new_AGEMA_signal_7406, new_AGEMA_signal_7405, ColumnOutput[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_12_U1 ( .s (new_AGEMA_signal_11461), .b ({new_AGEMA_signal_6954, new_AGEMA_signal_6953, new_AGEMA_signal_6952, MixColumnsOutput[12]}), .a ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, new_AGEMA_signal_5932, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_7410, new_AGEMA_signal_7409, new_AGEMA_signal_7408, ColumnOutput[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_13_U1 ( .s (new_AGEMA_signal_11461), .b ({new_AGEMA_signal_6567, new_AGEMA_signal_6566, new_AGEMA_signal_6565, MixColumnsOutput[13]}), .a ({new_AGEMA_signal_5931, new_AGEMA_signal_5930, new_AGEMA_signal_5929, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_6981, new_AGEMA_signal_6980, new_AGEMA_signal_6979, ColumnOutput[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_14_U1 ( .s (new_AGEMA_signal_11461), .b ({new_AGEMA_signal_6564, new_AGEMA_signal_6563, new_AGEMA_signal_6562, MixColumnsOutput[14]}), .a ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, new_AGEMA_signal_5926, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_6984, new_AGEMA_signal_6983, new_AGEMA_signal_6982, ColumnOutput[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_15_U1 ( .s (new_AGEMA_signal_11461), .b ({new_AGEMA_signal_6561, new_AGEMA_signal_6560, new_AGEMA_signal_6559, MixColumnsOutput[15]}), .a ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_6987, new_AGEMA_signal_6986, new_AGEMA_signal_6985, ColumnOutput[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_16_U1 ( .s (new_AGEMA_signal_11461), .b ({new_AGEMA_signal_6558, new_AGEMA_signal_6557, new_AGEMA_signal_6556, MixColumnsOutput[16]}), .a ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, new_AGEMA_signal_5866, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_6990, new_AGEMA_signal_6989, new_AGEMA_signal_6988, ColumnOutput[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_17_U1 ( .s (new_AGEMA_signal_11461), .b ({new_AGEMA_signal_6951, new_AGEMA_signal_6950, new_AGEMA_signal_6949, MixColumnsOutput[17]}), .a ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, new_AGEMA_signal_5962, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_7413, new_AGEMA_signal_7412, new_AGEMA_signal_7411, ColumnOutput[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_18_U1 ( .s (new_AGEMA_signal_11461), .b ({new_AGEMA_signal_6552, new_AGEMA_signal_6551, new_AGEMA_signal_6550, MixColumnsOutput[18]}), .a ({new_AGEMA_signal_5961, new_AGEMA_signal_5960, new_AGEMA_signal_5959, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_6993, new_AGEMA_signal_6992, new_AGEMA_signal_6991, ColumnOutput[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_19_U1 ( .s (new_AGEMA_signal_11461), .b ({new_AGEMA_signal_6948, new_AGEMA_signal_6947, new_AGEMA_signal_6946, MixColumnsOutput[19]}), .a ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, new_AGEMA_signal_5956, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, new_AGEMA_signal_7414, ColumnOutput[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_20_U1 ( .s (new_AGEMA_signal_11469), .b ({new_AGEMA_signal_6942, new_AGEMA_signal_6941, new_AGEMA_signal_6940, MixColumnsOutput[20]}), .a ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, new_AGEMA_signal_5953, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_7419, new_AGEMA_signal_7418, new_AGEMA_signal_7417, ColumnOutput[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_21_U1 ( .s (new_AGEMA_signal_11469), .b ({new_AGEMA_signal_6540, new_AGEMA_signal_6539, new_AGEMA_signal_6538, MixColumnsOutput[21]}), .a ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, new_AGEMA_signal_5950, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_6996, new_AGEMA_signal_6995, new_AGEMA_signal_6994, ColumnOutput[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_22_U1 ( .s (new_AGEMA_signal_11469), .b ({new_AGEMA_signal_6537, new_AGEMA_signal_6536, new_AGEMA_signal_6535, MixColumnsOutput[22]}), .a ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, new_AGEMA_signal_5947, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_6999, new_AGEMA_signal_6998, new_AGEMA_signal_6997, ColumnOutput[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_23_U1 ( .s (new_AGEMA_signal_11469), .b ({new_AGEMA_signal_6534, new_AGEMA_signal_6533, new_AGEMA_signal_6532, MixColumnsOutput[23]}), .a ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_7002, new_AGEMA_signal_7001, new_AGEMA_signal_7000, ColumnOutput[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_24_U1 ( .s (new_AGEMA_signal_11469), .b ({new_AGEMA_signal_6531, new_AGEMA_signal_6530, new_AGEMA_signal_6529, MixColumnsOutput[24]}), .a ({new_AGEMA_signal_5901, new_AGEMA_signal_5900, new_AGEMA_signal_5899, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_7005, new_AGEMA_signal_7004, new_AGEMA_signal_7003, ColumnOutput[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_25_U1 ( .s (new_AGEMA_signal_11469), .b ({new_AGEMA_signal_6939, new_AGEMA_signal_6938, new_AGEMA_signal_6937, MixColumnsOutput[25]}), .a ({new_AGEMA_signal_5985, new_AGEMA_signal_5984, new_AGEMA_signal_5983, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_7422, new_AGEMA_signal_7421, new_AGEMA_signal_7420, ColumnOutput[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_26_U1 ( .s (new_AGEMA_signal_11469), .b ({new_AGEMA_signal_6525, new_AGEMA_signal_6524, new_AGEMA_signal_6523, MixColumnsOutput[26]}), .a ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, new_AGEMA_signal_5980, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_7008, new_AGEMA_signal_7007, new_AGEMA_signal_7006, ColumnOutput[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_27_U1 ( .s (new_AGEMA_signal_11469), .b ({new_AGEMA_signal_6936, new_AGEMA_signal_6935, new_AGEMA_signal_6934, MixColumnsOutput[27]}), .a ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, new_AGEMA_signal_5977, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_7425, new_AGEMA_signal_7424, new_AGEMA_signal_7423, ColumnOutput[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_28_U1 ( .s (new_AGEMA_signal_11469), .b ({new_AGEMA_signal_6933, new_AGEMA_signal_6932, new_AGEMA_signal_6931, MixColumnsOutput[28]}), .a ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, new_AGEMA_signal_5974, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_7428, new_AGEMA_signal_7427, new_AGEMA_signal_7426, ColumnOutput[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_29_U1 ( .s (new_AGEMA_signal_11469), .b ({new_AGEMA_signal_6516, new_AGEMA_signal_6515, new_AGEMA_signal_6514, MixColumnsOutput[29]}), .a ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_7011, new_AGEMA_signal_7010, new_AGEMA_signal_7009, ColumnOutput[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_30_U1 ( .s (new_AGEMA_signal_11469), .b ({new_AGEMA_signal_6510, new_AGEMA_signal_6509, new_AGEMA_signal_6508, MixColumnsOutput[30]}), .a ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, new_AGEMA_signal_5968, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_7014, new_AGEMA_signal_7013, new_AGEMA_signal_7012, ColumnOutput[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxMCOut_mux_inst_31_U1 ( .s (new_AGEMA_signal_11469), .b ({new_AGEMA_signal_6507, new_AGEMA_signal_6506, new_AGEMA_signal_6505, MixColumnsOutput[31]}), .a ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, new_AGEMA_signal_5965, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_7017, new_AGEMA_signal_7016, new_AGEMA_signal_7015, ColumnOutput[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_0_U1 ( .s (new_AGEMA_signal_11473), .b ({new_AGEMA_signal_6960, new_AGEMA_signal_6959, new_AGEMA_signal_6958, ColumnOutput[0]}), .a ({new_AGEMA_signal_11489, new_AGEMA_signal_11485, new_AGEMA_signal_11481, new_AGEMA_signal_11477}), .c ({new_AGEMA_signal_7431, new_AGEMA_signal_7430, new_AGEMA_signal_7429, RoundOutput[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_1_U1 ( .s (new_AGEMA_signal_11493), .b ({new_AGEMA_signal_7395, new_AGEMA_signal_7394, new_AGEMA_signal_7393, ColumnOutput[1]}), .a ({new_AGEMA_signal_11509, new_AGEMA_signal_11505, new_AGEMA_signal_11501, new_AGEMA_signal_11497}), .c ({new_AGEMA_signal_7911, new_AGEMA_signal_7910, new_AGEMA_signal_7909, RoundOutput[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_2_U1 ( .s (new_AGEMA_signal_11513), .b ({new_AGEMA_signal_6963, new_AGEMA_signal_6962, new_AGEMA_signal_6961, ColumnOutput[2]}), .a ({new_AGEMA_signal_11529, new_AGEMA_signal_11525, new_AGEMA_signal_11521, new_AGEMA_signal_11517}), .c ({new_AGEMA_signal_7434, new_AGEMA_signal_7433, new_AGEMA_signal_7432, RoundOutput[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_3_U1 ( .s (new_AGEMA_signal_11533), .b ({new_AGEMA_signal_7398, new_AGEMA_signal_7397, new_AGEMA_signal_7396, ColumnOutput[3]}), .a ({new_AGEMA_signal_11549, new_AGEMA_signal_11545, new_AGEMA_signal_11541, new_AGEMA_signal_11537}), .c ({new_AGEMA_signal_7914, new_AGEMA_signal_7913, new_AGEMA_signal_7912, RoundOutput[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_4_U1 ( .s (new_AGEMA_signal_11553), .b ({new_AGEMA_signal_7401, new_AGEMA_signal_7400, new_AGEMA_signal_7399, ColumnOutput[4]}), .a ({new_AGEMA_signal_11569, new_AGEMA_signal_11565, new_AGEMA_signal_11561, new_AGEMA_signal_11557}), .c ({new_AGEMA_signal_7917, new_AGEMA_signal_7916, new_AGEMA_signal_7915, RoundOutput[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_5_U1 ( .s (new_AGEMA_signal_11573), .b ({new_AGEMA_signal_6966, new_AGEMA_signal_6965, new_AGEMA_signal_6964, ColumnOutput[5]}), .a ({new_AGEMA_signal_11589, new_AGEMA_signal_11585, new_AGEMA_signal_11581, new_AGEMA_signal_11577}), .c ({new_AGEMA_signal_7437, new_AGEMA_signal_7436, new_AGEMA_signal_7435, RoundOutput[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_6_U1 ( .s (new_AGEMA_signal_11593), .b ({new_AGEMA_signal_6969, new_AGEMA_signal_6968, new_AGEMA_signal_6967, ColumnOutput[6]}), .a ({new_AGEMA_signal_11609, new_AGEMA_signal_11605, new_AGEMA_signal_11601, new_AGEMA_signal_11597}), .c ({new_AGEMA_signal_7440, new_AGEMA_signal_7439, new_AGEMA_signal_7438, RoundOutput[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_7_U1 ( .s (new_AGEMA_signal_11493), .b ({new_AGEMA_signal_6972, new_AGEMA_signal_6971, new_AGEMA_signal_6970, ColumnOutput[7]}), .a ({new_AGEMA_signal_11625, new_AGEMA_signal_11621, new_AGEMA_signal_11617, new_AGEMA_signal_11613}), .c ({new_AGEMA_signal_7443, new_AGEMA_signal_7442, new_AGEMA_signal_7441, RoundOutput[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_8_U1 ( .s (new_AGEMA_signal_11553), .b ({new_AGEMA_signal_6975, new_AGEMA_signal_6974, new_AGEMA_signal_6973, ColumnOutput[8]}), .a ({new_AGEMA_signal_11641, new_AGEMA_signal_11637, new_AGEMA_signal_11633, new_AGEMA_signal_11629}), .c ({new_AGEMA_signal_7446, new_AGEMA_signal_7445, new_AGEMA_signal_7444, RoundOutput[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_9_U1 ( .s (new_AGEMA_signal_11493), .b ({new_AGEMA_signal_7404, new_AGEMA_signal_7403, new_AGEMA_signal_7402, ColumnOutput[9]}), .a ({new_AGEMA_signal_11657, new_AGEMA_signal_11653, new_AGEMA_signal_11649, new_AGEMA_signal_11645}), .c ({new_AGEMA_signal_7920, new_AGEMA_signal_7919, new_AGEMA_signal_7918, RoundOutput[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_10_U1 ( .s (new_AGEMA_signal_11473), .b ({new_AGEMA_signal_6978, new_AGEMA_signal_6977, new_AGEMA_signal_6976, ColumnOutput[10]}), .a ({new_AGEMA_signal_11673, new_AGEMA_signal_11669, new_AGEMA_signal_11665, new_AGEMA_signal_11661}), .c ({new_AGEMA_signal_7449, new_AGEMA_signal_7448, new_AGEMA_signal_7447, RoundOutput[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_11_U1 ( .s (new_AGEMA_signal_11473), .b ({new_AGEMA_signal_7407, new_AGEMA_signal_7406, new_AGEMA_signal_7405, ColumnOutput[11]}), .a ({new_AGEMA_signal_11689, new_AGEMA_signal_11685, new_AGEMA_signal_11681, new_AGEMA_signal_11677}), .c ({new_AGEMA_signal_7923, new_AGEMA_signal_7922, new_AGEMA_signal_7921, RoundOutput[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_12_U1 ( .s (new_AGEMA_signal_11473), .b ({new_AGEMA_signal_7410, new_AGEMA_signal_7409, new_AGEMA_signal_7408, ColumnOutput[12]}), .a ({new_AGEMA_signal_11705, new_AGEMA_signal_11701, new_AGEMA_signal_11697, new_AGEMA_signal_11693}), .c ({new_AGEMA_signal_7926, new_AGEMA_signal_7925, new_AGEMA_signal_7924, RoundOutput[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_13_U1 ( .s (new_AGEMA_signal_11473), .b ({new_AGEMA_signal_6981, new_AGEMA_signal_6980, new_AGEMA_signal_6979, ColumnOutput[13]}), .a ({new_AGEMA_signal_11721, new_AGEMA_signal_11717, new_AGEMA_signal_11713, new_AGEMA_signal_11709}), .c ({new_AGEMA_signal_7452, new_AGEMA_signal_7451, new_AGEMA_signal_7450, RoundOutput[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_14_U1 ( .s (new_AGEMA_signal_11473), .b ({new_AGEMA_signal_6984, new_AGEMA_signal_6983, new_AGEMA_signal_6982, ColumnOutput[14]}), .a ({new_AGEMA_signal_11737, new_AGEMA_signal_11733, new_AGEMA_signal_11729, new_AGEMA_signal_11725}), .c ({new_AGEMA_signal_7455, new_AGEMA_signal_7454, new_AGEMA_signal_7453, RoundOutput[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_15_U1 ( .s (new_AGEMA_signal_11473), .b ({new_AGEMA_signal_6987, new_AGEMA_signal_6986, new_AGEMA_signal_6985, ColumnOutput[15]}), .a ({new_AGEMA_signal_11753, new_AGEMA_signal_11749, new_AGEMA_signal_11745, new_AGEMA_signal_11741}), .c ({new_AGEMA_signal_7458, new_AGEMA_signal_7457, new_AGEMA_signal_7456, RoundOutput[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_16_U1 ( .s (new_AGEMA_signal_11473), .b ({new_AGEMA_signal_6990, new_AGEMA_signal_6989, new_AGEMA_signal_6988, ColumnOutput[16]}), .a ({new_AGEMA_signal_11769, new_AGEMA_signal_11765, new_AGEMA_signal_11761, new_AGEMA_signal_11757}), .c ({new_AGEMA_signal_7461, new_AGEMA_signal_7460, new_AGEMA_signal_7459, RoundOutput[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_17_U1 ( .s (new_AGEMA_signal_11473), .b ({new_AGEMA_signal_7413, new_AGEMA_signal_7412, new_AGEMA_signal_7411, ColumnOutput[17]}), .a ({new_AGEMA_signal_11785, new_AGEMA_signal_11781, new_AGEMA_signal_11777, new_AGEMA_signal_11773}), .c ({new_AGEMA_signal_7929, new_AGEMA_signal_7928, new_AGEMA_signal_7927, RoundOutput[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_18_U1 ( .s (new_AGEMA_signal_11473), .b ({new_AGEMA_signal_6993, new_AGEMA_signal_6992, new_AGEMA_signal_6991, ColumnOutput[18]}), .a ({new_AGEMA_signal_11801, new_AGEMA_signal_11797, new_AGEMA_signal_11793, new_AGEMA_signal_11789}), .c ({new_AGEMA_signal_7464, new_AGEMA_signal_7463, new_AGEMA_signal_7462, RoundOutput[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_19_U1 ( .s (new_AGEMA_signal_11473), .b ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, new_AGEMA_signal_7414, ColumnOutput[19]}), .a ({new_AGEMA_signal_11817, new_AGEMA_signal_11813, new_AGEMA_signal_11809, new_AGEMA_signal_11805}), .c ({new_AGEMA_signal_7932, new_AGEMA_signal_7931, new_AGEMA_signal_7930, RoundOutput[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_20_U1 ( .s (new_AGEMA_signal_11513), .b ({new_AGEMA_signal_7419, new_AGEMA_signal_7418, new_AGEMA_signal_7417, ColumnOutput[20]}), .a ({new_AGEMA_signal_11833, new_AGEMA_signal_11829, new_AGEMA_signal_11825, new_AGEMA_signal_11821}), .c ({new_AGEMA_signal_7935, new_AGEMA_signal_7934, new_AGEMA_signal_7933, RoundOutput[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_21_U1 ( .s (new_AGEMA_signal_11533), .b ({new_AGEMA_signal_6996, new_AGEMA_signal_6995, new_AGEMA_signal_6994, ColumnOutput[21]}), .a ({new_AGEMA_signal_11849, new_AGEMA_signal_11845, new_AGEMA_signal_11841, new_AGEMA_signal_11837}), .c ({new_AGEMA_signal_7467, new_AGEMA_signal_7466, new_AGEMA_signal_7465, RoundOutput[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_22_U1 ( .s (new_AGEMA_signal_11553), .b ({new_AGEMA_signal_6999, new_AGEMA_signal_6998, new_AGEMA_signal_6997, ColumnOutput[22]}), .a ({new_AGEMA_signal_11865, new_AGEMA_signal_11861, new_AGEMA_signal_11857, new_AGEMA_signal_11853}), .c ({new_AGEMA_signal_7470, new_AGEMA_signal_7469, new_AGEMA_signal_7468, RoundOutput[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_23_U1 ( .s (new_AGEMA_signal_11573), .b ({new_AGEMA_signal_7002, new_AGEMA_signal_7001, new_AGEMA_signal_7000, ColumnOutput[23]}), .a ({new_AGEMA_signal_11881, new_AGEMA_signal_11877, new_AGEMA_signal_11873, new_AGEMA_signal_11869}), .c ({new_AGEMA_signal_7473, new_AGEMA_signal_7472, new_AGEMA_signal_7471, RoundOutput[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_24_U1 ( .s (new_AGEMA_signal_11593), .b ({new_AGEMA_signal_7005, new_AGEMA_signal_7004, new_AGEMA_signal_7003, ColumnOutput[24]}), .a ({new_AGEMA_signal_11897, new_AGEMA_signal_11893, new_AGEMA_signal_11889, new_AGEMA_signal_11885}), .c ({new_AGEMA_signal_7476, new_AGEMA_signal_7475, new_AGEMA_signal_7474, RoundOutput[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_25_U1 ( .s (new_AGEMA_signal_11553), .b ({new_AGEMA_signal_7422, new_AGEMA_signal_7421, new_AGEMA_signal_7420, ColumnOutput[25]}), .a ({new_AGEMA_signal_11913, new_AGEMA_signal_11909, new_AGEMA_signal_11905, new_AGEMA_signal_11901}), .c ({new_AGEMA_signal_7938, new_AGEMA_signal_7937, new_AGEMA_signal_7936, RoundOutput[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_26_U1 ( .s (new_AGEMA_signal_11573), .b ({new_AGEMA_signal_7008, new_AGEMA_signal_7007, new_AGEMA_signal_7006, ColumnOutput[26]}), .a ({new_AGEMA_signal_11929, new_AGEMA_signal_11925, new_AGEMA_signal_11921, new_AGEMA_signal_11917}), .c ({new_AGEMA_signal_7479, new_AGEMA_signal_7478, new_AGEMA_signal_7477, RoundOutput[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_27_U1 ( .s (new_AGEMA_signal_11473), .b ({new_AGEMA_signal_7425, new_AGEMA_signal_7424, new_AGEMA_signal_7423, ColumnOutput[27]}), .a ({new_AGEMA_signal_11945, new_AGEMA_signal_11941, new_AGEMA_signal_11937, new_AGEMA_signal_11933}), .c ({new_AGEMA_signal_7941, new_AGEMA_signal_7940, new_AGEMA_signal_7939, RoundOutput[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_28_U1 ( .s (new_AGEMA_signal_11473), .b ({new_AGEMA_signal_7428, new_AGEMA_signal_7427, new_AGEMA_signal_7426, ColumnOutput[28]}), .a ({new_AGEMA_signal_11961, new_AGEMA_signal_11957, new_AGEMA_signal_11953, new_AGEMA_signal_11949}), .c ({new_AGEMA_signal_7944, new_AGEMA_signal_7943, new_AGEMA_signal_7942, RoundOutput[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_29_U1 ( .s (new_AGEMA_signal_11493), .b ({new_AGEMA_signal_7011, new_AGEMA_signal_7010, new_AGEMA_signal_7009, ColumnOutput[29]}), .a ({new_AGEMA_signal_11977, new_AGEMA_signal_11973, new_AGEMA_signal_11969, new_AGEMA_signal_11965}), .c ({new_AGEMA_signal_7482, new_AGEMA_signal_7481, new_AGEMA_signal_7480, RoundOutput[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_30_U1 ( .s (new_AGEMA_signal_11513), .b ({new_AGEMA_signal_7014, new_AGEMA_signal_7013, new_AGEMA_signal_7012, ColumnOutput[30]}), .a ({new_AGEMA_signal_11993, new_AGEMA_signal_11989, new_AGEMA_signal_11985, new_AGEMA_signal_11981}), .c ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, new_AGEMA_signal_7483, RoundOutput[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxRound_mux_inst_31_U1 ( .s (new_AGEMA_signal_11533), .b ({new_AGEMA_signal_7017, new_AGEMA_signal_7016, new_AGEMA_signal_7015, ColumnOutput[31]}), .a ({new_AGEMA_signal_12009, new_AGEMA_signal_12005, new_AGEMA_signal_12001, new_AGEMA_signal_11997}), .c ({new_AGEMA_signal_7488, new_AGEMA_signal_7487, new_AGEMA_signal_7486, RoundOutput[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7299, new_AGEMA_signal_7298, new_AGEMA_signal_7297, RoundKeyOutput[0]}), .a ({new_AGEMA_signal_12025, new_AGEMA_signal_12021, new_AGEMA_signal_12017, new_AGEMA_signal_12013}), .c ({new_AGEMA_signal_7494, new_AGEMA_signal_7493, new_AGEMA_signal_7492, KeyReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7704, new_AGEMA_signal_7703, new_AGEMA_signal_7702, RoundKeyOutput[1]}), .a ({new_AGEMA_signal_12041, new_AGEMA_signal_12037, new_AGEMA_signal_12033, new_AGEMA_signal_12029}), .c ({new_AGEMA_signal_7950, new_AGEMA_signal_7949, new_AGEMA_signal_7948, KeyReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7707, new_AGEMA_signal_7706, new_AGEMA_signal_7705, RoundKeyOutput[2]}), .a ({new_AGEMA_signal_12057, new_AGEMA_signal_12053, new_AGEMA_signal_12049, new_AGEMA_signal_12045}), .c ({new_AGEMA_signal_7956, new_AGEMA_signal_7955, new_AGEMA_signal_7954, KeyReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7710, new_AGEMA_signal_7709, new_AGEMA_signal_7708, RoundKeyOutput[3]}), .a ({new_AGEMA_signal_12073, new_AGEMA_signal_12069, new_AGEMA_signal_12065, new_AGEMA_signal_12061}), .c ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, new_AGEMA_signal_7960, KeyReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7713, new_AGEMA_signal_7712, new_AGEMA_signal_7711, RoundKeyOutput[4]}), .a ({new_AGEMA_signal_12089, new_AGEMA_signal_12085, new_AGEMA_signal_12081, new_AGEMA_signal_12077}), .c ({new_AGEMA_signal_7968, new_AGEMA_signal_7967, new_AGEMA_signal_7966, KeyReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7716, new_AGEMA_signal_7715, new_AGEMA_signal_7714, RoundKeyOutput[5]}), .a ({new_AGEMA_signal_12105, new_AGEMA_signal_12101, new_AGEMA_signal_12097, new_AGEMA_signal_12093}), .c ({new_AGEMA_signal_7974, new_AGEMA_signal_7973, new_AGEMA_signal_7972, KeyReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7719, new_AGEMA_signal_7718, new_AGEMA_signal_7717, RoundKeyOutput[6]}), .a ({new_AGEMA_signal_12121, new_AGEMA_signal_12117, new_AGEMA_signal_12113, new_AGEMA_signal_12109}), .c ({new_AGEMA_signal_7980, new_AGEMA_signal_7979, new_AGEMA_signal_7978, KeyReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7722, new_AGEMA_signal_7721, new_AGEMA_signal_7720, RoundKeyOutput[7]}), .a ({new_AGEMA_signal_12137, new_AGEMA_signal_12133, new_AGEMA_signal_12129, new_AGEMA_signal_12125}), .c ({new_AGEMA_signal_7986, new_AGEMA_signal_7985, new_AGEMA_signal_7984, KeyReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, new_AGEMA_signal_7300, RoundKeyOutput[8]}), .a ({new_AGEMA_signal_12153, new_AGEMA_signal_12149, new_AGEMA_signal_12145, new_AGEMA_signal_12141}), .c ({new_AGEMA_signal_7500, new_AGEMA_signal_7499, new_AGEMA_signal_7498, KeyReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7725, new_AGEMA_signal_7724, new_AGEMA_signal_7723, RoundKeyOutput[9]}), .a ({new_AGEMA_signal_12169, new_AGEMA_signal_12165, new_AGEMA_signal_12161, new_AGEMA_signal_12157}), .c ({new_AGEMA_signal_7992, new_AGEMA_signal_7991, new_AGEMA_signal_7990, KeyReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7728, new_AGEMA_signal_7727, new_AGEMA_signal_7726, RoundKeyOutput[10]}), .a ({new_AGEMA_signal_12185, new_AGEMA_signal_12181, new_AGEMA_signal_12177, new_AGEMA_signal_12173}), .c ({new_AGEMA_signal_7998, new_AGEMA_signal_7997, new_AGEMA_signal_7996, KeyReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7731, new_AGEMA_signal_7730, new_AGEMA_signal_7729, RoundKeyOutput[11]}), .a ({new_AGEMA_signal_12201, new_AGEMA_signal_12197, new_AGEMA_signal_12193, new_AGEMA_signal_12189}), .c ({new_AGEMA_signal_8004, new_AGEMA_signal_8003, new_AGEMA_signal_8002, KeyReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7734, new_AGEMA_signal_7733, new_AGEMA_signal_7732, RoundKeyOutput[12]}), .a ({new_AGEMA_signal_12217, new_AGEMA_signal_12213, new_AGEMA_signal_12209, new_AGEMA_signal_12205}), .c ({new_AGEMA_signal_8010, new_AGEMA_signal_8009, new_AGEMA_signal_8008, KeyReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7737, new_AGEMA_signal_7736, new_AGEMA_signal_7735, RoundKeyOutput[13]}), .a ({new_AGEMA_signal_12233, new_AGEMA_signal_12229, new_AGEMA_signal_12225, new_AGEMA_signal_12221}), .c ({new_AGEMA_signal_8016, new_AGEMA_signal_8015, new_AGEMA_signal_8014, KeyReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7740, new_AGEMA_signal_7739, new_AGEMA_signal_7738, RoundKeyOutput[14]}), .a ({new_AGEMA_signal_12249, new_AGEMA_signal_12245, new_AGEMA_signal_12241, new_AGEMA_signal_12237}), .c ({new_AGEMA_signal_8022, new_AGEMA_signal_8021, new_AGEMA_signal_8020, KeyReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7743, new_AGEMA_signal_7742, new_AGEMA_signal_7741, RoundKeyOutput[15]}), .a ({new_AGEMA_signal_12265, new_AGEMA_signal_12261, new_AGEMA_signal_12257, new_AGEMA_signal_12253}), .c ({new_AGEMA_signal_8028, new_AGEMA_signal_8027, new_AGEMA_signal_8026, KeyReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7305, new_AGEMA_signal_7304, new_AGEMA_signal_7303, RoundKeyOutput[16]}), .a ({new_AGEMA_signal_12281, new_AGEMA_signal_12277, new_AGEMA_signal_12273, new_AGEMA_signal_12269}), .c ({new_AGEMA_signal_7506, new_AGEMA_signal_7505, new_AGEMA_signal_7504, KeyReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7746, new_AGEMA_signal_7745, new_AGEMA_signal_7744, RoundKeyOutput[17]}), .a ({new_AGEMA_signal_12297, new_AGEMA_signal_12293, new_AGEMA_signal_12289, new_AGEMA_signal_12285}), .c ({new_AGEMA_signal_8034, new_AGEMA_signal_8033, new_AGEMA_signal_8032, KeyReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7749, new_AGEMA_signal_7748, new_AGEMA_signal_7747, RoundKeyOutput[18]}), .a ({new_AGEMA_signal_12313, new_AGEMA_signal_12309, new_AGEMA_signal_12305, new_AGEMA_signal_12301}), .c ({new_AGEMA_signal_8040, new_AGEMA_signal_8039, new_AGEMA_signal_8038, KeyReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7752, new_AGEMA_signal_7751, new_AGEMA_signal_7750, RoundKeyOutput[19]}), .a ({new_AGEMA_signal_12329, new_AGEMA_signal_12325, new_AGEMA_signal_12321, new_AGEMA_signal_12317}), .c ({new_AGEMA_signal_8046, new_AGEMA_signal_8045, new_AGEMA_signal_8044, KeyReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7755, new_AGEMA_signal_7754, new_AGEMA_signal_7753, RoundKeyOutput[20]}), .a ({new_AGEMA_signal_12345, new_AGEMA_signal_12341, new_AGEMA_signal_12337, new_AGEMA_signal_12333}), .c ({new_AGEMA_signal_8052, new_AGEMA_signal_8051, new_AGEMA_signal_8050, KeyReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7758, new_AGEMA_signal_7757, new_AGEMA_signal_7756, RoundKeyOutput[21]}), .a ({new_AGEMA_signal_12361, new_AGEMA_signal_12357, new_AGEMA_signal_12353, new_AGEMA_signal_12349}), .c ({new_AGEMA_signal_8058, new_AGEMA_signal_8057, new_AGEMA_signal_8056, KeyReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7761, new_AGEMA_signal_7760, new_AGEMA_signal_7759, RoundKeyOutput[22]}), .a ({new_AGEMA_signal_12377, new_AGEMA_signal_12373, new_AGEMA_signal_12369, new_AGEMA_signal_12365}), .c ({new_AGEMA_signal_8064, new_AGEMA_signal_8063, new_AGEMA_signal_8062, KeyReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7764, new_AGEMA_signal_7763, new_AGEMA_signal_7762, RoundKeyOutput[23]}), .a ({new_AGEMA_signal_12393, new_AGEMA_signal_12389, new_AGEMA_signal_12385, new_AGEMA_signal_12381}), .c ({new_AGEMA_signal_8070, new_AGEMA_signal_8069, new_AGEMA_signal_8068, KeyReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7767, new_AGEMA_signal_7766, new_AGEMA_signal_7765, RoundKeyOutput[24]}), .a ({new_AGEMA_signal_12409, new_AGEMA_signal_12405, new_AGEMA_signal_12401, new_AGEMA_signal_12397}), .c ({new_AGEMA_signal_8076, new_AGEMA_signal_8075, new_AGEMA_signal_8074, KeyReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_8121, new_AGEMA_signal_8120, new_AGEMA_signal_8119, RoundKeyOutput[25]}), .a ({new_AGEMA_signal_12425, new_AGEMA_signal_12421, new_AGEMA_signal_12417, new_AGEMA_signal_12413}), .c ({new_AGEMA_signal_8217, new_AGEMA_signal_8216, new_AGEMA_signal_8215, KeyReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_8124, new_AGEMA_signal_8123, new_AGEMA_signal_8122, RoundKeyOutput[26]}), .a ({new_AGEMA_signal_12441, new_AGEMA_signal_12437, new_AGEMA_signal_12433, new_AGEMA_signal_12429}), .c ({new_AGEMA_signal_8223, new_AGEMA_signal_8222, new_AGEMA_signal_8221, KeyReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_8127, new_AGEMA_signal_8126, new_AGEMA_signal_8125, RoundKeyOutput[27]}), .a ({new_AGEMA_signal_12457, new_AGEMA_signal_12453, new_AGEMA_signal_12449, new_AGEMA_signal_12445}), .c ({new_AGEMA_signal_8229, new_AGEMA_signal_8228, new_AGEMA_signal_8227, KeyReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_8130, new_AGEMA_signal_8129, new_AGEMA_signal_8128, RoundKeyOutput[28]}), .a ({new_AGEMA_signal_12473, new_AGEMA_signal_12469, new_AGEMA_signal_12465, new_AGEMA_signal_12461}), .c ({new_AGEMA_signal_8235, new_AGEMA_signal_8234, new_AGEMA_signal_8233, KeyReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_8133, new_AGEMA_signal_8132, new_AGEMA_signal_8131, RoundKeyOutput[29]}), .a ({new_AGEMA_signal_12489, new_AGEMA_signal_12485, new_AGEMA_signal_12481, new_AGEMA_signal_12477}), .c ({new_AGEMA_signal_8241, new_AGEMA_signal_8240, new_AGEMA_signal_8239, KeyReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_8136, new_AGEMA_signal_8135, new_AGEMA_signal_8134, RoundKeyOutput[30]}), .a ({new_AGEMA_signal_12505, new_AGEMA_signal_12501, new_AGEMA_signal_12497, new_AGEMA_signal_12493}), .c ({new_AGEMA_signal_8247, new_AGEMA_signal_8246, new_AGEMA_signal_8245, KeyReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_8139, new_AGEMA_signal_8138, new_AGEMA_signal_8137, RoundKeyOutput[31]}), .a ({new_AGEMA_signal_12521, new_AGEMA_signal_12517, new_AGEMA_signal_12513, new_AGEMA_signal_12509}), .c ({new_AGEMA_signal_8253, new_AGEMA_signal_8252, new_AGEMA_signal_8251, KeyReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6828, new_AGEMA_signal_6827, new_AGEMA_signal_6826, RoundKeyOutput[32]}), .a ({new_AGEMA_signal_12537, new_AGEMA_signal_12533, new_AGEMA_signal_12529, new_AGEMA_signal_12525}), .c ({new_AGEMA_signal_7023, new_AGEMA_signal_7022, new_AGEMA_signal_7021, KeyReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7308, new_AGEMA_signal_7307, new_AGEMA_signal_7306, RoundKeyOutput[33]}), .a ({new_AGEMA_signal_12553, new_AGEMA_signal_12549, new_AGEMA_signal_12545, new_AGEMA_signal_12541}), .c ({new_AGEMA_signal_7512, new_AGEMA_signal_7511, new_AGEMA_signal_7510, KeyReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7311, new_AGEMA_signal_7310, new_AGEMA_signal_7309, RoundKeyOutput[34]}), .a ({new_AGEMA_signal_12569, new_AGEMA_signal_12565, new_AGEMA_signal_12561, new_AGEMA_signal_12557}), .c ({new_AGEMA_signal_7518, new_AGEMA_signal_7517, new_AGEMA_signal_7516, KeyReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7314, new_AGEMA_signal_7313, new_AGEMA_signal_7312, RoundKeyOutput[35]}), .a ({new_AGEMA_signal_12585, new_AGEMA_signal_12581, new_AGEMA_signal_12577, new_AGEMA_signal_12573}), .c ({new_AGEMA_signal_7524, new_AGEMA_signal_7523, new_AGEMA_signal_7522, KeyReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7317, new_AGEMA_signal_7316, new_AGEMA_signal_7315, RoundKeyOutput[36]}), .a ({new_AGEMA_signal_12601, new_AGEMA_signal_12597, new_AGEMA_signal_12593, new_AGEMA_signal_12589}), .c ({new_AGEMA_signal_7530, new_AGEMA_signal_7529, new_AGEMA_signal_7528, KeyReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7320, new_AGEMA_signal_7319, new_AGEMA_signal_7318, RoundKeyOutput[37]}), .a ({new_AGEMA_signal_12617, new_AGEMA_signal_12613, new_AGEMA_signal_12609, new_AGEMA_signal_12605}), .c ({new_AGEMA_signal_7536, new_AGEMA_signal_7535, new_AGEMA_signal_7534, KeyReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7323, new_AGEMA_signal_7322, new_AGEMA_signal_7321, RoundKeyOutput[38]}), .a ({new_AGEMA_signal_12633, new_AGEMA_signal_12629, new_AGEMA_signal_12625, new_AGEMA_signal_12621}), .c ({new_AGEMA_signal_7542, new_AGEMA_signal_7541, new_AGEMA_signal_7540, KeyReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7326, new_AGEMA_signal_7325, new_AGEMA_signal_7324, RoundKeyOutput[39]}), .a ({new_AGEMA_signal_12649, new_AGEMA_signal_12645, new_AGEMA_signal_12641, new_AGEMA_signal_12637}), .c ({new_AGEMA_signal_7548, new_AGEMA_signal_7547, new_AGEMA_signal_7546, KeyReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6831, new_AGEMA_signal_6830, new_AGEMA_signal_6829, RoundKeyOutput[40]}), .a ({new_AGEMA_signal_12665, new_AGEMA_signal_12661, new_AGEMA_signal_12657, new_AGEMA_signal_12653}), .c ({new_AGEMA_signal_7029, new_AGEMA_signal_7028, new_AGEMA_signal_7027, KeyReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7329, new_AGEMA_signal_7328, new_AGEMA_signal_7327, RoundKeyOutput[41]}), .a ({new_AGEMA_signal_12681, new_AGEMA_signal_12677, new_AGEMA_signal_12673, new_AGEMA_signal_12669}), .c ({new_AGEMA_signal_7554, new_AGEMA_signal_7553, new_AGEMA_signal_7552, KeyReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7332, new_AGEMA_signal_7331, new_AGEMA_signal_7330, RoundKeyOutput[42]}), .a ({new_AGEMA_signal_12697, new_AGEMA_signal_12693, new_AGEMA_signal_12689, new_AGEMA_signal_12685}), .c ({new_AGEMA_signal_7560, new_AGEMA_signal_7559, new_AGEMA_signal_7558, KeyReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7335, new_AGEMA_signal_7334, new_AGEMA_signal_7333, RoundKeyOutput[43]}), .a ({new_AGEMA_signal_12713, new_AGEMA_signal_12709, new_AGEMA_signal_12705, new_AGEMA_signal_12701}), .c ({new_AGEMA_signal_7566, new_AGEMA_signal_7565, new_AGEMA_signal_7564, KeyReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7338, new_AGEMA_signal_7337, new_AGEMA_signal_7336, RoundKeyOutput[44]}), .a ({new_AGEMA_signal_12729, new_AGEMA_signal_12725, new_AGEMA_signal_12721, new_AGEMA_signal_12717}), .c ({new_AGEMA_signal_7572, new_AGEMA_signal_7571, new_AGEMA_signal_7570, KeyReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7341, new_AGEMA_signal_7340, new_AGEMA_signal_7339, RoundKeyOutput[45]}), .a ({new_AGEMA_signal_12745, new_AGEMA_signal_12741, new_AGEMA_signal_12737, new_AGEMA_signal_12733}), .c ({new_AGEMA_signal_7578, new_AGEMA_signal_7577, new_AGEMA_signal_7576, KeyReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, new_AGEMA_signal_7342, RoundKeyOutput[46]}), .a ({new_AGEMA_signal_12761, new_AGEMA_signal_12757, new_AGEMA_signal_12753, new_AGEMA_signal_12749}), .c ({new_AGEMA_signal_7584, new_AGEMA_signal_7583, new_AGEMA_signal_7582, KeyReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7347, new_AGEMA_signal_7346, new_AGEMA_signal_7345, RoundKeyOutput[47]}), .a ({new_AGEMA_signal_12777, new_AGEMA_signal_12773, new_AGEMA_signal_12769, new_AGEMA_signal_12765}), .c ({new_AGEMA_signal_7590, new_AGEMA_signal_7589, new_AGEMA_signal_7588, KeyReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6834, new_AGEMA_signal_6833, new_AGEMA_signal_6832, RoundKeyOutput[48]}), .a ({new_AGEMA_signal_12793, new_AGEMA_signal_12789, new_AGEMA_signal_12785, new_AGEMA_signal_12781}), .c ({new_AGEMA_signal_7035, new_AGEMA_signal_7034, new_AGEMA_signal_7033, KeyReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7350, new_AGEMA_signal_7349, new_AGEMA_signal_7348, RoundKeyOutput[49]}), .a ({new_AGEMA_signal_12809, new_AGEMA_signal_12805, new_AGEMA_signal_12801, new_AGEMA_signal_12797}), .c ({new_AGEMA_signal_7596, new_AGEMA_signal_7595, new_AGEMA_signal_7594, KeyReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7353, new_AGEMA_signal_7352, new_AGEMA_signal_7351, RoundKeyOutput[50]}), .a ({new_AGEMA_signal_12825, new_AGEMA_signal_12821, new_AGEMA_signal_12817, new_AGEMA_signal_12813}), .c ({new_AGEMA_signal_7602, new_AGEMA_signal_7601, new_AGEMA_signal_7600, KeyReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7356, new_AGEMA_signal_7355, new_AGEMA_signal_7354, RoundKeyOutput[51]}), .a ({new_AGEMA_signal_12841, new_AGEMA_signal_12837, new_AGEMA_signal_12833, new_AGEMA_signal_12829}), .c ({new_AGEMA_signal_7608, new_AGEMA_signal_7607, new_AGEMA_signal_7606, KeyReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7359, new_AGEMA_signal_7358, new_AGEMA_signal_7357, RoundKeyOutput[52]}), .a ({new_AGEMA_signal_12857, new_AGEMA_signal_12853, new_AGEMA_signal_12849, new_AGEMA_signal_12845}), .c ({new_AGEMA_signal_7614, new_AGEMA_signal_7613, new_AGEMA_signal_7612, KeyReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7362, new_AGEMA_signal_7361, new_AGEMA_signal_7360, RoundKeyOutput[53]}), .a ({new_AGEMA_signal_12873, new_AGEMA_signal_12869, new_AGEMA_signal_12865, new_AGEMA_signal_12861}), .c ({new_AGEMA_signal_7620, new_AGEMA_signal_7619, new_AGEMA_signal_7618, KeyReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7365, new_AGEMA_signal_7364, new_AGEMA_signal_7363, RoundKeyOutput[54]}), .a ({new_AGEMA_signal_12889, new_AGEMA_signal_12885, new_AGEMA_signal_12881, new_AGEMA_signal_12877}), .c ({new_AGEMA_signal_7626, new_AGEMA_signal_7625, new_AGEMA_signal_7624, KeyReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, new_AGEMA_signal_7366, RoundKeyOutput[55]}), .a ({new_AGEMA_signal_12905, new_AGEMA_signal_12901, new_AGEMA_signal_12897, new_AGEMA_signal_12893}), .c ({new_AGEMA_signal_7632, new_AGEMA_signal_7631, new_AGEMA_signal_7630, KeyReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7371, new_AGEMA_signal_7370, new_AGEMA_signal_7369, RoundKeyOutput[56]}), .a ({new_AGEMA_signal_12921, new_AGEMA_signal_12917, new_AGEMA_signal_12913, new_AGEMA_signal_12909}), .c ({new_AGEMA_signal_7638, new_AGEMA_signal_7637, new_AGEMA_signal_7636, KeyReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7770, new_AGEMA_signal_7769, new_AGEMA_signal_7768, RoundKeyOutput[57]}), .a ({new_AGEMA_signal_12937, new_AGEMA_signal_12933, new_AGEMA_signal_12929, new_AGEMA_signal_12925}), .c ({new_AGEMA_signal_8082, new_AGEMA_signal_8081, new_AGEMA_signal_8080, KeyReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7773, new_AGEMA_signal_7772, new_AGEMA_signal_7771, RoundKeyOutput[58]}), .a ({new_AGEMA_signal_12953, new_AGEMA_signal_12949, new_AGEMA_signal_12945, new_AGEMA_signal_12941}), .c ({new_AGEMA_signal_8088, new_AGEMA_signal_8087, new_AGEMA_signal_8086, KeyReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7776, new_AGEMA_signal_7775, new_AGEMA_signal_7774, RoundKeyOutput[59]}), .a ({new_AGEMA_signal_12969, new_AGEMA_signal_12965, new_AGEMA_signal_12961, new_AGEMA_signal_12957}), .c ({new_AGEMA_signal_8094, new_AGEMA_signal_8093, new_AGEMA_signal_8092, KeyReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7779, new_AGEMA_signal_7778, new_AGEMA_signal_7777, RoundKeyOutput[60]}), .a ({new_AGEMA_signal_12985, new_AGEMA_signal_12981, new_AGEMA_signal_12977, new_AGEMA_signal_12973}), .c ({new_AGEMA_signal_8100, new_AGEMA_signal_8099, new_AGEMA_signal_8098, KeyReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7782, new_AGEMA_signal_7781, new_AGEMA_signal_7780, RoundKeyOutput[61]}), .a ({new_AGEMA_signal_13001, new_AGEMA_signal_12997, new_AGEMA_signal_12993, new_AGEMA_signal_12989}), .c ({new_AGEMA_signal_8106, new_AGEMA_signal_8105, new_AGEMA_signal_8104, KeyReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7785, new_AGEMA_signal_7784, new_AGEMA_signal_7783, RoundKeyOutput[62]}), .a ({new_AGEMA_signal_13017, new_AGEMA_signal_13013, new_AGEMA_signal_13009, new_AGEMA_signal_13005}), .c ({new_AGEMA_signal_8112, new_AGEMA_signal_8111, new_AGEMA_signal_8110, KeyReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7788, new_AGEMA_signal_7787, new_AGEMA_signal_7786, RoundKeyOutput[63]}), .a ({new_AGEMA_signal_13033, new_AGEMA_signal_13029, new_AGEMA_signal_13025, new_AGEMA_signal_13021}), .c ({new_AGEMA_signal_8118, new_AGEMA_signal_8117, new_AGEMA_signal_8116, KeyReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6411, new_AGEMA_signal_6410, new_AGEMA_signal_6409, RoundKeyOutput[64]}), .a ({new_AGEMA_signal_13049, new_AGEMA_signal_13045, new_AGEMA_signal_13041, new_AGEMA_signal_13037}), .c ({new_AGEMA_signal_6585, new_AGEMA_signal_6584, new_AGEMA_signal_6583, KeyReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6837, new_AGEMA_signal_6836, new_AGEMA_signal_6835, RoundKeyOutput[65]}), .a ({new_AGEMA_signal_13065, new_AGEMA_signal_13061, new_AGEMA_signal_13057, new_AGEMA_signal_13053}), .c ({new_AGEMA_signal_7041, new_AGEMA_signal_7040, new_AGEMA_signal_7039, KeyReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6840, new_AGEMA_signal_6839, new_AGEMA_signal_6838, RoundKeyOutput[66]}), .a ({new_AGEMA_signal_13081, new_AGEMA_signal_13077, new_AGEMA_signal_13073, new_AGEMA_signal_13069}), .c ({new_AGEMA_signal_7047, new_AGEMA_signal_7046, new_AGEMA_signal_7045, KeyReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6843, new_AGEMA_signal_6842, new_AGEMA_signal_6841, RoundKeyOutput[67]}), .a ({new_AGEMA_signal_13097, new_AGEMA_signal_13093, new_AGEMA_signal_13089, new_AGEMA_signal_13085}), .c ({new_AGEMA_signal_7053, new_AGEMA_signal_7052, new_AGEMA_signal_7051, KeyReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6846, new_AGEMA_signal_6845, new_AGEMA_signal_6844, RoundKeyOutput[68]}), .a ({new_AGEMA_signal_13113, new_AGEMA_signal_13109, new_AGEMA_signal_13105, new_AGEMA_signal_13101}), .c ({new_AGEMA_signal_7059, new_AGEMA_signal_7058, new_AGEMA_signal_7057, KeyReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6849, new_AGEMA_signal_6848, new_AGEMA_signal_6847, RoundKeyOutput[69]}), .a ({new_AGEMA_signal_13129, new_AGEMA_signal_13125, new_AGEMA_signal_13121, new_AGEMA_signal_13117}), .c ({new_AGEMA_signal_7065, new_AGEMA_signal_7064, new_AGEMA_signal_7063, KeyReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6852, new_AGEMA_signal_6851, new_AGEMA_signal_6850, RoundKeyOutput[70]}), .a ({new_AGEMA_signal_13145, new_AGEMA_signal_13141, new_AGEMA_signal_13137, new_AGEMA_signal_13133}), .c ({new_AGEMA_signal_7071, new_AGEMA_signal_7070, new_AGEMA_signal_7069, KeyReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6855, new_AGEMA_signal_6854, new_AGEMA_signal_6853, RoundKeyOutput[71]}), .a ({new_AGEMA_signal_13161, new_AGEMA_signal_13157, new_AGEMA_signal_13153, new_AGEMA_signal_13149}), .c ({new_AGEMA_signal_7077, new_AGEMA_signal_7076, new_AGEMA_signal_7075, KeyReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6414, new_AGEMA_signal_6413, new_AGEMA_signal_6412, RoundKeyOutput[72]}), .a ({new_AGEMA_signal_13177, new_AGEMA_signal_13173, new_AGEMA_signal_13169, new_AGEMA_signal_13165}), .c ({new_AGEMA_signal_6591, new_AGEMA_signal_6590, new_AGEMA_signal_6589, KeyReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6858, new_AGEMA_signal_6857, new_AGEMA_signal_6856, RoundKeyOutput[73]}), .a ({new_AGEMA_signal_13193, new_AGEMA_signal_13189, new_AGEMA_signal_13185, new_AGEMA_signal_13181}), .c ({new_AGEMA_signal_7083, new_AGEMA_signal_7082, new_AGEMA_signal_7081, KeyReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6861, new_AGEMA_signal_6860, new_AGEMA_signal_6859, RoundKeyOutput[74]}), .a ({new_AGEMA_signal_13209, new_AGEMA_signal_13205, new_AGEMA_signal_13201, new_AGEMA_signal_13197}), .c ({new_AGEMA_signal_7089, new_AGEMA_signal_7088, new_AGEMA_signal_7087, KeyReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6864, new_AGEMA_signal_6863, new_AGEMA_signal_6862, RoundKeyOutput[75]}), .a ({new_AGEMA_signal_13225, new_AGEMA_signal_13221, new_AGEMA_signal_13217, new_AGEMA_signal_13213}), .c ({new_AGEMA_signal_7095, new_AGEMA_signal_7094, new_AGEMA_signal_7093, KeyReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6867, new_AGEMA_signal_6866, new_AGEMA_signal_6865, RoundKeyOutput[76]}), .a ({new_AGEMA_signal_13241, new_AGEMA_signal_13237, new_AGEMA_signal_13233, new_AGEMA_signal_13229}), .c ({new_AGEMA_signal_7101, new_AGEMA_signal_7100, new_AGEMA_signal_7099, KeyReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6870, new_AGEMA_signal_6869, new_AGEMA_signal_6868, RoundKeyOutput[77]}), .a ({new_AGEMA_signal_13257, new_AGEMA_signal_13253, new_AGEMA_signal_13249, new_AGEMA_signal_13245}), .c ({new_AGEMA_signal_7107, new_AGEMA_signal_7106, new_AGEMA_signal_7105, KeyReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6873, new_AGEMA_signal_6872, new_AGEMA_signal_6871, RoundKeyOutput[78]}), .a ({new_AGEMA_signal_13273, new_AGEMA_signal_13269, new_AGEMA_signal_13265, new_AGEMA_signal_13261}), .c ({new_AGEMA_signal_7113, new_AGEMA_signal_7112, new_AGEMA_signal_7111, KeyReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6876, new_AGEMA_signal_6875, new_AGEMA_signal_6874, RoundKeyOutput[79]}), .a ({new_AGEMA_signal_13289, new_AGEMA_signal_13285, new_AGEMA_signal_13281, new_AGEMA_signal_13277}), .c ({new_AGEMA_signal_7119, new_AGEMA_signal_7118, new_AGEMA_signal_7117, KeyReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6417, new_AGEMA_signal_6416, new_AGEMA_signal_6415, RoundKeyOutput[80]}), .a ({new_AGEMA_signal_13305, new_AGEMA_signal_13301, new_AGEMA_signal_13297, new_AGEMA_signal_13293}), .c ({new_AGEMA_signal_6597, new_AGEMA_signal_6596, new_AGEMA_signal_6595, KeyReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6879, new_AGEMA_signal_6878, new_AGEMA_signal_6877, RoundKeyOutput[81]}), .a ({new_AGEMA_signal_13321, new_AGEMA_signal_13317, new_AGEMA_signal_13313, new_AGEMA_signal_13309}), .c ({new_AGEMA_signal_7125, new_AGEMA_signal_7124, new_AGEMA_signal_7123, KeyReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6882, new_AGEMA_signal_6881, new_AGEMA_signal_6880, RoundKeyOutput[82]}), .a ({new_AGEMA_signal_13337, new_AGEMA_signal_13333, new_AGEMA_signal_13329, new_AGEMA_signal_13325}), .c ({new_AGEMA_signal_7131, new_AGEMA_signal_7130, new_AGEMA_signal_7129, KeyReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6885, new_AGEMA_signal_6884, new_AGEMA_signal_6883, RoundKeyOutput[83]}), .a ({new_AGEMA_signal_13353, new_AGEMA_signal_13349, new_AGEMA_signal_13345, new_AGEMA_signal_13341}), .c ({new_AGEMA_signal_7137, new_AGEMA_signal_7136, new_AGEMA_signal_7135, KeyReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6888, new_AGEMA_signal_6887, new_AGEMA_signal_6886, RoundKeyOutput[84]}), .a ({new_AGEMA_signal_13369, new_AGEMA_signal_13365, new_AGEMA_signal_13361, new_AGEMA_signal_13357}), .c ({new_AGEMA_signal_7143, new_AGEMA_signal_7142, new_AGEMA_signal_7141, KeyReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6891, new_AGEMA_signal_6890, new_AGEMA_signal_6889, RoundKeyOutput[85]}), .a ({new_AGEMA_signal_13385, new_AGEMA_signal_13381, new_AGEMA_signal_13377, new_AGEMA_signal_13373}), .c ({new_AGEMA_signal_7149, new_AGEMA_signal_7148, new_AGEMA_signal_7147, KeyReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6894, new_AGEMA_signal_6893, new_AGEMA_signal_6892, RoundKeyOutput[86]}), .a ({new_AGEMA_signal_13401, new_AGEMA_signal_13397, new_AGEMA_signal_13393, new_AGEMA_signal_13389}), .c ({new_AGEMA_signal_7155, new_AGEMA_signal_7154, new_AGEMA_signal_7153, KeyReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6897, new_AGEMA_signal_6896, new_AGEMA_signal_6895, RoundKeyOutput[87]}), .a ({new_AGEMA_signal_13417, new_AGEMA_signal_13413, new_AGEMA_signal_13409, new_AGEMA_signal_13405}), .c ({new_AGEMA_signal_7161, new_AGEMA_signal_7160, new_AGEMA_signal_7159, KeyReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6900, new_AGEMA_signal_6899, new_AGEMA_signal_6898, RoundKeyOutput[88]}), .a ({new_AGEMA_signal_13433, new_AGEMA_signal_13429, new_AGEMA_signal_13425, new_AGEMA_signal_13421}), .c ({new_AGEMA_signal_7167, new_AGEMA_signal_7166, new_AGEMA_signal_7165, KeyReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7374, new_AGEMA_signal_7373, new_AGEMA_signal_7372, RoundKeyOutput[89]}), .a ({new_AGEMA_signal_13449, new_AGEMA_signal_13445, new_AGEMA_signal_13441, new_AGEMA_signal_13437}), .c ({new_AGEMA_signal_7644, new_AGEMA_signal_7643, new_AGEMA_signal_7642, KeyReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7377, new_AGEMA_signal_7376, new_AGEMA_signal_7375, RoundKeyOutput[90]}), .a ({new_AGEMA_signal_13465, new_AGEMA_signal_13461, new_AGEMA_signal_13457, new_AGEMA_signal_13453}), .c ({new_AGEMA_signal_7650, new_AGEMA_signal_7649, new_AGEMA_signal_7648, KeyReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7380, new_AGEMA_signal_7379, new_AGEMA_signal_7378, RoundKeyOutput[91]}), .a ({new_AGEMA_signal_13481, new_AGEMA_signal_13477, new_AGEMA_signal_13473, new_AGEMA_signal_13469}), .c ({new_AGEMA_signal_7656, new_AGEMA_signal_7655, new_AGEMA_signal_7654, KeyReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7383, new_AGEMA_signal_7382, new_AGEMA_signal_7381, RoundKeyOutput[92]}), .a ({new_AGEMA_signal_13497, new_AGEMA_signal_13493, new_AGEMA_signal_13489, new_AGEMA_signal_13485}), .c ({new_AGEMA_signal_7662, new_AGEMA_signal_7661, new_AGEMA_signal_7660, KeyReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7386, new_AGEMA_signal_7385, new_AGEMA_signal_7384, RoundKeyOutput[93]}), .a ({new_AGEMA_signal_13513, new_AGEMA_signal_13509, new_AGEMA_signal_13505, new_AGEMA_signal_13501}), .c ({new_AGEMA_signal_7668, new_AGEMA_signal_7667, new_AGEMA_signal_7666, KeyReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7389, new_AGEMA_signal_7388, new_AGEMA_signal_7387, RoundKeyOutput[94]}), .a ({new_AGEMA_signal_13529, new_AGEMA_signal_13525, new_AGEMA_signal_13521, new_AGEMA_signal_13517}), .c ({new_AGEMA_signal_7674, new_AGEMA_signal_7673, new_AGEMA_signal_7672, KeyReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_7392, new_AGEMA_signal_7391, new_AGEMA_signal_7390, RoundKeyOutput[95]}), .a ({new_AGEMA_signal_13545, new_AGEMA_signal_13541, new_AGEMA_signal_13537, new_AGEMA_signal_13533}), .c ({new_AGEMA_signal_7680, new_AGEMA_signal_7679, new_AGEMA_signal_7678, KeyReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6192, new_AGEMA_signal_6191, new_AGEMA_signal_6190, RoundKeyOutput[96]}), .a ({new_AGEMA_signal_13561, new_AGEMA_signal_13557, new_AGEMA_signal_13553, new_AGEMA_signal_13549}), .c ({new_AGEMA_signal_6300, new_AGEMA_signal_6299, new_AGEMA_signal_6298, KeyReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6420, new_AGEMA_signal_6419, new_AGEMA_signal_6418, RoundKeyOutput[97]}), .a ({new_AGEMA_signal_13577, new_AGEMA_signal_13573, new_AGEMA_signal_13569, new_AGEMA_signal_13565}), .c ({new_AGEMA_signal_6603, new_AGEMA_signal_6602, new_AGEMA_signal_6601, KeyReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6423, new_AGEMA_signal_6422, new_AGEMA_signal_6421, RoundKeyOutput[98]}), .a ({new_AGEMA_signal_13593, new_AGEMA_signal_13589, new_AGEMA_signal_13585, new_AGEMA_signal_13581}), .c ({new_AGEMA_signal_6609, new_AGEMA_signal_6608, new_AGEMA_signal_6607, KeyReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6426, new_AGEMA_signal_6425, new_AGEMA_signal_6424, RoundKeyOutput[99]}), .a ({new_AGEMA_signal_13609, new_AGEMA_signal_13605, new_AGEMA_signal_13601, new_AGEMA_signal_13597}), .c ({new_AGEMA_signal_6615, new_AGEMA_signal_6614, new_AGEMA_signal_6613, KeyReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6429, new_AGEMA_signal_6428, new_AGEMA_signal_6427, RoundKeyOutput[100]}), .a ({new_AGEMA_signal_13625, new_AGEMA_signal_13621, new_AGEMA_signal_13617, new_AGEMA_signal_13613}), .c ({new_AGEMA_signal_6621, new_AGEMA_signal_6620, new_AGEMA_signal_6619, KeyReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6432, new_AGEMA_signal_6431, new_AGEMA_signal_6430, RoundKeyOutput[101]}), .a ({new_AGEMA_signal_13641, new_AGEMA_signal_13637, new_AGEMA_signal_13633, new_AGEMA_signal_13629}), .c ({new_AGEMA_signal_6627, new_AGEMA_signal_6626, new_AGEMA_signal_6625, KeyReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6435, new_AGEMA_signal_6434, new_AGEMA_signal_6433, RoundKeyOutput[102]}), .a ({new_AGEMA_signal_13657, new_AGEMA_signal_13653, new_AGEMA_signal_13649, new_AGEMA_signal_13645}), .c ({new_AGEMA_signal_6633, new_AGEMA_signal_6632, new_AGEMA_signal_6631, KeyReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6438, new_AGEMA_signal_6437, new_AGEMA_signal_6436, RoundKeyOutput[103]}), .a ({new_AGEMA_signal_13673, new_AGEMA_signal_13669, new_AGEMA_signal_13665, new_AGEMA_signal_13661}), .c ({new_AGEMA_signal_6639, new_AGEMA_signal_6638, new_AGEMA_signal_6637, KeyReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6195, new_AGEMA_signal_6194, new_AGEMA_signal_6193, RoundKeyOutput[104]}), .a ({new_AGEMA_signal_13689, new_AGEMA_signal_13685, new_AGEMA_signal_13681, new_AGEMA_signal_13677}), .c ({new_AGEMA_signal_6306, new_AGEMA_signal_6305, new_AGEMA_signal_6304, KeyReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6441, new_AGEMA_signal_6440, new_AGEMA_signal_6439, RoundKeyOutput[105]}), .a ({new_AGEMA_signal_13705, new_AGEMA_signal_13701, new_AGEMA_signal_13697, new_AGEMA_signal_13693}), .c ({new_AGEMA_signal_6645, new_AGEMA_signal_6644, new_AGEMA_signal_6643, KeyReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6444, new_AGEMA_signal_6443, new_AGEMA_signal_6442, RoundKeyOutput[106]}), .a ({new_AGEMA_signal_13721, new_AGEMA_signal_13717, new_AGEMA_signal_13713, new_AGEMA_signal_13709}), .c ({new_AGEMA_signal_6651, new_AGEMA_signal_6650, new_AGEMA_signal_6649, KeyReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6447, new_AGEMA_signal_6446, new_AGEMA_signal_6445, RoundKeyOutput[107]}), .a ({new_AGEMA_signal_13737, new_AGEMA_signal_13733, new_AGEMA_signal_13729, new_AGEMA_signal_13725}), .c ({new_AGEMA_signal_6657, new_AGEMA_signal_6656, new_AGEMA_signal_6655, KeyReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6450, new_AGEMA_signal_6449, new_AGEMA_signal_6448, RoundKeyOutput[108]}), .a ({new_AGEMA_signal_13753, new_AGEMA_signal_13749, new_AGEMA_signal_13745, new_AGEMA_signal_13741}), .c ({new_AGEMA_signal_6663, new_AGEMA_signal_6662, new_AGEMA_signal_6661, KeyReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6453, new_AGEMA_signal_6452, new_AGEMA_signal_6451, RoundKeyOutput[109]}), .a ({new_AGEMA_signal_13769, new_AGEMA_signal_13765, new_AGEMA_signal_13761, new_AGEMA_signal_13757}), .c ({new_AGEMA_signal_6669, new_AGEMA_signal_6668, new_AGEMA_signal_6667, KeyReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6456, new_AGEMA_signal_6455, new_AGEMA_signal_6454, RoundKeyOutput[110]}), .a ({new_AGEMA_signal_13785, new_AGEMA_signal_13781, new_AGEMA_signal_13777, new_AGEMA_signal_13773}), .c ({new_AGEMA_signal_6675, new_AGEMA_signal_6674, new_AGEMA_signal_6673, KeyReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6459, new_AGEMA_signal_6458, new_AGEMA_signal_6457, RoundKeyOutput[111]}), .a ({new_AGEMA_signal_13801, new_AGEMA_signal_13797, new_AGEMA_signal_13793, new_AGEMA_signal_13789}), .c ({new_AGEMA_signal_6681, new_AGEMA_signal_6680, new_AGEMA_signal_6679, KeyReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6198, new_AGEMA_signal_6197, new_AGEMA_signal_6196, RoundKeyOutput[112]}), .a ({new_AGEMA_signal_13817, new_AGEMA_signal_13813, new_AGEMA_signal_13809, new_AGEMA_signal_13805}), .c ({new_AGEMA_signal_6312, new_AGEMA_signal_6311, new_AGEMA_signal_6310, KeyReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6462, new_AGEMA_signal_6461, new_AGEMA_signal_6460, RoundKeyOutput[113]}), .a ({new_AGEMA_signal_13833, new_AGEMA_signal_13829, new_AGEMA_signal_13825, new_AGEMA_signal_13821}), .c ({new_AGEMA_signal_6687, new_AGEMA_signal_6686, new_AGEMA_signal_6685, KeyReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6465, new_AGEMA_signal_6464, new_AGEMA_signal_6463, RoundKeyOutput[114]}), .a ({new_AGEMA_signal_13849, new_AGEMA_signal_13845, new_AGEMA_signal_13841, new_AGEMA_signal_13837}), .c ({new_AGEMA_signal_6693, new_AGEMA_signal_6692, new_AGEMA_signal_6691, KeyReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6468, new_AGEMA_signal_6467, new_AGEMA_signal_6466, RoundKeyOutput[115]}), .a ({new_AGEMA_signal_13865, new_AGEMA_signal_13861, new_AGEMA_signal_13857, new_AGEMA_signal_13853}), .c ({new_AGEMA_signal_6699, new_AGEMA_signal_6698, new_AGEMA_signal_6697, KeyReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6471, new_AGEMA_signal_6470, new_AGEMA_signal_6469, RoundKeyOutput[116]}), .a ({new_AGEMA_signal_13881, new_AGEMA_signal_13877, new_AGEMA_signal_13873, new_AGEMA_signal_13869}), .c ({new_AGEMA_signal_6705, new_AGEMA_signal_6704, new_AGEMA_signal_6703, KeyReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6474, new_AGEMA_signal_6473, new_AGEMA_signal_6472, RoundKeyOutput[117]}), .a ({new_AGEMA_signal_13897, new_AGEMA_signal_13893, new_AGEMA_signal_13889, new_AGEMA_signal_13885}), .c ({new_AGEMA_signal_6711, new_AGEMA_signal_6710, new_AGEMA_signal_6709, KeyReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6477, new_AGEMA_signal_6476, new_AGEMA_signal_6475, RoundKeyOutput[118]}), .a ({new_AGEMA_signal_13913, new_AGEMA_signal_13909, new_AGEMA_signal_13905, new_AGEMA_signal_13901}), .c ({new_AGEMA_signal_6717, new_AGEMA_signal_6716, new_AGEMA_signal_6715, KeyReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6480, new_AGEMA_signal_6479, new_AGEMA_signal_6478, RoundKeyOutput[119]}), .a ({new_AGEMA_signal_13929, new_AGEMA_signal_13925, new_AGEMA_signal_13921, new_AGEMA_signal_13917}), .c ({new_AGEMA_signal_6723, new_AGEMA_signal_6722, new_AGEMA_signal_6721, KeyReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6483, new_AGEMA_signal_6482, new_AGEMA_signal_6481, RoundKeyOutput[120]}), .a ({new_AGEMA_signal_13945, new_AGEMA_signal_13941, new_AGEMA_signal_13937, new_AGEMA_signal_13933}), .c ({new_AGEMA_signal_6729, new_AGEMA_signal_6728, new_AGEMA_signal_6727, KeyReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6903, new_AGEMA_signal_6902, new_AGEMA_signal_6901, RoundKeyOutput[121]}), .a ({new_AGEMA_signal_13961, new_AGEMA_signal_13957, new_AGEMA_signal_13953, new_AGEMA_signal_13949}), .c ({new_AGEMA_signal_7173, new_AGEMA_signal_7172, new_AGEMA_signal_7171, KeyReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6906, new_AGEMA_signal_6905, new_AGEMA_signal_6904, RoundKeyOutput[122]}), .a ({new_AGEMA_signal_13977, new_AGEMA_signal_13973, new_AGEMA_signal_13969, new_AGEMA_signal_13965}), .c ({new_AGEMA_signal_7179, new_AGEMA_signal_7178, new_AGEMA_signal_7177, KeyReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6909, new_AGEMA_signal_6908, new_AGEMA_signal_6907, RoundKeyOutput[123]}), .a ({new_AGEMA_signal_13993, new_AGEMA_signal_13989, new_AGEMA_signal_13985, new_AGEMA_signal_13981}), .c ({new_AGEMA_signal_7185, new_AGEMA_signal_7184, new_AGEMA_signal_7183, KeyReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6912, new_AGEMA_signal_6911, new_AGEMA_signal_6910, RoundKeyOutput[124]}), .a ({new_AGEMA_signal_14009, new_AGEMA_signal_14005, new_AGEMA_signal_14001, new_AGEMA_signal_13997}), .c ({new_AGEMA_signal_7191, new_AGEMA_signal_7190, new_AGEMA_signal_7189, KeyReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6915, new_AGEMA_signal_6914, new_AGEMA_signal_6913, RoundKeyOutput[125]}), .a ({new_AGEMA_signal_14025, new_AGEMA_signal_14021, new_AGEMA_signal_14017, new_AGEMA_signal_14013}), .c ({new_AGEMA_signal_7197, new_AGEMA_signal_7196, new_AGEMA_signal_7195, KeyReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6918, new_AGEMA_signal_6917, new_AGEMA_signal_6916, RoundKeyOutput[126]}), .a ({new_AGEMA_signal_14041, new_AGEMA_signal_14037, new_AGEMA_signal_14033, new_AGEMA_signal_14029}), .c ({new_AGEMA_signal_7203, new_AGEMA_signal_7202, new_AGEMA_signal_7201, KeyReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (new_AGEMA_signal_10081), .b ({new_AGEMA_signal_6921, new_AGEMA_signal_6920, new_AGEMA_signal_6919, RoundKeyOutput[127]}), .a ({new_AGEMA_signal_14057, new_AGEMA_signal_14053, new_AGEMA_signal_14049, new_AGEMA_signal_14045}), .c ({new_AGEMA_signal_7209, new_AGEMA_signal_7208, new_AGEMA_signal_7207, KeyReg_Inst_ff_SDE_127_next_state}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U128 ( .a ({new_AGEMA_signal_14073, new_AGEMA_signal_14069, new_AGEMA_signal_14065, new_AGEMA_signal_14061}), .b ({new_AGEMA_signal_6735, new_AGEMA_signal_6734, new_AGEMA_signal_6733, KeyExpansionOutput[41]}), .c ({new_AGEMA_signal_7212, new_AGEMA_signal_7211, new_AGEMA_signal_7210, KeyExpansionOutput[9]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U127 ( .a ({new_AGEMA_signal_14089, new_AGEMA_signal_14085, new_AGEMA_signal_14081, new_AGEMA_signal_14077}), .b ({new_AGEMA_signal_6318, new_AGEMA_signal_6317, new_AGEMA_signal_6316, KeyExpansionOutput[40]}), .c ({new_AGEMA_signal_6732, new_AGEMA_signal_6731, new_AGEMA_signal_6730, KeyExpansionOutput[8]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U126 ( .a ({new_AGEMA_signal_14105, new_AGEMA_signal_14101, new_AGEMA_signal_14097, new_AGEMA_signal_14093}), .b ({new_AGEMA_signal_6738, new_AGEMA_signal_6737, new_AGEMA_signal_6736, KeyExpansionOutput[39]}), .c ({new_AGEMA_signal_7215, new_AGEMA_signal_7214, new_AGEMA_signal_7213, KeyExpansionOutput[7]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U125 ( .a ({new_AGEMA_signal_14121, new_AGEMA_signal_14117, new_AGEMA_signal_14113, new_AGEMA_signal_14109}), .b ({new_AGEMA_signal_6741, new_AGEMA_signal_6740, new_AGEMA_signal_6739, KeyExpansionOutput[38]}), .c ({new_AGEMA_signal_7218, new_AGEMA_signal_7217, new_AGEMA_signal_7216, KeyExpansionOutput[6]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U124 ( .a ({new_AGEMA_signal_14137, new_AGEMA_signal_14133, new_AGEMA_signal_14129, new_AGEMA_signal_14125}), .b ({new_AGEMA_signal_6744, new_AGEMA_signal_6743, new_AGEMA_signal_6742, KeyExpansionOutput[37]}), .c ({new_AGEMA_signal_7221, new_AGEMA_signal_7220, new_AGEMA_signal_7219, KeyExpansionOutput[5]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U123 ( .a ({new_AGEMA_signal_14153, new_AGEMA_signal_14149, new_AGEMA_signal_14145, new_AGEMA_signal_14141}), .b ({new_AGEMA_signal_6747, new_AGEMA_signal_6746, new_AGEMA_signal_6745, KeyExpansionOutput[36]}), .c ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, new_AGEMA_signal_7222, KeyExpansionOutput[4]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U122 ( .a ({new_AGEMA_signal_14169, new_AGEMA_signal_14165, new_AGEMA_signal_14161, new_AGEMA_signal_14157}), .b ({new_AGEMA_signal_6315, new_AGEMA_signal_6314, new_AGEMA_signal_6313, KeyExpansionOutput[73]}), .c ({new_AGEMA_signal_6735, new_AGEMA_signal_6734, new_AGEMA_signal_6733, KeyExpansionOutput[41]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U121 ( .a ({new_AGEMA_signal_14185, new_AGEMA_signal_14181, new_AGEMA_signal_14177, new_AGEMA_signal_14173}), .b ({new_AGEMA_signal_6153, new_AGEMA_signal_6152, new_AGEMA_signal_6151, KeyExpansionOutput[105]}), .c ({new_AGEMA_signal_6315, new_AGEMA_signal_6314, new_AGEMA_signal_6313, KeyExpansionOutput[73]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U120 ( .a ({new_AGEMA_signal_14201, new_AGEMA_signal_14197, new_AGEMA_signal_14193, new_AGEMA_signal_14189}), .b ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, new_AGEMA_signal_6094, KeyExpansionOutput[72]}), .c ({new_AGEMA_signal_6318, new_AGEMA_signal_6317, new_AGEMA_signal_6316, KeyExpansionOutput[40]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U119 ( .a ({new_AGEMA_signal_14217, new_AGEMA_signal_14213, new_AGEMA_signal_14209, new_AGEMA_signal_14205}), .b ({new_AGEMA_signal_5991, new_AGEMA_signal_5990, new_AGEMA_signal_5989, KeyExpansionOutput[104]}), .c ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, new_AGEMA_signal_6094, KeyExpansionOutput[72]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U118 ( .a ({new_AGEMA_signal_14233, new_AGEMA_signal_14229, new_AGEMA_signal_14225, new_AGEMA_signal_14221}), .b ({new_AGEMA_signal_6750, new_AGEMA_signal_6749, new_AGEMA_signal_6748, KeyExpansionOutput[35]}), .c ({new_AGEMA_signal_7227, new_AGEMA_signal_7226, new_AGEMA_signal_7225, KeyExpansionOutput[3]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U117 ( .a ({new_AGEMA_signal_14249, new_AGEMA_signal_14245, new_AGEMA_signal_14241, new_AGEMA_signal_14237}), .b ({new_AGEMA_signal_6321, new_AGEMA_signal_6320, new_AGEMA_signal_6319, KeyExpansionOutput[71]}), .c ({new_AGEMA_signal_6738, new_AGEMA_signal_6737, new_AGEMA_signal_6736, KeyExpansionOutput[39]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U116 ( .a ({new_AGEMA_signal_14265, new_AGEMA_signal_14261, new_AGEMA_signal_14257, new_AGEMA_signal_14253}), .b ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, new_AGEMA_signal_6154, KeyExpansionOutput[103]}), .c ({new_AGEMA_signal_6321, new_AGEMA_signal_6320, new_AGEMA_signal_6319, KeyExpansionOutput[71]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U115 ( .a ({new_AGEMA_signal_14281, new_AGEMA_signal_14277, new_AGEMA_signal_14273, new_AGEMA_signal_14269}), .b ({new_AGEMA_signal_6324, new_AGEMA_signal_6323, new_AGEMA_signal_6322, KeyExpansionOutput[70]}), .c ({new_AGEMA_signal_6741, new_AGEMA_signal_6740, new_AGEMA_signal_6739, KeyExpansionOutput[38]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U114 ( .a ({new_AGEMA_signal_14297, new_AGEMA_signal_14293, new_AGEMA_signal_14289, new_AGEMA_signal_14285}), .b ({new_AGEMA_signal_6159, new_AGEMA_signal_6158, new_AGEMA_signal_6157, KeyExpansionOutput[102]}), .c ({new_AGEMA_signal_6324, new_AGEMA_signal_6323, new_AGEMA_signal_6322, KeyExpansionOutput[70]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U113 ( .a ({new_AGEMA_signal_14313, new_AGEMA_signal_14309, new_AGEMA_signal_14305, new_AGEMA_signal_14301}), .b ({new_AGEMA_signal_6327, new_AGEMA_signal_6326, new_AGEMA_signal_6325, KeyExpansionOutput[69]}), .c ({new_AGEMA_signal_6744, new_AGEMA_signal_6743, new_AGEMA_signal_6742, KeyExpansionOutput[37]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U112 ( .a ({new_AGEMA_signal_14329, new_AGEMA_signal_14325, new_AGEMA_signal_14321, new_AGEMA_signal_14317}), .b ({new_AGEMA_signal_6162, new_AGEMA_signal_6161, new_AGEMA_signal_6160, KeyExpansionOutput[101]}), .c ({new_AGEMA_signal_6327, new_AGEMA_signal_6326, new_AGEMA_signal_6325, KeyExpansionOutput[69]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U111 ( .a ({new_AGEMA_signal_14345, new_AGEMA_signal_14341, new_AGEMA_signal_14337, new_AGEMA_signal_14333}), .b ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, new_AGEMA_signal_6328, KeyExpansionOutput[68]}), .c ({new_AGEMA_signal_6747, new_AGEMA_signal_6746, new_AGEMA_signal_6745, KeyExpansionOutput[36]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U110 ( .a ({new_AGEMA_signal_14361, new_AGEMA_signal_14357, new_AGEMA_signal_14353, new_AGEMA_signal_14349}), .b ({new_AGEMA_signal_6165, new_AGEMA_signal_6164, new_AGEMA_signal_6163, KeyExpansionOutput[100]}), .c ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, new_AGEMA_signal_6328, KeyExpansionOutput[68]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U109 ( .a ({new_AGEMA_signal_14377, new_AGEMA_signal_14373, new_AGEMA_signal_14369, new_AGEMA_signal_14365}), .b ({new_AGEMA_signal_6333, new_AGEMA_signal_6332, new_AGEMA_signal_6331, KeyExpansionOutput[67]}), .c ({new_AGEMA_signal_6750, new_AGEMA_signal_6749, new_AGEMA_signal_6748, KeyExpansionOutput[35]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U108 ( .a ({new_AGEMA_signal_14393, new_AGEMA_signal_14389, new_AGEMA_signal_14385, new_AGEMA_signal_14381}), .b ({new_AGEMA_signal_6099, new_AGEMA_signal_6098, new_AGEMA_signal_6097, KeyExpansionOutput[99]}), .c ({new_AGEMA_signal_6333, new_AGEMA_signal_6332, new_AGEMA_signal_6331, KeyExpansionOutput[67]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U107 ( .a ({new_AGEMA_signal_14409, new_AGEMA_signal_14405, new_AGEMA_signal_14401, new_AGEMA_signal_14397}), .b ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, new_AGEMA_signal_5977, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_6099, new_AGEMA_signal_6098, new_AGEMA_signal_6097, KeyExpansionOutput[99]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U106 ( .a ({new_AGEMA_signal_14425, new_AGEMA_signal_14421, new_AGEMA_signal_14417, new_AGEMA_signal_14413}), .b ({new_AGEMA_signal_7230, new_AGEMA_signal_7229, new_AGEMA_signal_7228, KeyExpansionOutput[63]}), .c ({new_AGEMA_signal_7683, new_AGEMA_signal_7682, new_AGEMA_signal_7681, KeyExpansionOutput[31]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U105 ( .a ({new_AGEMA_signal_14441, new_AGEMA_signal_14437, new_AGEMA_signal_14433, new_AGEMA_signal_14429}), .b ({new_AGEMA_signal_6753, new_AGEMA_signal_6752, new_AGEMA_signal_6751, KeyExpansionOutput[95]}), .c ({new_AGEMA_signal_7230, new_AGEMA_signal_7229, new_AGEMA_signal_7228, KeyExpansionOutput[63]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U104 ( .a ({new_AGEMA_signal_14457, new_AGEMA_signal_14453, new_AGEMA_signal_14449, new_AGEMA_signal_14445}), .b ({new_AGEMA_signal_6381, new_AGEMA_signal_6380, new_AGEMA_signal_6379, KeyExpansionOutput[127]}), .c ({new_AGEMA_signal_6753, new_AGEMA_signal_6752, new_AGEMA_signal_6751, KeyExpansionOutput[95]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U103 ( .a ({new_AGEMA_signal_14473, new_AGEMA_signal_14469, new_AGEMA_signal_14465, new_AGEMA_signal_14461}), .b ({new_AGEMA_signal_7233, new_AGEMA_signal_7232, new_AGEMA_signal_7231, KeyExpansionOutput[62]}), .c ({new_AGEMA_signal_7686, new_AGEMA_signal_7685, new_AGEMA_signal_7684, KeyExpansionOutput[30]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U102 ( .a ({new_AGEMA_signal_14489, new_AGEMA_signal_14485, new_AGEMA_signal_14481, new_AGEMA_signal_14477}), .b ({new_AGEMA_signal_6756, new_AGEMA_signal_6755, new_AGEMA_signal_6754, KeyExpansionOutput[94]}), .c ({new_AGEMA_signal_7233, new_AGEMA_signal_7232, new_AGEMA_signal_7231, KeyExpansionOutput[62]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U101 ( .a ({new_AGEMA_signal_14505, new_AGEMA_signal_14501, new_AGEMA_signal_14497, new_AGEMA_signal_14493}), .b ({new_AGEMA_signal_6384, new_AGEMA_signal_6383, new_AGEMA_signal_6382, KeyExpansionOutput[126]}), .c ({new_AGEMA_signal_6756, new_AGEMA_signal_6755, new_AGEMA_signal_6754, KeyExpansionOutput[94]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U100 ( .a ({new_AGEMA_signal_14521, new_AGEMA_signal_14517, new_AGEMA_signal_14513, new_AGEMA_signal_14509}), .b ({new_AGEMA_signal_6759, new_AGEMA_signal_6758, new_AGEMA_signal_6757, KeyExpansionOutput[34]}), .c ({new_AGEMA_signal_7236, new_AGEMA_signal_7235, new_AGEMA_signal_7234, KeyExpansionOutput[2]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U99 ( .a ({new_AGEMA_signal_14537, new_AGEMA_signal_14533, new_AGEMA_signal_14529, new_AGEMA_signal_14525}), .b ({new_AGEMA_signal_6336, new_AGEMA_signal_6335, new_AGEMA_signal_6334, KeyExpansionOutput[66]}), .c ({new_AGEMA_signal_6759, new_AGEMA_signal_6758, new_AGEMA_signal_6757, KeyExpansionOutput[34]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U98 ( .a ({new_AGEMA_signal_14553, new_AGEMA_signal_14549, new_AGEMA_signal_14545, new_AGEMA_signal_14541}), .b ({new_AGEMA_signal_6102, new_AGEMA_signal_6101, new_AGEMA_signal_6100, KeyExpansionOutput[98]}), .c ({new_AGEMA_signal_6336, new_AGEMA_signal_6335, new_AGEMA_signal_6334, KeyExpansionOutput[66]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U97 ( .a ({new_AGEMA_signal_14569, new_AGEMA_signal_14565, new_AGEMA_signal_14561, new_AGEMA_signal_14557}), .b ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, new_AGEMA_signal_5980, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_6102, new_AGEMA_signal_6101, new_AGEMA_signal_6100, KeyExpansionOutput[98]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U96 ( .a ({new_AGEMA_signal_14585, new_AGEMA_signal_14581, new_AGEMA_signal_14577, new_AGEMA_signal_14573}), .b ({new_AGEMA_signal_7239, new_AGEMA_signal_7238, new_AGEMA_signal_7237, KeyExpansionOutput[61]}), .c ({new_AGEMA_signal_7689, new_AGEMA_signal_7688, new_AGEMA_signal_7687, KeyExpansionOutput[29]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U95 ( .a ({new_AGEMA_signal_14601, new_AGEMA_signal_14597, new_AGEMA_signal_14593, new_AGEMA_signal_14589}), .b ({new_AGEMA_signal_6762, new_AGEMA_signal_6761, new_AGEMA_signal_6760, KeyExpansionOutput[93]}), .c ({new_AGEMA_signal_7239, new_AGEMA_signal_7238, new_AGEMA_signal_7237, KeyExpansionOutput[61]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U94 ( .a ({new_AGEMA_signal_14617, new_AGEMA_signal_14613, new_AGEMA_signal_14609, new_AGEMA_signal_14605}), .b ({new_AGEMA_signal_6387, new_AGEMA_signal_6386, new_AGEMA_signal_6385, KeyExpansionOutput[125]}), .c ({new_AGEMA_signal_6762, new_AGEMA_signal_6761, new_AGEMA_signal_6760, KeyExpansionOutput[93]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U93 ( .a ({new_AGEMA_signal_14633, new_AGEMA_signal_14629, new_AGEMA_signal_14625, new_AGEMA_signal_14621}), .b ({new_AGEMA_signal_7242, new_AGEMA_signal_7241, new_AGEMA_signal_7240, KeyExpansionOutput[60]}), .c ({new_AGEMA_signal_7692, new_AGEMA_signal_7691, new_AGEMA_signal_7690, KeyExpansionOutput[28]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U92 ( .a ({new_AGEMA_signal_14649, new_AGEMA_signal_14645, new_AGEMA_signal_14641, new_AGEMA_signal_14637}), .b ({new_AGEMA_signal_6765, new_AGEMA_signal_6764, new_AGEMA_signal_6763, KeyExpansionOutput[92]}), .c ({new_AGEMA_signal_7242, new_AGEMA_signal_7241, new_AGEMA_signal_7240, KeyExpansionOutput[60]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U91 ( .a ({new_AGEMA_signal_14665, new_AGEMA_signal_14661, new_AGEMA_signal_14657, new_AGEMA_signal_14653}), .b ({new_AGEMA_signal_6390, new_AGEMA_signal_6389, new_AGEMA_signal_6388, KeyExpansionOutput[124]}), .c ({new_AGEMA_signal_6765, new_AGEMA_signal_6764, new_AGEMA_signal_6763, KeyExpansionOutput[92]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U90 ( .a ({new_AGEMA_signal_14681, new_AGEMA_signal_14677, new_AGEMA_signal_14673, new_AGEMA_signal_14669}), .b ({new_AGEMA_signal_7245, new_AGEMA_signal_7244, new_AGEMA_signal_7243, KeyExpansionOutput[59]}), .c ({new_AGEMA_signal_7695, new_AGEMA_signal_7694, new_AGEMA_signal_7693, KeyExpansionOutput[27]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U89 ( .a ({new_AGEMA_signal_14697, new_AGEMA_signal_14693, new_AGEMA_signal_14689, new_AGEMA_signal_14685}), .b ({new_AGEMA_signal_6768, new_AGEMA_signal_6767, new_AGEMA_signal_6766, KeyExpansionOutput[91]}), .c ({new_AGEMA_signal_7245, new_AGEMA_signal_7244, new_AGEMA_signal_7243, KeyExpansionOutput[59]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U88 ( .a ({new_AGEMA_signal_14713, new_AGEMA_signal_14709, new_AGEMA_signal_14705, new_AGEMA_signal_14701}), .b ({new_AGEMA_signal_6393, new_AGEMA_signal_6392, new_AGEMA_signal_6391, KeyExpansionOutput[123]}), .c ({new_AGEMA_signal_6768, new_AGEMA_signal_6767, new_AGEMA_signal_6766, KeyExpansionOutput[91]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U87 ( .a ({new_AGEMA_signal_14729, new_AGEMA_signal_14725, new_AGEMA_signal_14721, new_AGEMA_signal_14717}), .b ({new_AGEMA_signal_7248, new_AGEMA_signal_7247, new_AGEMA_signal_7246, KeyExpansionOutput[58]}), .c ({new_AGEMA_signal_7698, new_AGEMA_signal_7697, new_AGEMA_signal_7696, KeyExpansionOutput[26]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U86 ( .a ({new_AGEMA_signal_14745, new_AGEMA_signal_14741, new_AGEMA_signal_14737, new_AGEMA_signal_14733}), .b ({new_AGEMA_signal_6771, new_AGEMA_signal_6770, new_AGEMA_signal_6769, KeyExpansionOutput[90]}), .c ({new_AGEMA_signal_7248, new_AGEMA_signal_7247, new_AGEMA_signal_7246, KeyExpansionOutput[58]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U85 ( .a ({new_AGEMA_signal_14761, new_AGEMA_signal_14757, new_AGEMA_signal_14753, new_AGEMA_signal_14749}), .b ({new_AGEMA_signal_6396, new_AGEMA_signal_6395, new_AGEMA_signal_6394, KeyExpansionOutput[122]}), .c ({new_AGEMA_signal_6771, new_AGEMA_signal_6770, new_AGEMA_signal_6769, KeyExpansionOutput[90]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U84 ( .a ({new_AGEMA_signal_14777, new_AGEMA_signal_14773, new_AGEMA_signal_14769, new_AGEMA_signal_14765}), .b ({new_AGEMA_signal_7251, new_AGEMA_signal_7250, new_AGEMA_signal_7249, KeyExpansionOutput[57]}), .c ({new_AGEMA_signal_7701, new_AGEMA_signal_7700, new_AGEMA_signal_7699, KeyExpansionOutput[25]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U83 ( .a ({new_AGEMA_signal_14793, new_AGEMA_signal_14789, new_AGEMA_signal_14785, new_AGEMA_signal_14781}), .b ({new_AGEMA_signal_6774, new_AGEMA_signal_6773, new_AGEMA_signal_6772, KeyExpansionOutput[89]}), .c ({new_AGEMA_signal_7251, new_AGEMA_signal_7250, new_AGEMA_signal_7249, KeyExpansionOutput[57]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U82 ( .a ({new_AGEMA_signal_14809, new_AGEMA_signal_14805, new_AGEMA_signal_14801, new_AGEMA_signal_14797}), .b ({new_AGEMA_signal_6399, new_AGEMA_signal_6398, new_AGEMA_signal_6397, KeyExpansionOutput[121]}), .c ({new_AGEMA_signal_6774, new_AGEMA_signal_6773, new_AGEMA_signal_6772, KeyExpansionOutput[89]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U81 ( .a ({new_AGEMA_signal_14825, new_AGEMA_signal_14821, new_AGEMA_signal_14817, new_AGEMA_signal_14813}), .b ({new_AGEMA_signal_6777, new_AGEMA_signal_6776, new_AGEMA_signal_6775, KeyExpansionOutput[56]}), .c ({new_AGEMA_signal_7254, new_AGEMA_signal_7253, new_AGEMA_signal_7252, KeyExpansionOutput[24]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U80 ( .a ({new_AGEMA_signal_14841, new_AGEMA_signal_14837, new_AGEMA_signal_14833, new_AGEMA_signal_14829}), .b ({new_AGEMA_signal_6339, new_AGEMA_signal_6338, new_AGEMA_signal_6337, KeyExpansionOutput[88]}), .c ({new_AGEMA_signal_6777, new_AGEMA_signal_6776, new_AGEMA_signal_6775, KeyExpansionOutput[56]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U79 ( .a ({new_AGEMA_signal_14857, new_AGEMA_signal_14853, new_AGEMA_signal_14849, new_AGEMA_signal_14845}), .b ({new_AGEMA_signal_6111, new_AGEMA_signal_6110, new_AGEMA_signal_6109, KeyExpansionOutput[120]}), .c ({new_AGEMA_signal_6339, new_AGEMA_signal_6338, new_AGEMA_signal_6337, KeyExpansionOutput[88]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U78 ( .a ({new_AGEMA_signal_14873, new_AGEMA_signal_14869, new_AGEMA_signal_14865, new_AGEMA_signal_14861}), .b ({new_AGEMA_signal_6780, new_AGEMA_signal_6779, new_AGEMA_signal_6778, KeyExpansionOutput[55]}), .c ({new_AGEMA_signal_7257, new_AGEMA_signal_7256, new_AGEMA_signal_7255, KeyExpansionOutput[23]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U77 ( .a ({new_AGEMA_signal_14889, new_AGEMA_signal_14885, new_AGEMA_signal_14881, new_AGEMA_signal_14877}), .b ({new_AGEMA_signal_6342, new_AGEMA_signal_6341, new_AGEMA_signal_6340, KeyExpansionOutput[87]}), .c ({new_AGEMA_signal_6780, new_AGEMA_signal_6779, new_AGEMA_signal_6778, KeyExpansionOutput[55]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U76 ( .a ({new_AGEMA_signal_14905, new_AGEMA_signal_14901, new_AGEMA_signal_14897, new_AGEMA_signal_14893}), .b ({new_AGEMA_signal_6114, new_AGEMA_signal_6113, new_AGEMA_signal_6112, KeyExpansionOutput[119]}), .c ({new_AGEMA_signal_6342, new_AGEMA_signal_6341, new_AGEMA_signal_6340, KeyExpansionOutput[87]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U75 ( .a ({new_AGEMA_signal_14921, new_AGEMA_signal_14917, new_AGEMA_signal_14913, new_AGEMA_signal_14909}), .b ({new_AGEMA_signal_6783, new_AGEMA_signal_6782, new_AGEMA_signal_6781, KeyExpansionOutput[54]}), .c ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, new_AGEMA_signal_7258, KeyExpansionOutput[22]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U74 ( .a ({new_AGEMA_signal_14937, new_AGEMA_signal_14933, new_AGEMA_signal_14929, new_AGEMA_signal_14925}), .b ({new_AGEMA_signal_6345, new_AGEMA_signal_6344, new_AGEMA_signal_6343, KeyExpansionOutput[86]}), .c ({new_AGEMA_signal_6783, new_AGEMA_signal_6782, new_AGEMA_signal_6781, KeyExpansionOutput[54]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U73 ( .a ({new_AGEMA_signal_14953, new_AGEMA_signal_14949, new_AGEMA_signal_14945, new_AGEMA_signal_14941}), .b ({new_AGEMA_signal_6117, new_AGEMA_signal_6116, new_AGEMA_signal_6115, KeyExpansionOutput[118]}), .c ({new_AGEMA_signal_6345, new_AGEMA_signal_6344, new_AGEMA_signal_6343, KeyExpansionOutput[86]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U72 ( .a ({new_AGEMA_signal_14969, new_AGEMA_signal_14965, new_AGEMA_signal_14961, new_AGEMA_signal_14957}), .b ({new_AGEMA_signal_6786, new_AGEMA_signal_6785, new_AGEMA_signal_6784, KeyExpansionOutput[53]}), .c ({new_AGEMA_signal_7263, new_AGEMA_signal_7262, new_AGEMA_signal_7261, KeyExpansionOutput[21]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U71 ( .a ({new_AGEMA_signal_14985, new_AGEMA_signal_14981, new_AGEMA_signal_14977, new_AGEMA_signal_14973}), .b ({new_AGEMA_signal_6348, new_AGEMA_signal_6347, new_AGEMA_signal_6346, KeyExpansionOutput[85]}), .c ({new_AGEMA_signal_6786, new_AGEMA_signal_6785, new_AGEMA_signal_6784, KeyExpansionOutput[53]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U70 ( .a ({new_AGEMA_signal_15001, new_AGEMA_signal_14997, new_AGEMA_signal_14993, new_AGEMA_signal_14989}), .b ({new_AGEMA_signal_6120, new_AGEMA_signal_6119, new_AGEMA_signal_6118, KeyExpansionOutput[117]}), .c ({new_AGEMA_signal_6348, new_AGEMA_signal_6347, new_AGEMA_signal_6346, KeyExpansionOutput[85]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U69 ( .a ({new_AGEMA_signal_15017, new_AGEMA_signal_15013, new_AGEMA_signal_15009, new_AGEMA_signal_15005}), .b ({new_AGEMA_signal_6789, new_AGEMA_signal_6788, new_AGEMA_signal_6787, KeyExpansionOutput[52]}), .c ({new_AGEMA_signal_7266, new_AGEMA_signal_7265, new_AGEMA_signal_7264, KeyExpansionOutput[20]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U68 ( .a ({new_AGEMA_signal_15033, new_AGEMA_signal_15029, new_AGEMA_signal_15025, new_AGEMA_signal_15021}), .b ({new_AGEMA_signal_6351, new_AGEMA_signal_6350, new_AGEMA_signal_6349, KeyExpansionOutput[84]}), .c ({new_AGEMA_signal_6789, new_AGEMA_signal_6788, new_AGEMA_signal_6787, KeyExpansionOutput[52]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U67 ( .a ({new_AGEMA_signal_15049, new_AGEMA_signal_15045, new_AGEMA_signal_15041, new_AGEMA_signal_15037}), .b ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, new_AGEMA_signal_6121, KeyExpansionOutput[116]}), .c ({new_AGEMA_signal_6351, new_AGEMA_signal_6350, new_AGEMA_signal_6349, KeyExpansionOutput[84]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U66 ( .a ({new_AGEMA_signal_15065, new_AGEMA_signal_15061, new_AGEMA_signal_15057, new_AGEMA_signal_15053}), .b ({new_AGEMA_signal_6792, new_AGEMA_signal_6791, new_AGEMA_signal_6790, KeyExpansionOutput[33]}), .c ({new_AGEMA_signal_7269, new_AGEMA_signal_7268, new_AGEMA_signal_7267, KeyExpansionOutput[1]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U65 ( .a ({new_AGEMA_signal_15081, new_AGEMA_signal_15077, new_AGEMA_signal_15073, new_AGEMA_signal_15069}), .b ({new_AGEMA_signal_6354, new_AGEMA_signal_6353, new_AGEMA_signal_6352, KeyExpansionOutput[65]}), .c ({new_AGEMA_signal_6792, new_AGEMA_signal_6791, new_AGEMA_signal_6790, KeyExpansionOutput[33]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U64 ( .a ({new_AGEMA_signal_15097, new_AGEMA_signal_15093, new_AGEMA_signal_15089, new_AGEMA_signal_15085}), .b ({new_AGEMA_signal_6105, new_AGEMA_signal_6104, new_AGEMA_signal_6103, KeyExpansionOutput[97]}), .c ({new_AGEMA_signal_6354, new_AGEMA_signal_6353, new_AGEMA_signal_6352, KeyExpansionOutput[65]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U63 ( .a ({new_AGEMA_signal_15113, new_AGEMA_signal_15109, new_AGEMA_signal_15105, new_AGEMA_signal_15101}), .b ({new_AGEMA_signal_5985, new_AGEMA_signal_5984, new_AGEMA_signal_5983, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_6105, new_AGEMA_signal_6104, new_AGEMA_signal_6103, KeyExpansionOutput[97]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U62 ( .a ({new_AGEMA_signal_15129, new_AGEMA_signal_15125, new_AGEMA_signal_15121, new_AGEMA_signal_15117}), .b ({new_AGEMA_signal_6795, new_AGEMA_signal_6794, new_AGEMA_signal_6793, KeyExpansionOutput[51]}), .c ({new_AGEMA_signal_7272, new_AGEMA_signal_7271, new_AGEMA_signal_7270, KeyExpansionOutput[19]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U61 ( .a ({new_AGEMA_signal_15145, new_AGEMA_signal_15141, new_AGEMA_signal_15137, new_AGEMA_signal_15133}), .b ({new_AGEMA_signal_6357, new_AGEMA_signal_6356, new_AGEMA_signal_6355, KeyExpansionOutput[83]}), .c ({new_AGEMA_signal_6795, new_AGEMA_signal_6794, new_AGEMA_signal_6793, KeyExpansionOutput[51]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U60 ( .a ({new_AGEMA_signal_15161, new_AGEMA_signal_15157, new_AGEMA_signal_15153, new_AGEMA_signal_15149}), .b ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, new_AGEMA_signal_6124, KeyExpansionOutput[115]}), .c ({new_AGEMA_signal_6357, new_AGEMA_signal_6356, new_AGEMA_signal_6355, KeyExpansionOutput[83]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U59 ( .a ({new_AGEMA_signal_15177, new_AGEMA_signal_15173, new_AGEMA_signal_15169, new_AGEMA_signal_15165}), .b ({new_AGEMA_signal_6798, new_AGEMA_signal_6797, new_AGEMA_signal_6796, KeyExpansionOutput[50]}), .c ({new_AGEMA_signal_7275, new_AGEMA_signal_7274, new_AGEMA_signal_7273, KeyExpansionOutput[18]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U58 ( .a ({new_AGEMA_signal_15193, new_AGEMA_signal_15189, new_AGEMA_signal_15185, new_AGEMA_signal_15181}), .b ({new_AGEMA_signal_6360, new_AGEMA_signal_6359, new_AGEMA_signal_6358, KeyExpansionOutput[82]}), .c ({new_AGEMA_signal_6798, new_AGEMA_signal_6797, new_AGEMA_signal_6796, KeyExpansionOutput[50]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U57 ( .a ({new_AGEMA_signal_15209, new_AGEMA_signal_15205, new_AGEMA_signal_15201, new_AGEMA_signal_15197}), .b ({new_AGEMA_signal_6129, new_AGEMA_signal_6128, new_AGEMA_signal_6127, KeyExpansionOutput[114]}), .c ({new_AGEMA_signal_6360, new_AGEMA_signal_6359, new_AGEMA_signal_6358, KeyExpansionOutput[82]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U56 ( .a ({new_AGEMA_signal_15225, new_AGEMA_signal_15221, new_AGEMA_signal_15217, new_AGEMA_signal_15213}), .b ({new_AGEMA_signal_6801, new_AGEMA_signal_6800, new_AGEMA_signal_6799, KeyExpansionOutput[49]}), .c ({new_AGEMA_signal_7278, new_AGEMA_signal_7277, new_AGEMA_signal_7276, KeyExpansionOutput[17]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U55 ( .a ({new_AGEMA_signal_15241, new_AGEMA_signal_15237, new_AGEMA_signal_15233, new_AGEMA_signal_15229}), .b ({new_AGEMA_signal_6363, new_AGEMA_signal_6362, new_AGEMA_signal_6361, KeyExpansionOutput[81]}), .c ({new_AGEMA_signal_6801, new_AGEMA_signal_6800, new_AGEMA_signal_6799, KeyExpansionOutput[49]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U54 ( .a ({new_AGEMA_signal_15257, new_AGEMA_signal_15253, new_AGEMA_signal_15249, new_AGEMA_signal_15245}), .b ({new_AGEMA_signal_6132, new_AGEMA_signal_6131, new_AGEMA_signal_6130, KeyExpansionOutput[113]}), .c ({new_AGEMA_signal_6363, new_AGEMA_signal_6362, new_AGEMA_signal_6361, KeyExpansionOutput[81]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U53 ( .a ({new_AGEMA_signal_15273, new_AGEMA_signal_15269, new_AGEMA_signal_15265, new_AGEMA_signal_15261}), .b ({new_AGEMA_signal_6366, new_AGEMA_signal_6365, new_AGEMA_signal_6364, KeyExpansionOutput[48]}), .c ({new_AGEMA_signal_6804, new_AGEMA_signal_6803, new_AGEMA_signal_6802, KeyExpansionOutput[16]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U52 ( .a ({new_AGEMA_signal_15289, new_AGEMA_signal_15285, new_AGEMA_signal_15281, new_AGEMA_signal_15277}), .b ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, new_AGEMA_signal_6106, KeyExpansionOutput[80]}), .c ({new_AGEMA_signal_6366, new_AGEMA_signal_6365, new_AGEMA_signal_6364, KeyExpansionOutput[48]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U51 ( .a ({new_AGEMA_signal_15305, new_AGEMA_signal_15301, new_AGEMA_signal_15297, new_AGEMA_signal_15293}), .b ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, new_AGEMA_signal_5986, KeyExpansionOutput[112]}), .c ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, new_AGEMA_signal_6106, KeyExpansionOutput[80]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U50 ( .a ({new_AGEMA_signal_15321, new_AGEMA_signal_15317, new_AGEMA_signal_15313, new_AGEMA_signal_15309}), .b ({new_AGEMA_signal_6807, new_AGEMA_signal_6806, new_AGEMA_signal_6805, KeyExpansionOutput[47]}), .c ({new_AGEMA_signal_7281, new_AGEMA_signal_7280, new_AGEMA_signal_7279, KeyExpansionOutput[15]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U49 ( .a ({new_AGEMA_signal_15337, new_AGEMA_signal_15333, new_AGEMA_signal_15329, new_AGEMA_signal_15325}), .b ({new_AGEMA_signal_6369, new_AGEMA_signal_6368, new_AGEMA_signal_6367, KeyExpansionOutput[79]}), .c ({new_AGEMA_signal_6807, new_AGEMA_signal_6806, new_AGEMA_signal_6805, KeyExpansionOutput[47]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U48 ( .a ({new_AGEMA_signal_15353, new_AGEMA_signal_15349, new_AGEMA_signal_15345, new_AGEMA_signal_15341}), .b ({new_AGEMA_signal_6135, new_AGEMA_signal_6134, new_AGEMA_signal_6133, KeyExpansionOutput[111]}), .c ({new_AGEMA_signal_6369, new_AGEMA_signal_6368, new_AGEMA_signal_6367, KeyExpansionOutput[79]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U47 ( .a ({new_AGEMA_signal_15369, new_AGEMA_signal_15365, new_AGEMA_signal_15361, new_AGEMA_signal_15357}), .b ({new_AGEMA_signal_6810, new_AGEMA_signal_6809, new_AGEMA_signal_6808, KeyExpansionOutput[46]}), .c ({new_AGEMA_signal_7284, new_AGEMA_signal_7283, new_AGEMA_signal_7282, KeyExpansionOutput[14]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U46 ( .a ({new_AGEMA_signal_15385, new_AGEMA_signal_15381, new_AGEMA_signal_15377, new_AGEMA_signal_15373}), .b ({new_AGEMA_signal_6372, new_AGEMA_signal_6371, new_AGEMA_signal_6370, KeyExpansionOutput[78]}), .c ({new_AGEMA_signal_6810, new_AGEMA_signal_6809, new_AGEMA_signal_6808, KeyExpansionOutput[46]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U45 ( .a ({new_AGEMA_signal_15401, new_AGEMA_signal_15397, new_AGEMA_signal_15393, new_AGEMA_signal_15389}), .b ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, new_AGEMA_signal_6136, KeyExpansionOutput[110]}), .c ({new_AGEMA_signal_6372, new_AGEMA_signal_6371, new_AGEMA_signal_6370, KeyExpansionOutput[78]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U44 ( .a ({new_AGEMA_signal_15417, new_AGEMA_signal_15413, new_AGEMA_signal_15409, new_AGEMA_signal_15405}), .b ({new_AGEMA_signal_6813, new_AGEMA_signal_6812, new_AGEMA_signal_6811, KeyExpansionOutput[45]}), .c ({new_AGEMA_signal_7287, new_AGEMA_signal_7286, new_AGEMA_signal_7285, KeyExpansionOutput[13]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U43 ( .a ({new_AGEMA_signal_15433, new_AGEMA_signal_15429, new_AGEMA_signal_15425, new_AGEMA_signal_15421}), .b ({new_AGEMA_signal_6375, new_AGEMA_signal_6374, new_AGEMA_signal_6373, KeyExpansionOutput[77]}), .c ({new_AGEMA_signal_6813, new_AGEMA_signal_6812, new_AGEMA_signal_6811, KeyExpansionOutput[45]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U42 ( .a ({new_AGEMA_signal_15449, new_AGEMA_signal_15445, new_AGEMA_signal_15441, new_AGEMA_signal_15437}), .b ({new_AGEMA_signal_6141, new_AGEMA_signal_6140, new_AGEMA_signal_6139, KeyExpansionOutput[109]}), .c ({new_AGEMA_signal_6375, new_AGEMA_signal_6374, new_AGEMA_signal_6373, KeyExpansionOutput[77]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U41 ( .a ({new_AGEMA_signal_15465, new_AGEMA_signal_15461, new_AGEMA_signal_15457, new_AGEMA_signal_15453}), .b ({new_AGEMA_signal_6816, new_AGEMA_signal_6815, new_AGEMA_signal_6814, KeyExpansionOutput[44]}), .c ({new_AGEMA_signal_7290, new_AGEMA_signal_7289, new_AGEMA_signal_7288, KeyExpansionOutput[12]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U40 ( .a ({new_AGEMA_signal_15481, new_AGEMA_signal_15477, new_AGEMA_signal_15473, new_AGEMA_signal_15469}), .b ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, new_AGEMA_signal_6376, KeyExpansionOutput[76]}), .c ({new_AGEMA_signal_6816, new_AGEMA_signal_6815, new_AGEMA_signal_6814, KeyExpansionOutput[44]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U39 ( .a ({new_AGEMA_signal_15497, new_AGEMA_signal_15493, new_AGEMA_signal_15489, new_AGEMA_signal_15485}), .b ({new_AGEMA_signal_6144, new_AGEMA_signal_6143, new_AGEMA_signal_6142, KeyExpansionOutput[108]}), .c ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, new_AGEMA_signal_6376, KeyExpansionOutput[76]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U38 ( .a ({new_AGEMA_signal_15513, new_AGEMA_signal_15509, new_AGEMA_signal_15505, new_AGEMA_signal_15501}), .b ({new_AGEMA_signal_6171, new_AGEMA_signal_6170, new_AGEMA_signal_6169, KeyExpansionIns_tmp[31]}), .c ({new_AGEMA_signal_6381, new_AGEMA_signal_6380, new_AGEMA_signal_6379, KeyExpansionOutput[127]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U37 ( .a ({new_AGEMA_signal_15529, new_AGEMA_signal_15525, new_AGEMA_signal_15521, new_AGEMA_signal_15517}), .b ({new_AGEMA_signal_6174, new_AGEMA_signal_6173, new_AGEMA_signal_6172, KeyExpansionIns_tmp[30]}), .c ({new_AGEMA_signal_6384, new_AGEMA_signal_6383, new_AGEMA_signal_6382, KeyExpansionOutput[126]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U36 ( .a ({new_AGEMA_signal_15545, new_AGEMA_signal_15541, new_AGEMA_signal_15537, new_AGEMA_signal_15533}), .b ({new_AGEMA_signal_6177, new_AGEMA_signal_6176, new_AGEMA_signal_6175, KeyExpansionIns_tmp[29]}), .c ({new_AGEMA_signal_6387, new_AGEMA_signal_6386, new_AGEMA_signal_6385, KeyExpansionOutput[125]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U35 ( .a ({new_AGEMA_signal_15561, new_AGEMA_signal_15557, new_AGEMA_signal_15553, new_AGEMA_signal_15549}), .b ({new_AGEMA_signal_6180, new_AGEMA_signal_6179, new_AGEMA_signal_6178, KeyExpansionIns_tmp[28]}), .c ({new_AGEMA_signal_6390, new_AGEMA_signal_6389, new_AGEMA_signal_6388, KeyExpansionOutput[124]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U34 ( .a ({new_AGEMA_signal_15577, new_AGEMA_signal_15573, new_AGEMA_signal_15569, new_AGEMA_signal_15565}), .b ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, new_AGEMA_signal_6181, KeyExpansionIns_tmp[27]}), .c ({new_AGEMA_signal_6393, new_AGEMA_signal_6392, new_AGEMA_signal_6391, KeyExpansionOutput[123]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U33 ( .a ({new_AGEMA_signal_15593, new_AGEMA_signal_15589, new_AGEMA_signal_15585, new_AGEMA_signal_15581}), .b ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, new_AGEMA_signal_6184, KeyExpansionIns_tmp[26]}), .c ({new_AGEMA_signal_6396, new_AGEMA_signal_6395, new_AGEMA_signal_6394, KeyExpansionOutput[122]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U32 ( .a ({new_AGEMA_signal_15609, new_AGEMA_signal_15605, new_AGEMA_signal_15601, new_AGEMA_signal_15597}), .b ({new_AGEMA_signal_6189, new_AGEMA_signal_6188, new_AGEMA_signal_6187, KeyExpansionIns_tmp[25]}), .c ({new_AGEMA_signal_6399, new_AGEMA_signal_6398, new_AGEMA_signal_6397, KeyExpansionOutput[121]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U31 ( .a ({new_AGEMA_signal_15625, new_AGEMA_signal_15621, new_AGEMA_signal_15617, new_AGEMA_signal_15613}), .b ({new_AGEMA_signal_5997, new_AGEMA_signal_5996, new_AGEMA_signal_5995, KeyExpansionIns_tmp[24]}), .c ({new_AGEMA_signal_6111, new_AGEMA_signal_6110, new_AGEMA_signal_6109, KeyExpansionOutput[120]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U30 ( .a ({new_AGEMA_signal_15641, new_AGEMA_signal_15637, new_AGEMA_signal_15633, new_AGEMA_signal_15629}), .b ({new_AGEMA_signal_6819, new_AGEMA_signal_6818, new_AGEMA_signal_6817, KeyExpansionOutput[43]}), .c ({new_AGEMA_signal_7293, new_AGEMA_signal_7292, new_AGEMA_signal_7291, KeyExpansionOutput[11]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U29 ( .a ({new_AGEMA_signal_15657, new_AGEMA_signal_15653, new_AGEMA_signal_15649, new_AGEMA_signal_15645}), .b ({new_AGEMA_signal_6402, new_AGEMA_signal_6401, new_AGEMA_signal_6400, KeyExpansionOutput[75]}), .c ({new_AGEMA_signal_6819, new_AGEMA_signal_6818, new_AGEMA_signal_6817, KeyExpansionOutput[43]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U28 ( .a ({new_AGEMA_signal_15673, new_AGEMA_signal_15669, new_AGEMA_signal_15665, new_AGEMA_signal_15661}), .b ({new_AGEMA_signal_6147, new_AGEMA_signal_6146, new_AGEMA_signal_6145, KeyExpansionOutput[107]}), .c ({new_AGEMA_signal_6402, new_AGEMA_signal_6401, new_AGEMA_signal_6400, KeyExpansionOutput[75]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U27 ( .a ({new_AGEMA_signal_15689, new_AGEMA_signal_15685, new_AGEMA_signal_15681, new_AGEMA_signal_15677}), .b ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_6114, new_AGEMA_signal_6113, new_AGEMA_signal_6112, KeyExpansionOutput[119]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U26 ( .a ({new_AGEMA_signal_15705, new_AGEMA_signal_15701, new_AGEMA_signal_15697, new_AGEMA_signal_15693}), .b ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, new_AGEMA_signal_5926, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_6117, new_AGEMA_signal_6116, new_AGEMA_signal_6115, KeyExpansionOutput[118]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U25 ( .a ({new_AGEMA_signal_15721, new_AGEMA_signal_15717, new_AGEMA_signal_15713, new_AGEMA_signal_15709}), .b ({new_AGEMA_signal_5931, new_AGEMA_signal_5930, new_AGEMA_signal_5929, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_6120, new_AGEMA_signal_6119, new_AGEMA_signal_6118, KeyExpansionOutput[117]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U24 ( .a ({new_AGEMA_signal_15737, new_AGEMA_signal_15733, new_AGEMA_signal_15729, new_AGEMA_signal_15725}), .b ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, new_AGEMA_signal_5932, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, new_AGEMA_signal_6121, KeyExpansionOutput[116]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U23 ( .a ({new_AGEMA_signal_15753, new_AGEMA_signal_15749, new_AGEMA_signal_15745, new_AGEMA_signal_15741}), .b ({new_AGEMA_signal_5937, new_AGEMA_signal_5936, new_AGEMA_signal_5935, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, new_AGEMA_signal_6124, KeyExpansionOutput[115]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U22 ( .a ({new_AGEMA_signal_15769, new_AGEMA_signal_15765, new_AGEMA_signal_15761, new_AGEMA_signal_15757}), .b ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, new_AGEMA_signal_5938, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_6129, new_AGEMA_signal_6128, new_AGEMA_signal_6127, KeyExpansionOutput[114]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U21 ( .a ({new_AGEMA_signal_15785, new_AGEMA_signal_15781, new_AGEMA_signal_15777, new_AGEMA_signal_15773}), .b ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_6132, new_AGEMA_signal_6131, new_AGEMA_signal_6130, KeyExpansionOutput[113]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U20 ( .a ({new_AGEMA_signal_15801, new_AGEMA_signal_15797, new_AGEMA_signal_15793, new_AGEMA_signal_15789}), .b ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, new_AGEMA_signal_5833, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, new_AGEMA_signal_5986, KeyExpansionOutput[112]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U19 ( .a ({new_AGEMA_signal_15817, new_AGEMA_signal_15813, new_AGEMA_signal_15809, new_AGEMA_signal_15805}), .b ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_6135, new_AGEMA_signal_6134, new_AGEMA_signal_6133, KeyExpansionOutput[111]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U18 ( .a ({new_AGEMA_signal_15833, new_AGEMA_signal_15829, new_AGEMA_signal_15825, new_AGEMA_signal_15821}), .b ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, new_AGEMA_signal_5947, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, new_AGEMA_signal_6136, KeyExpansionOutput[110]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U17 ( .a ({new_AGEMA_signal_15849, new_AGEMA_signal_15845, new_AGEMA_signal_15841, new_AGEMA_signal_15837}), .b ({new_AGEMA_signal_6822, new_AGEMA_signal_6821, new_AGEMA_signal_6820, KeyExpansionOutput[42]}), .c ({new_AGEMA_signal_7296, new_AGEMA_signal_7295, new_AGEMA_signal_7294, KeyExpansionOutput[10]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U16 ( .a ({new_AGEMA_signal_15865, new_AGEMA_signal_15861, new_AGEMA_signal_15857, new_AGEMA_signal_15853}), .b ({new_AGEMA_signal_6405, new_AGEMA_signal_6404, new_AGEMA_signal_6403, KeyExpansionOutput[74]}), .c ({new_AGEMA_signal_6822, new_AGEMA_signal_6821, new_AGEMA_signal_6820, KeyExpansionOutput[42]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U15 ( .a ({new_AGEMA_signal_15881, new_AGEMA_signal_15877, new_AGEMA_signal_15873, new_AGEMA_signal_15869}), .b ({new_AGEMA_signal_6150, new_AGEMA_signal_6149, new_AGEMA_signal_6148, KeyExpansionOutput[106]}), .c ({new_AGEMA_signal_6405, new_AGEMA_signal_6404, new_AGEMA_signal_6403, KeyExpansionOutput[74]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U14 ( .a ({new_AGEMA_signal_15897, new_AGEMA_signal_15893, new_AGEMA_signal_15889, new_AGEMA_signal_15885}), .b ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, new_AGEMA_signal_5950, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_6141, new_AGEMA_signal_6140, new_AGEMA_signal_6139, KeyExpansionOutput[109]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U13 ( .a ({new_AGEMA_signal_15913, new_AGEMA_signal_15909, new_AGEMA_signal_15905, new_AGEMA_signal_15901}), .b ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, new_AGEMA_signal_5953, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_6144, new_AGEMA_signal_6143, new_AGEMA_signal_6142, KeyExpansionOutput[108]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U12 ( .a ({new_AGEMA_signal_15929, new_AGEMA_signal_15925, new_AGEMA_signal_15921, new_AGEMA_signal_15917}), .b ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, new_AGEMA_signal_5956, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_6147, new_AGEMA_signal_6146, new_AGEMA_signal_6145, KeyExpansionOutput[107]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U11 ( .a ({new_AGEMA_signal_15945, new_AGEMA_signal_15941, new_AGEMA_signal_15937, new_AGEMA_signal_15933}), .b ({new_AGEMA_signal_5961, new_AGEMA_signal_5960, new_AGEMA_signal_5959, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_6150, new_AGEMA_signal_6149, new_AGEMA_signal_6148, KeyExpansionOutput[106]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U10 ( .a ({new_AGEMA_signal_15961, new_AGEMA_signal_15957, new_AGEMA_signal_15953, new_AGEMA_signal_15949}), .b ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, new_AGEMA_signal_5962, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_6153, new_AGEMA_signal_6152, new_AGEMA_signal_6151, KeyExpansionOutput[105]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U9 ( .a ({new_AGEMA_signal_15977, new_AGEMA_signal_15973, new_AGEMA_signal_15969, new_AGEMA_signal_15965}), .b ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, new_AGEMA_signal_5866, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_5991, new_AGEMA_signal_5990, new_AGEMA_signal_5989, KeyExpansionOutput[104]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U8 ( .a ({new_AGEMA_signal_15993, new_AGEMA_signal_15989, new_AGEMA_signal_15985, new_AGEMA_signal_15981}), .b ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, new_AGEMA_signal_5965, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, new_AGEMA_signal_6154, KeyExpansionOutput[103]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U7 ( .a ({new_AGEMA_signal_16009, new_AGEMA_signal_16005, new_AGEMA_signal_16001, new_AGEMA_signal_15997}), .b ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, new_AGEMA_signal_5968, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_6159, new_AGEMA_signal_6158, new_AGEMA_signal_6157, KeyExpansionOutput[102]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U6 ( .a ({new_AGEMA_signal_16025, new_AGEMA_signal_16021, new_AGEMA_signal_16017, new_AGEMA_signal_16013}), .b ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_6162, new_AGEMA_signal_6161, new_AGEMA_signal_6160, KeyExpansionOutput[101]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U5 ( .a ({new_AGEMA_signal_16041, new_AGEMA_signal_16037, new_AGEMA_signal_16033, new_AGEMA_signal_16029}), .b ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, new_AGEMA_signal_5974, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_6165, new_AGEMA_signal_6164, new_AGEMA_signal_6163, KeyExpansionOutput[100]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U4 ( .a ({new_AGEMA_signal_16057, new_AGEMA_signal_16053, new_AGEMA_signal_16049, new_AGEMA_signal_16045}), .b ({new_AGEMA_signal_6408, new_AGEMA_signal_6407, new_AGEMA_signal_6406, KeyExpansionOutput[32]}), .c ({new_AGEMA_signal_6825, new_AGEMA_signal_6824, new_AGEMA_signal_6823, KeyExpansionOutput[0]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U3 ( .a ({new_AGEMA_signal_16073, new_AGEMA_signal_16069, new_AGEMA_signal_16065, new_AGEMA_signal_16061}), .b ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, new_AGEMA_signal_6166, KeyExpansionOutput[64]}), .c ({new_AGEMA_signal_6408, new_AGEMA_signal_6407, new_AGEMA_signal_6406, KeyExpansionOutput[32]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U2 ( .a ({new_AGEMA_signal_16089, new_AGEMA_signal_16085, new_AGEMA_signal_16081, new_AGEMA_signal_16077}), .b ({new_AGEMA_signal_5994, new_AGEMA_signal_5993, new_AGEMA_signal_5992, KeyExpansionOutput[96]}), .c ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, new_AGEMA_signal_6166, KeyExpansionOutput[64]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_U1 ( .a ({new_AGEMA_signal_16105, new_AGEMA_signal_16101, new_AGEMA_signal_16097, new_AGEMA_signal_16093}), .b ({new_AGEMA_signal_5901, new_AGEMA_signal_5900, new_AGEMA_signal_5899, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_5994, new_AGEMA_signal_5993, new_AGEMA_signal_5992, KeyExpansionOutput[96]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U8 ( .a ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_16109}), .b ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, new_AGEMA_signal_5902, MixColumnsIns_DoubleBytes[0]}), .c ({new_AGEMA_signal_6171, new_AGEMA_signal_6170, new_AGEMA_signal_6169, KeyExpansionIns_tmp[31]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U7 ( .a ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_16113}), .b ({new_AGEMA_signal_5907, new_AGEMA_signal_5906, new_AGEMA_signal_5905, MixColumnsIns_DoubleBytes[7]}), .c ({new_AGEMA_signal_6174, new_AGEMA_signal_6173, new_AGEMA_signal_6172, KeyExpansionIns_tmp[30]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U6 ( .a ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_16117}), .b ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, new_AGEMA_signal_5908, MixColumnsIns_DoubleBytes[6]}), .c ({new_AGEMA_signal_6177, new_AGEMA_signal_6176, new_AGEMA_signal_6175, KeyExpansionIns_tmp[29]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U5 ( .a ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_16121}), .b ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, MixColumnsIns_DoubleBytes[5]}), .c ({new_AGEMA_signal_6180, new_AGEMA_signal_6179, new_AGEMA_signal_6178, KeyExpansionIns_tmp[28]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U4 ( .a ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_16125}), .b ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, new_AGEMA_signal_5914, SubBytesOutput[3]}), .c ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, new_AGEMA_signal_6181, KeyExpansionIns_tmp[27]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U3 ( .a ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_16129}), .b ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesOutput[2]}), .c ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, new_AGEMA_signal_6184, KeyExpansionIns_tmp[26]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U2 ( .a ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_16133}), .b ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, new_AGEMA_signal_5920, MixColumnsIns_DoubleBytes[2]}), .c ({new_AGEMA_signal_6189, new_AGEMA_signal_6188, new_AGEMA_signal_6187, KeyExpansionIns_tmp[25]}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U1 ( .a ({1'b0, 1'b0, 1'b0, new_AGEMA_signal_16137}), .b ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, new_AGEMA_signal_5800, SubBytesOutput[0]}), .c ({new_AGEMA_signal_5997, new_AGEMA_signal_5996, new_AGEMA_signal_5995, KeyExpansionIns_tmp[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_0_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_16057, new_AGEMA_signal_16053, new_AGEMA_signal_16049, new_AGEMA_signal_16045}), .a ({new_AGEMA_signal_6825, new_AGEMA_signal_6824, new_AGEMA_signal_6823, KeyExpansionOutput[0]}), .c ({new_AGEMA_signal_7299, new_AGEMA_signal_7298, new_AGEMA_signal_7297, RoundKeyOutput[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_1_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_15065, new_AGEMA_signal_15061, new_AGEMA_signal_15057, new_AGEMA_signal_15053}), .a ({new_AGEMA_signal_7269, new_AGEMA_signal_7268, new_AGEMA_signal_7267, KeyExpansionOutput[1]}), .c ({new_AGEMA_signal_7704, new_AGEMA_signal_7703, new_AGEMA_signal_7702, RoundKeyOutput[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_2_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_14521, new_AGEMA_signal_14517, new_AGEMA_signal_14513, new_AGEMA_signal_14509}), .a ({new_AGEMA_signal_7236, new_AGEMA_signal_7235, new_AGEMA_signal_7234, KeyExpansionOutput[2]}), .c ({new_AGEMA_signal_7707, new_AGEMA_signal_7706, new_AGEMA_signal_7705, RoundKeyOutput[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_3_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_14233, new_AGEMA_signal_14229, new_AGEMA_signal_14225, new_AGEMA_signal_14221}), .a ({new_AGEMA_signal_7227, new_AGEMA_signal_7226, new_AGEMA_signal_7225, KeyExpansionOutput[3]}), .c ({new_AGEMA_signal_7710, new_AGEMA_signal_7709, new_AGEMA_signal_7708, RoundKeyOutput[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_4_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_14153, new_AGEMA_signal_14149, new_AGEMA_signal_14145, new_AGEMA_signal_14141}), .a ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, new_AGEMA_signal_7222, KeyExpansionOutput[4]}), .c ({new_AGEMA_signal_7713, new_AGEMA_signal_7712, new_AGEMA_signal_7711, RoundKeyOutput[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_5_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_14137, new_AGEMA_signal_14133, new_AGEMA_signal_14129, new_AGEMA_signal_14125}), .a ({new_AGEMA_signal_7221, new_AGEMA_signal_7220, new_AGEMA_signal_7219, KeyExpansionOutput[5]}), .c ({new_AGEMA_signal_7716, new_AGEMA_signal_7715, new_AGEMA_signal_7714, RoundKeyOutput[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_6_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_14121, new_AGEMA_signal_14117, new_AGEMA_signal_14113, new_AGEMA_signal_14109}), .a ({new_AGEMA_signal_7218, new_AGEMA_signal_7217, new_AGEMA_signal_7216, KeyExpansionOutput[6]}), .c ({new_AGEMA_signal_7719, new_AGEMA_signal_7718, new_AGEMA_signal_7717, RoundKeyOutput[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_7_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_14105, new_AGEMA_signal_14101, new_AGEMA_signal_14097, new_AGEMA_signal_14093}), .a ({new_AGEMA_signal_7215, new_AGEMA_signal_7214, new_AGEMA_signal_7213, KeyExpansionOutput[7]}), .c ({new_AGEMA_signal_7722, new_AGEMA_signal_7721, new_AGEMA_signal_7720, RoundKeyOutput[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_8_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_14089, new_AGEMA_signal_14085, new_AGEMA_signal_14081, new_AGEMA_signal_14077}), .a ({new_AGEMA_signal_6732, new_AGEMA_signal_6731, new_AGEMA_signal_6730, KeyExpansionOutput[8]}), .c ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, new_AGEMA_signal_7300, RoundKeyOutput[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_9_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_14073, new_AGEMA_signal_14069, new_AGEMA_signal_14065, new_AGEMA_signal_14061}), .a ({new_AGEMA_signal_7212, new_AGEMA_signal_7211, new_AGEMA_signal_7210, KeyExpansionOutput[9]}), .c ({new_AGEMA_signal_7725, new_AGEMA_signal_7724, new_AGEMA_signal_7723, RoundKeyOutput[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_10_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_15849, new_AGEMA_signal_15845, new_AGEMA_signal_15841, new_AGEMA_signal_15837}), .a ({new_AGEMA_signal_7296, new_AGEMA_signal_7295, new_AGEMA_signal_7294, KeyExpansionOutput[10]}), .c ({new_AGEMA_signal_7728, new_AGEMA_signal_7727, new_AGEMA_signal_7726, RoundKeyOutput[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_11_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_15641, new_AGEMA_signal_15637, new_AGEMA_signal_15633, new_AGEMA_signal_15629}), .a ({new_AGEMA_signal_7293, new_AGEMA_signal_7292, new_AGEMA_signal_7291, KeyExpansionOutput[11]}), .c ({new_AGEMA_signal_7731, new_AGEMA_signal_7730, new_AGEMA_signal_7729, RoundKeyOutput[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_12_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_15465, new_AGEMA_signal_15461, new_AGEMA_signal_15457, new_AGEMA_signal_15453}), .a ({new_AGEMA_signal_7290, new_AGEMA_signal_7289, new_AGEMA_signal_7288, KeyExpansionOutput[12]}), .c ({new_AGEMA_signal_7734, new_AGEMA_signal_7733, new_AGEMA_signal_7732, RoundKeyOutput[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_13_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_15417, new_AGEMA_signal_15413, new_AGEMA_signal_15409, new_AGEMA_signal_15405}), .a ({new_AGEMA_signal_7287, new_AGEMA_signal_7286, new_AGEMA_signal_7285, KeyExpansionOutput[13]}), .c ({new_AGEMA_signal_7737, new_AGEMA_signal_7736, new_AGEMA_signal_7735, RoundKeyOutput[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_14_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_15369, new_AGEMA_signal_15365, new_AGEMA_signal_15361, new_AGEMA_signal_15357}), .a ({new_AGEMA_signal_7284, new_AGEMA_signal_7283, new_AGEMA_signal_7282, KeyExpansionOutput[14]}), .c ({new_AGEMA_signal_7740, new_AGEMA_signal_7739, new_AGEMA_signal_7738, RoundKeyOutput[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_15_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_15321, new_AGEMA_signal_15317, new_AGEMA_signal_15313, new_AGEMA_signal_15309}), .a ({new_AGEMA_signal_7281, new_AGEMA_signal_7280, new_AGEMA_signal_7279, KeyExpansionOutput[15]}), .c ({new_AGEMA_signal_7743, new_AGEMA_signal_7742, new_AGEMA_signal_7741, RoundKeyOutput[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_16_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_15273, new_AGEMA_signal_15269, new_AGEMA_signal_15265, new_AGEMA_signal_15261}), .a ({new_AGEMA_signal_6804, new_AGEMA_signal_6803, new_AGEMA_signal_6802, KeyExpansionOutput[16]}), .c ({new_AGEMA_signal_7305, new_AGEMA_signal_7304, new_AGEMA_signal_7303, RoundKeyOutput[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_17_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_15225, new_AGEMA_signal_15221, new_AGEMA_signal_15217, new_AGEMA_signal_15213}), .a ({new_AGEMA_signal_7278, new_AGEMA_signal_7277, new_AGEMA_signal_7276, KeyExpansionOutput[17]}), .c ({new_AGEMA_signal_7746, new_AGEMA_signal_7745, new_AGEMA_signal_7744, RoundKeyOutput[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_18_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_15177, new_AGEMA_signal_15173, new_AGEMA_signal_15169, new_AGEMA_signal_15165}), .a ({new_AGEMA_signal_7275, new_AGEMA_signal_7274, new_AGEMA_signal_7273, KeyExpansionOutput[18]}), .c ({new_AGEMA_signal_7749, new_AGEMA_signal_7748, new_AGEMA_signal_7747, RoundKeyOutput[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_19_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_15129, new_AGEMA_signal_15125, new_AGEMA_signal_15121, new_AGEMA_signal_15117}), .a ({new_AGEMA_signal_7272, new_AGEMA_signal_7271, new_AGEMA_signal_7270, KeyExpansionOutput[19]}), .c ({new_AGEMA_signal_7752, new_AGEMA_signal_7751, new_AGEMA_signal_7750, RoundKeyOutput[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_20_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_15017, new_AGEMA_signal_15013, new_AGEMA_signal_15009, new_AGEMA_signal_15005}), .a ({new_AGEMA_signal_7266, new_AGEMA_signal_7265, new_AGEMA_signal_7264, KeyExpansionOutput[20]}), .c ({new_AGEMA_signal_7755, new_AGEMA_signal_7754, new_AGEMA_signal_7753, RoundKeyOutput[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_21_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_14969, new_AGEMA_signal_14965, new_AGEMA_signal_14961, new_AGEMA_signal_14957}), .a ({new_AGEMA_signal_7263, new_AGEMA_signal_7262, new_AGEMA_signal_7261, KeyExpansionOutput[21]}), .c ({new_AGEMA_signal_7758, new_AGEMA_signal_7757, new_AGEMA_signal_7756, RoundKeyOutput[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_22_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_14921, new_AGEMA_signal_14917, new_AGEMA_signal_14913, new_AGEMA_signal_14909}), .a ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, new_AGEMA_signal_7258, KeyExpansionOutput[22]}), .c ({new_AGEMA_signal_7761, new_AGEMA_signal_7760, new_AGEMA_signal_7759, RoundKeyOutput[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_23_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_14873, new_AGEMA_signal_14869, new_AGEMA_signal_14865, new_AGEMA_signal_14861}), .a ({new_AGEMA_signal_7257, new_AGEMA_signal_7256, new_AGEMA_signal_7255, KeyExpansionOutput[23]}), .c ({new_AGEMA_signal_7764, new_AGEMA_signal_7763, new_AGEMA_signal_7762, RoundKeyOutput[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_24_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_14825, new_AGEMA_signal_14821, new_AGEMA_signal_14817, new_AGEMA_signal_14813}), .a ({new_AGEMA_signal_7254, new_AGEMA_signal_7253, new_AGEMA_signal_7252, KeyExpansionOutput[24]}), .c ({new_AGEMA_signal_7767, new_AGEMA_signal_7766, new_AGEMA_signal_7765, RoundKeyOutput[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_25_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_14777, new_AGEMA_signal_14773, new_AGEMA_signal_14769, new_AGEMA_signal_14765}), .a ({new_AGEMA_signal_7701, new_AGEMA_signal_7700, new_AGEMA_signal_7699, KeyExpansionOutput[25]}), .c ({new_AGEMA_signal_8121, new_AGEMA_signal_8120, new_AGEMA_signal_8119, RoundKeyOutput[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_26_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_14729, new_AGEMA_signal_14725, new_AGEMA_signal_14721, new_AGEMA_signal_14717}), .a ({new_AGEMA_signal_7698, new_AGEMA_signal_7697, new_AGEMA_signal_7696, KeyExpansionOutput[26]}), .c ({new_AGEMA_signal_8124, new_AGEMA_signal_8123, new_AGEMA_signal_8122, RoundKeyOutput[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_27_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_14681, new_AGEMA_signal_14677, new_AGEMA_signal_14673, new_AGEMA_signal_14669}), .a ({new_AGEMA_signal_7695, new_AGEMA_signal_7694, new_AGEMA_signal_7693, KeyExpansionOutput[27]}), .c ({new_AGEMA_signal_8127, new_AGEMA_signal_8126, new_AGEMA_signal_8125, RoundKeyOutput[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_28_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_14633, new_AGEMA_signal_14629, new_AGEMA_signal_14625, new_AGEMA_signal_14621}), .a ({new_AGEMA_signal_7692, new_AGEMA_signal_7691, new_AGEMA_signal_7690, KeyExpansionOutput[28]}), .c ({new_AGEMA_signal_8130, new_AGEMA_signal_8129, new_AGEMA_signal_8128, RoundKeyOutput[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_29_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_14585, new_AGEMA_signal_14581, new_AGEMA_signal_14577, new_AGEMA_signal_14573}), .a ({new_AGEMA_signal_7689, new_AGEMA_signal_7688, new_AGEMA_signal_7687, KeyExpansionOutput[29]}), .c ({new_AGEMA_signal_8133, new_AGEMA_signal_8132, new_AGEMA_signal_8131, RoundKeyOutput[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_30_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_14473, new_AGEMA_signal_14469, new_AGEMA_signal_14465, new_AGEMA_signal_14461}), .a ({new_AGEMA_signal_7686, new_AGEMA_signal_7685, new_AGEMA_signal_7684, KeyExpansionOutput[30]}), .c ({new_AGEMA_signal_8136, new_AGEMA_signal_8135, new_AGEMA_signal_8134, RoundKeyOutput[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_31_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_14425, new_AGEMA_signal_14421, new_AGEMA_signal_14417, new_AGEMA_signal_14413}), .a ({new_AGEMA_signal_7683, new_AGEMA_signal_7682, new_AGEMA_signal_7681, KeyExpansionOutput[31]}), .c ({new_AGEMA_signal_8139, new_AGEMA_signal_8138, new_AGEMA_signal_8137, RoundKeyOutput[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_32_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_16073, new_AGEMA_signal_16069, new_AGEMA_signal_16065, new_AGEMA_signal_16061}), .a ({new_AGEMA_signal_6408, new_AGEMA_signal_6407, new_AGEMA_signal_6406, KeyExpansionOutput[32]}), .c ({new_AGEMA_signal_6828, new_AGEMA_signal_6827, new_AGEMA_signal_6826, RoundKeyOutput[32]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_33_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_15081, new_AGEMA_signal_15077, new_AGEMA_signal_15073, new_AGEMA_signal_15069}), .a ({new_AGEMA_signal_6792, new_AGEMA_signal_6791, new_AGEMA_signal_6790, KeyExpansionOutput[33]}), .c ({new_AGEMA_signal_7308, new_AGEMA_signal_7307, new_AGEMA_signal_7306, RoundKeyOutput[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_34_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_14537, new_AGEMA_signal_14533, new_AGEMA_signal_14529, new_AGEMA_signal_14525}), .a ({new_AGEMA_signal_6759, new_AGEMA_signal_6758, new_AGEMA_signal_6757, KeyExpansionOutput[34]}), .c ({new_AGEMA_signal_7311, new_AGEMA_signal_7310, new_AGEMA_signal_7309, RoundKeyOutput[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_35_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_14377, new_AGEMA_signal_14373, new_AGEMA_signal_14369, new_AGEMA_signal_14365}), .a ({new_AGEMA_signal_6750, new_AGEMA_signal_6749, new_AGEMA_signal_6748, KeyExpansionOutput[35]}), .c ({new_AGEMA_signal_7314, new_AGEMA_signal_7313, new_AGEMA_signal_7312, RoundKeyOutput[35]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_36_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_14345, new_AGEMA_signal_14341, new_AGEMA_signal_14337, new_AGEMA_signal_14333}), .a ({new_AGEMA_signal_6747, new_AGEMA_signal_6746, new_AGEMA_signal_6745, KeyExpansionOutput[36]}), .c ({new_AGEMA_signal_7317, new_AGEMA_signal_7316, new_AGEMA_signal_7315, RoundKeyOutput[36]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_37_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_14313, new_AGEMA_signal_14309, new_AGEMA_signal_14305, new_AGEMA_signal_14301}), .a ({new_AGEMA_signal_6744, new_AGEMA_signal_6743, new_AGEMA_signal_6742, KeyExpansionOutput[37]}), .c ({new_AGEMA_signal_7320, new_AGEMA_signal_7319, new_AGEMA_signal_7318, RoundKeyOutput[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_38_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_14281, new_AGEMA_signal_14277, new_AGEMA_signal_14273, new_AGEMA_signal_14269}), .a ({new_AGEMA_signal_6741, new_AGEMA_signal_6740, new_AGEMA_signal_6739, KeyExpansionOutput[38]}), .c ({new_AGEMA_signal_7323, new_AGEMA_signal_7322, new_AGEMA_signal_7321, RoundKeyOutput[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_39_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_14249, new_AGEMA_signal_14245, new_AGEMA_signal_14241, new_AGEMA_signal_14237}), .a ({new_AGEMA_signal_6738, new_AGEMA_signal_6737, new_AGEMA_signal_6736, KeyExpansionOutput[39]}), .c ({new_AGEMA_signal_7326, new_AGEMA_signal_7325, new_AGEMA_signal_7324, RoundKeyOutput[39]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_40_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_14201, new_AGEMA_signal_14197, new_AGEMA_signal_14193, new_AGEMA_signal_14189}), .a ({new_AGEMA_signal_6318, new_AGEMA_signal_6317, new_AGEMA_signal_6316, KeyExpansionOutput[40]}), .c ({new_AGEMA_signal_6831, new_AGEMA_signal_6830, new_AGEMA_signal_6829, RoundKeyOutput[40]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_41_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_14169, new_AGEMA_signal_14165, new_AGEMA_signal_14161, new_AGEMA_signal_14157}), .a ({new_AGEMA_signal_6735, new_AGEMA_signal_6734, new_AGEMA_signal_6733, KeyExpansionOutput[41]}), .c ({new_AGEMA_signal_7329, new_AGEMA_signal_7328, new_AGEMA_signal_7327, RoundKeyOutput[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_42_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_15865, new_AGEMA_signal_15861, new_AGEMA_signal_15857, new_AGEMA_signal_15853}), .a ({new_AGEMA_signal_6822, new_AGEMA_signal_6821, new_AGEMA_signal_6820, KeyExpansionOutput[42]}), .c ({new_AGEMA_signal_7332, new_AGEMA_signal_7331, new_AGEMA_signal_7330, RoundKeyOutput[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_43_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_15657, new_AGEMA_signal_15653, new_AGEMA_signal_15649, new_AGEMA_signal_15645}), .a ({new_AGEMA_signal_6819, new_AGEMA_signal_6818, new_AGEMA_signal_6817, KeyExpansionOutput[43]}), .c ({new_AGEMA_signal_7335, new_AGEMA_signal_7334, new_AGEMA_signal_7333, RoundKeyOutput[43]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_44_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_15481, new_AGEMA_signal_15477, new_AGEMA_signal_15473, new_AGEMA_signal_15469}), .a ({new_AGEMA_signal_6816, new_AGEMA_signal_6815, new_AGEMA_signal_6814, KeyExpansionOutput[44]}), .c ({new_AGEMA_signal_7338, new_AGEMA_signal_7337, new_AGEMA_signal_7336, RoundKeyOutput[44]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_45_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_15433, new_AGEMA_signal_15429, new_AGEMA_signal_15425, new_AGEMA_signal_15421}), .a ({new_AGEMA_signal_6813, new_AGEMA_signal_6812, new_AGEMA_signal_6811, KeyExpansionOutput[45]}), .c ({new_AGEMA_signal_7341, new_AGEMA_signal_7340, new_AGEMA_signal_7339, RoundKeyOutput[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_46_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_15385, new_AGEMA_signal_15381, new_AGEMA_signal_15377, new_AGEMA_signal_15373}), .a ({new_AGEMA_signal_6810, new_AGEMA_signal_6809, new_AGEMA_signal_6808, KeyExpansionOutput[46]}), .c ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, new_AGEMA_signal_7342, RoundKeyOutput[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_47_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_15337, new_AGEMA_signal_15333, new_AGEMA_signal_15329, new_AGEMA_signal_15325}), .a ({new_AGEMA_signal_6807, new_AGEMA_signal_6806, new_AGEMA_signal_6805, KeyExpansionOutput[47]}), .c ({new_AGEMA_signal_7347, new_AGEMA_signal_7346, new_AGEMA_signal_7345, RoundKeyOutput[47]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_48_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_15289, new_AGEMA_signal_15285, new_AGEMA_signal_15281, new_AGEMA_signal_15277}), .a ({new_AGEMA_signal_6366, new_AGEMA_signal_6365, new_AGEMA_signal_6364, KeyExpansionOutput[48]}), .c ({new_AGEMA_signal_6834, new_AGEMA_signal_6833, new_AGEMA_signal_6832, RoundKeyOutput[48]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_49_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_15241, new_AGEMA_signal_15237, new_AGEMA_signal_15233, new_AGEMA_signal_15229}), .a ({new_AGEMA_signal_6801, new_AGEMA_signal_6800, new_AGEMA_signal_6799, KeyExpansionOutput[49]}), .c ({new_AGEMA_signal_7350, new_AGEMA_signal_7349, new_AGEMA_signal_7348, RoundKeyOutput[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_50_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_15193, new_AGEMA_signal_15189, new_AGEMA_signal_15185, new_AGEMA_signal_15181}), .a ({new_AGEMA_signal_6798, new_AGEMA_signal_6797, new_AGEMA_signal_6796, KeyExpansionOutput[50]}), .c ({new_AGEMA_signal_7353, new_AGEMA_signal_7352, new_AGEMA_signal_7351, RoundKeyOutput[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_51_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_15145, new_AGEMA_signal_15141, new_AGEMA_signal_15137, new_AGEMA_signal_15133}), .a ({new_AGEMA_signal_6795, new_AGEMA_signal_6794, new_AGEMA_signal_6793, KeyExpansionOutput[51]}), .c ({new_AGEMA_signal_7356, new_AGEMA_signal_7355, new_AGEMA_signal_7354, RoundKeyOutput[51]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_52_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_15033, new_AGEMA_signal_15029, new_AGEMA_signal_15025, new_AGEMA_signal_15021}), .a ({new_AGEMA_signal_6789, new_AGEMA_signal_6788, new_AGEMA_signal_6787, KeyExpansionOutput[52]}), .c ({new_AGEMA_signal_7359, new_AGEMA_signal_7358, new_AGEMA_signal_7357, RoundKeyOutput[52]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_53_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_14985, new_AGEMA_signal_14981, new_AGEMA_signal_14977, new_AGEMA_signal_14973}), .a ({new_AGEMA_signal_6786, new_AGEMA_signal_6785, new_AGEMA_signal_6784, KeyExpansionOutput[53]}), .c ({new_AGEMA_signal_7362, new_AGEMA_signal_7361, new_AGEMA_signal_7360, RoundKeyOutput[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_54_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_14937, new_AGEMA_signal_14933, new_AGEMA_signal_14929, new_AGEMA_signal_14925}), .a ({new_AGEMA_signal_6783, new_AGEMA_signal_6782, new_AGEMA_signal_6781, KeyExpansionOutput[54]}), .c ({new_AGEMA_signal_7365, new_AGEMA_signal_7364, new_AGEMA_signal_7363, RoundKeyOutput[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_55_U1 ( .s (new_AGEMA_signal_16161), .b ({new_AGEMA_signal_14889, new_AGEMA_signal_14885, new_AGEMA_signal_14881, new_AGEMA_signal_14877}), .a ({new_AGEMA_signal_6780, new_AGEMA_signal_6779, new_AGEMA_signal_6778, KeyExpansionOutput[55]}), .c ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, new_AGEMA_signal_7366, RoundKeyOutput[55]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_56_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_14841, new_AGEMA_signal_14837, new_AGEMA_signal_14833, new_AGEMA_signal_14829}), .a ({new_AGEMA_signal_6777, new_AGEMA_signal_6776, new_AGEMA_signal_6775, KeyExpansionOutput[56]}), .c ({new_AGEMA_signal_7371, new_AGEMA_signal_7370, new_AGEMA_signal_7369, RoundKeyOutput[56]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_57_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_14793, new_AGEMA_signal_14789, new_AGEMA_signal_14785, new_AGEMA_signal_14781}), .a ({new_AGEMA_signal_7251, new_AGEMA_signal_7250, new_AGEMA_signal_7249, KeyExpansionOutput[57]}), .c ({new_AGEMA_signal_7770, new_AGEMA_signal_7769, new_AGEMA_signal_7768, RoundKeyOutput[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_58_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_14745, new_AGEMA_signal_14741, new_AGEMA_signal_14737, new_AGEMA_signal_14733}), .a ({new_AGEMA_signal_7248, new_AGEMA_signal_7247, new_AGEMA_signal_7246, KeyExpansionOutput[58]}), .c ({new_AGEMA_signal_7773, new_AGEMA_signal_7772, new_AGEMA_signal_7771, RoundKeyOutput[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_59_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_14697, new_AGEMA_signal_14693, new_AGEMA_signal_14689, new_AGEMA_signal_14685}), .a ({new_AGEMA_signal_7245, new_AGEMA_signal_7244, new_AGEMA_signal_7243, KeyExpansionOutput[59]}), .c ({new_AGEMA_signal_7776, new_AGEMA_signal_7775, new_AGEMA_signal_7774, RoundKeyOutput[59]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_60_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_14649, new_AGEMA_signal_14645, new_AGEMA_signal_14641, new_AGEMA_signal_14637}), .a ({new_AGEMA_signal_7242, new_AGEMA_signal_7241, new_AGEMA_signal_7240, KeyExpansionOutput[60]}), .c ({new_AGEMA_signal_7779, new_AGEMA_signal_7778, new_AGEMA_signal_7777, RoundKeyOutput[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_61_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_14601, new_AGEMA_signal_14597, new_AGEMA_signal_14593, new_AGEMA_signal_14589}), .a ({new_AGEMA_signal_7239, new_AGEMA_signal_7238, new_AGEMA_signal_7237, KeyExpansionOutput[61]}), .c ({new_AGEMA_signal_7782, new_AGEMA_signal_7781, new_AGEMA_signal_7780, RoundKeyOutput[61]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_62_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_14489, new_AGEMA_signal_14485, new_AGEMA_signal_14481, new_AGEMA_signal_14477}), .a ({new_AGEMA_signal_7233, new_AGEMA_signal_7232, new_AGEMA_signal_7231, KeyExpansionOutput[62]}), .c ({new_AGEMA_signal_7785, new_AGEMA_signal_7784, new_AGEMA_signal_7783, RoundKeyOutput[62]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_63_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_14441, new_AGEMA_signal_14437, new_AGEMA_signal_14433, new_AGEMA_signal_14429}), .a ({new_AGEMA_signal_7230, new_AGEMA_signal_7229, new_AGEMA_signal_7228, KeyExpansionOutput[63]}), .c ({new_AGEMA_signal_7788, new_AGEMA_signal_7787, new_AGEMA_signal_7786, RoundKeyOutput[63]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_64_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_16089, new_AGEMA_signal_16085, new_AGEMA_signal_16081, new_AGEMA_signal_16077}), .a ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, new_AGEMA_signal_6166, KeyExpansionOutput[64]}), .c ({new_AGEMA_signal_6411, new_AGEMA_signal_6410, new_AGEMA_signal_6409, RoundKeyOutput[64]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_65_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_15097, new_AGEMA_signal_15093, new_AGEMA_signal_15089, new_AGEMA_signal_15085}), .a ({new_AGEMA_signal_6354, new_AGEMA_signal_6353, new_AGEMA_signal_6352, KeyExpansionOutput[65]}), .c ({new_AGEMA_signal_6837, new_AGEMA_signal_6836, new_AGEMA_signal_6835, RoundKeyOutput[65]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_66_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_14553, new_AGEMA_signal_14549, new_AGEMA_signal_14545, new_AGEMA_signal_14541}), .a ({new_AGEMA_signal_6336, new_AGEMA_signal_6335, new_AGEMA_signal_6334, KeyExpansionOutput[66]}), .c ({new_AGEMA_signal_6840, new_AGEMA_signal_6839, new_AGEMA_signal_6838, RoundKeyOutput[66]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_67_U1 ( .s (new_AGEMA_signal_16157), .b ({new_AGEMA_signal_14393, new_AGEMA_signal_14389, new_AGEMA_signal_14385, new_AGEMA_signal_14381}), .a ({new_AGEMA_signal_6333, new_AGEMA_signal_6332, new_AGEMA_signal_6331, KeyExpansionOutput[67]}), .c ({new_AGEMA_signal_6843, new_AGEMA_signal_6842, new_AGEMA_signal_6841, RoundKeyOutput[67]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_68_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_14361, new_AGEMA_signal_14357, new_AGEMA_signal_14353, new_AGEMA_signal_14349}), .a ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, new_AGEMA_signal_6328, KeyExpansionOutput[68]}), .c ({new_AGEMA_signal_6846, new_AGEMA_signal_6845, new_AGEMA_signal_6844, RoundKeyOutput[68]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_69_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_14329, new_AGEMA_signal_14325, new_AGEMA_signal_14321, new_AGEMA_signal_14317}), .a ({new_AGEMA_signal_6327, new_AGEMA_signal_6326, new_AGEMA_signal_6325, KeyExpansionOutput[69]}), .c ({new_AGEMA_signal_6849, new_AGEMA_signal_6848, new_AGEMA_signal_6847, RoundKeyOutput[69]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_70_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_14297, new_AGEMA_signal_14293, new_AGEMA_signal_14289, new_AGEMA_signal_14285}), .a ({new_AGEMA_signal_6324, new_AGEMA_signal_6323, new_AGEMA_signal_6322, KeyExpansionOutput[70]}), .c ({new_AGEMA_signal_6852, new_AGEMA_signal_6851, new_AGEMA_signal_6850, RoundKeyOutput[70]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_71_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_14265, new_AGEMA_signal_14261, new_AGEMA_signal_14257, new_AGEMA_signal_14253}), .a ({new_AGEMA_signal_6321, new_AGEMA_signal_6320, new_AGEMA_signal_6319, KeyExpansionOutput[71]}), .c ({new_AGEMA_signal_6855, new_AGEMA_signal_6854, new_AGEMA_signal_6853, RoundKeyOutput[71]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_72_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_14217, new_AGEMA_signal_14213, new_AGEMA_signal_14209, new_AGEMA_signal_14205}), .a ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, new_AGEMA_signal_6094, KeyExpansionOutput[72]}), .c ({new_AGEMA_signal_6414, new_AGEMA_signal_6413, new_AGEMA_signal_6412, RoundKeyOutput[72]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_73_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_14185, new_AGEMA_signal_14181, new_AGEMA_signal_14177, new_AGEMA_signal_14173}), .a ({new_AGEMA_signal_6315, new_AGEMA_signal_6314, new_AGEMA_signal_6313, KeyExpansionOutput[73]}), .c ({new_AGEMA_signal_6858, new_AGEMA_signal_6857, new_AGEMA_signal_6856, RoundKeyOutput[73]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_74_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_15881, new_AGEMA_signal_15877, new_AGEMA_signal_15873, new_AGEMA_signal_15869}), .a ({new_AGEMA_signal_6405, new_AGEMA_signal_6404, new_AGEMA_signal_6403, KeyExpansionOutput[74]}), .c ({new_AGEMA_signal_6861, new_AGEMA_signal_6860, new_AGEMA_signal_6859, RoundKeyOutput[74]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_75_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_15673, new_AGEMA_signal_15669, new_AGEMA_signal_15665, new_AGEMA_signal_15661}), .a ({new_AGEMA_signal_6402, new_AGEMA_signal_6401, new_AGEMA_signal_6400, KeyExpansionOutput[75]}), .c ({new_AGEMA_signal_6864, new_AGEMA_signal_6863, new_AGEMA_signal_6862, RoundKeyOutput[75]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_76_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_15497, new_AGEMA_signal_15493, new_AGEMA_signal_15489, new_AGEMA_signal_15485}), .a ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, new_AGEMA_signal_6376, KeyExpansionOutput[76]}), .c ({new_AGEMA_signal_6867, new_AGEMA_signal_6866, new_AGEMA_signal_6865, RoundKeyOutput[76]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_77_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_15449, new_AGEMA_signal_15445, new_AGEMA_signal_15441, new_AGEMA_signal_15437}), .a ({new_AGEMA_signal_6375, new_AGEMA_signal_6374, new_AGEMA_signal_6373, KeyExpansionOutput[77]}), .c ({new_AGEMA_signal_6870, new_AGEMA_signal_6869, new_AGEMA_signal_6868, RoundKeyOutput[77]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_78_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_15401, new_AGEMA_signal_15397, new_AGEMA_signal_15393, new_AGEMA_signal_15389}), .a ({new_AGEMA_signal_6372, new_AGEMA_signal_6371, new_AGEMA_signal_6370, KeyExpansionOutput[78]}), .c ({new_AGEMA_signal_6873, new_AGEMA_signal_6872, new_AGEMA_signal_6871, RoundKeyOutput[78]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_79_U1 ( .s (new_AGEMA_signal_16153), .b ({new_AGEMA_signal_15353, new_AGEMA_signal_15349, new_AGEMA_signal_15345, new_AGEMA_signal_15341}), .a ({new_AGEMA_signal_6369, new_AGEMA_signal_6368, new_AGEMA_signal_6367, KeyExpansionOutput[79]}), .c ({new_AGEMA_signal_6876, new_AGEMA_signal_6875, new_AGEMA_signal_6874, RoundKeyOutput[79]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_80_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_15305, new_AGEMA_signal_15301, new_AGEMA_signal_15297, new_AGEMA_signal_15293}), .a ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, new_AGEMA_signal_6106, KeyExpansionOutput[80]}), .c ({new_AGEMA_signal_6417, new_AGEMA_signal_6416, new_AGEMA_signal_6415, RoundKeyOutput[80]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_81_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_15257, new_AGEMA_signal_15253, new_AGEMA_signal_15249, new_AGEMA_signal_15245}), .a ({new_AGEMA_signal_6363, new_AGEMA_signal_6362, new_AGEMA_signal_6361, KeyExpansionOutput[81]}), .c ({new_AGEMA_signal_6879, new_AGEMA_signal_6878, new_AGEMA_signal_6877, RoundKeyOutput[81]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_82_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_15209, new_AGEMA_signal_15205, new_AGEMA_signal_15201, new_AGEMA_signal_15197}), .a ({new_AGEMA_signal_6360, new_AGEMA_signal_6359, new_AGEMA_signal_6358, KeyExpansionOutput[82]}), .c ({new_AGEMA_signal_6882, new_AGEMA_signal_6881, new_AGEMA_signal_6880, RoundKeyOutput[82]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_83_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_15161, new_AGEMA_signal_15157, new_AGEMA_signal_15153, new_AGEMA_signal_15149}), .a ({new_AGEMA_signal_6357, new_AGEMA_signal_6356, new_AGEMA_signal_6355, KeyExpansionOutput[83]}), .c ({new_AGEMA_signal_6885, new_AGEMA_signal_6884, new_AGEMA_signal_6883, RoundKeyOutput[83]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_84_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_15049, new_AGEMA_signal_15045, new_AGEMA_signal_15041, new_AGEMA_signal_15037}), .a ({new_AGEMA_signal_6351, new_AGEMA_signal_6350, new_AGEMA_signal_6349, KeyExpansionOutput[84]}), .c ({new_AGEMA_signal_6888, new_AGEMA_signal_6887, new_AGEMA_signal_6886, RoundKeyOutput[84]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_85_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_15001, new_AGEMA_signal_14997, new_AGEMA_signal_14993, new_AGEMA_signal_14989}), .a ({new_AGEMA_signal_6348, new_AGEMA_signal_6347, new_AGEMA_signal_6346, KeyExpansionOutput[85]}), .c ({new_AGEMA_signal_6891, new_AGEMA_signal_6890, new_AGEMA_signal_6889, RoundKeyOutput[85]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_86_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_14953, new_AGEMA_signal_14949, new_AGEMA_signal_14945, new_AGEMA_signal_14941}), .a ({new_AGEMA_signal_6345, new_AGEMA_signal_6344, new_AGEMA_signal_6343, KeyExpansionOutput[86]}), .c ({new_AGEMA_signal_6894, new_AGEMA_signal_6893, new_AGEMA_signal_6892, RoundKeyOutput[86]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_87_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_14905, new_AGEMA_signal_14901, new_AGEMA_signal_14897, new_AGEMA_signal_14893}), .a ({new_AGEMA_signal_6342, new_AGEMA_signal_6341, new_AGEMA_signal_6340, KeyExpansionOutput[87]}), .c ({new_AGEMA_signal_6897, new_AGEMA_signal_6896, new_AGEMA_signal_6895, RoundKeyOutput[87]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_88_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_14857, new_AGEMA_signal_14853, new_AGEMA_signal_14849, new_AGEMA_signal_14845}), .a ({new_AGEMA_signal_6339, new_AGEMA_signal_6338, new_AGEMA_signal_6337, KeyExpansionOutput[88]}), .c ({new_AGEMA_signal_6900, new_AGEMA_signal_6899, new_AGEMA_signal_6898, RoundKeyOutput[88]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_89_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_14809, new_AGEMA_signal_14805, new_AGEMA_signal_14801, new_AGEMA_signal_14797}), .a ({new_AGEMA_signal_6774, new_AGEMA_signal_6773, new_AGEMA_signal_6772, KeyExpansionOutput[89]}), .c ({new_AGEMA_signal_7374, new_AGEMA_signal_7373, new_AGEMA_signal_7372, RoundKeyOutput[89]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_90_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_14761, new_AGEMA_signal_14757, new_AGEMA_signal_14753, new_AGEMA_signal_14749}), .a ({new_AGEMA_signal_6771, new_AGEMA_signal_6770, new_AGEMA_signal_6769, KeyExpansionOutput[90]}), .c ({new_AGEMA_signal_7377, new_AGEMA_signal_7376, new_AGEMA_signal_7375, RoundKeyOutput[90]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_91_U1 ( .s (new_AGEMA_signal_16149), .b ({new_AGEMA_signal_14713, new_AGEMA_signal_14709, new_AGEMA_signal_14705, new_AGEMA_signal_14701}), .a ({new_AGEMA_signal_6768, new_AGEMA_signal_6767, new_AGEMA_signal_6766, KeyExpansionOutput[91]}), .c ({new_AGEMA_signal_7380, new_AGEMA_signal_7379, new_AGEMA_signal_7378, RoundKeyOutput[91]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_92_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_14665, new_AGEMA_signal_14661, new_AGEMA_signal_14657, new_AGEMA_signal_14653}), .a ({new_AGEMA_signal_6765, new_AGEMA_signal_6764, new_AGEMA_signal_6763, KeyExpansionOutput[92]}), .c ({new_AGEMA_signal_7383, new_AGEMA_signal_7382, new_AGEMA_signal_7381, RoundKeyOutput[92]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_93_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_14617, new_AGEMA_signal_14613, new_AGEMA_signal_14609, new_AGEMA_signal_14605}), .a ({new_AGEMA_signal_6762, new_AGEMA_signal_6761, new_AGEMA_signal_6760, KeyExpansionOutput[93]}), .c ({new_AGEMA_signal_7386, new_AGEMA_signal_7385, new_AGEMA_signal_7384, RoundKeyOutput[93]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_94_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_14505, new_AGEMA_signal_14501, new_AGEMA_signal_14497, new_AGEMA_signal_14493}), .a ({new_AGEMA_signal_6756, new_AGEMA_signal_6755, new_AGEMA_signal_6754, KeyExpansionOutput[94]}), .c ({new_AGEMA_signal_7389, new_AGEMA_signal_7388, new_AGEMA_signal_7387, RoundKeyOutput[94]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_95_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_14457, new_AGEMA_signal_14453, new_AGEMA_signal_14449, new_AGEMA_signal_14445}), .a ({new_AGEMA_signal_6753, new_AGEMA_signal_6752, new_AGEMA_signal_6751, KeyExpansionOutput[95]}), .c ({new_AGEMA_signal_7392, new_AGEMA_signal_7391, new_AGEMA_signal_7390, RoundKeyOutput[95]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_96_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_16105, new_AGEMA_signal_16101, new_AGEMA_signal_16097, new_AGEMA_signal_16093}), .a ({new_AGEMA_signal_5994, new_AGEMA_signal_5993, new_AGEMA_signal_5992, KeyExpansionOutput[96]}), .c ({new_AGEMA_signal_6192, new_AGEMA_signal_6191, new_AGEMA_signal_6190, RoundKeyOutput[96]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_97_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_15113, new_AGEMA_signal_15109, new_AGEMA_signal_15105, new_AGEMA_signal_15101}), .a ({new_AGEMA_signal_6105, new_AGEMA_signal_6104, new_AGEMA_signal_6103, KeyExpansionOutput[97]}), .c ({new_AGEMA_signal_6420, new_AGEMA_signal_6419, new_AGEMA_signal_6418, RoundKeyOutput[97]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_98_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_14569, new_AGEMA_signal_14565, new_AGEMA_signal_14561, new_AGEMA_signal_14557}), .a ({new_AGEMA_signal_6102, new_AGEMA_signal_6101, new_AGEMA_signal_6100, KeyExpansionOutput[98]}), .c ({new_AGEMA_signal_6423, new_AGEMA_signal_6422, new_AGEMA_signal_6421, RoundKeyOutput[98]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_99_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_14409, new_AGEMA_signal_14405, new_AGEMA_signal_14401, new_AGEMA_signal_14397}), .a ({new_AGEMA_signal_6099, new_AGEMA_signal_6098, new_AGEMA_signal_6097, KeyExpansionOutput[99]}), .c ({new_AGEMA_signal_6426, new_AGEMA_signal_6425, new_AGEMA_signal_6424, RoundKeyOutput[99]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_100_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_16041, new_AGEMA_signal_16037, new_AGEMA_signal_16033, new_AGEMA_signal_16029}), .a ({new_AGEMA_signal_6165, new_AGEMA_signal_6164, new_AGEMA_signal_6163, KeyExpansionOutput[100]}), .c ({new_AGEMA_signal_6429, new_AGEMA_signal_6428, new_AGEMA_signal_6427, RoundKeyOutput[100]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_101_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_16025, new_AGEMA_signal_16021, new_AGEMA_signal_16017, new_AGEMA_signal_16013}), .a ({new_AGEMA_signal_6162, new_AGEMA_signal_6161, new_AGEMA_signal_6160, KeyExpansionOutput[101]}), .c ({new_AGEMA_signal_6432, new_AGEMA_signal_6431, new_AGEMA_signal_6430, RoundKeyOutput[101]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_102_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_16009, new_AGEMA_signal_16005, new_AGEMA_signal_16001, new_AGEMA_signal_15997}), .a ({new_AGEMA_signal_6159, new_AGEMA_signal_6158, new_AGEMA_signal_6157, KeyExpansionOutput[102]}), .c ({new_AGEMA_signal_6435, new_AGEMA_signal_6434, new_AGEMA_signal_6433, RoundKeyOutput[102]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_103_U1 ( .s (new_AGEMA_signal_16145), .b ({new_AGEMA_signal_15993, new_AGEMA_signal_15989, new_AGEMA_signal_15985, new_AGEMA_signal_15981}), .a ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, new_AGEMA_signal_6154, KeyExpansionOutput[103]}), .c ({new_AGEMA_signal_6438, new_AGEMA_signal_6437, new_AGEMA_signal_6436, RoundKeyOutput[103]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_104_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_15977, new_AGEMA_signal_15973, new_AGEMA_signal_15969, new_AGEMA_signal_15965}), .a ({new_AGEMA_signal_5991, new_AGEMA_signal_5990, new_AGEMA_signal_5989, KeyExpansionOutput[104]}), .c ({new_AGEMA_signal_6195, new_AGEMA_signal_6194, new_AGEMA_signal_6193, RoundKeyOutput[104]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_105_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_15961, new_AGEMA_signal_15957, new_AGEMA_signal_15953, new_AGEMA_signal_15949}), .a ({new_AGEMA_signal_6153, new_AGEMA_signal_6152, new_AGEMA_signal_6151, KeyExpansionOutput[105]}), .c ({new_AGEMA_signal_6441, new_AGEMA_signal_6440, new_AGEMA_signal_6439, RoundKeyOutput[105]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_106_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_15945, new_AGEMA_signal_15941, new_AGEMA_signal_15937, new_AGEMA_signal_15933}), .a ({new_AGEMA_signal_6150, new_AGEMA_signal_6149, new_AGEMA_signal_6148, KeyExpansionOutput[106]}), .c ({new_AGEMA_signal_6444, new_AGEMA_signal_6443, new_AGEMA_signal_6442, RoundKeyOutput[106]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_107_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_15929, new_AGEMA_signal_15925, new_AGEMA_signal_15921, new_AGEMA_signal_15917}), .a ({new_AGEMA_signal_6147, new_AGEMA_signal_6146, new_AGEMA_signal_6145, KeyExpansionOutput[107]}), .c ({new_AGEMA_signal_6447, new_AGEMA_signal_6446, new_AGEMA_signal_6445, RoundKeyOutput[107]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_108_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_15913, new_AGEMA_signal_15909, new_AGEMA_signal_15905, new_AGEMA_signal_15901}), .a ({new_AGEMA_signal_6144, new_AGEMA_signal_6143, new_AGEMA_signal_6142, KeyExpansionOutput[108]}), .c ({new_AGEMA_signal_6450, new_AGEMA_signal_6449, new_AGEMA_signal_6448, RoundKeyOutput[108]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_109_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_15897, new_AGEMA_signal_15893, new_AGEMA_signal_15889, new_AGEMA_signal_15885}), .a ({new_AGEMA_signal_6141, new_AGEMA_signal_6140, new_AGEMA_signal_6139, KeyExpansionOutput[109]}), .c ({new_AGEMA_signal_6453, new_AGEMA_signal_6452, new_AGEMA_signal_6451, RoundKeyOutput[109]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_110_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_15833, new_AGEMA_signal_15829, new_AGEMA_signal_15825, new_AGEMA_signal_15821}), .a ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, new_AGEMA_signal_6136, KeyExpansionOutput[110]}), .c ({new_AGEMA_signal_6456, new_AGEMA_signal_6455, new_AGEMA_signal_6454, RoundKeyOutput[110]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_111_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_15817, new_AGEMA_signal_15813, new_AGEMA_signal_15809, new_AGEMA_signal_15805}), .a ({new_AGEMA_signal_6135, new_AGEMA_signal_6134, new_AGEMA_signal_6133, KeyExpansionOutput[111]}), .c ({new_AGEMA_signal_6459, new_AGEMA_signal_6458, new_AGEMA_signal_6457, RoundKeyOutput[111]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_112_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_15801, new_AGEMA_signal_15797, new_AGEMA_signal_15793, new_AGEMA_signal_15789}), .a ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, new_AGEMA_signal_5986, KeyExpansionOutput[112]}), .c ({new_AGEMA_signal_6198, new_AGEMA_signal_6197, new_AGEMA_signal_6196, RoundKeyOutput[112]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_113_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_15785, new_AGEMA_signal_15781, new_AGEMA_signal_15777, new_AGEMA_signal_15773}), .a ({new_AGEMA_signal_6132, new_AGEMA_signal_6131, new_AGEMA_signal_6130, KeyExpansionOutput[113]}), .c ({new_AGEMA_signal_6462, new_AGEMA_signal_6461, new_AGEMA_signal_6460, RoundKeyOutput[113]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_114_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_15769, new_AGEMA_signal_15765, new_AGEMA_signal_15761, new_AGEMA_signal_15757}), .a ({new_AGEMA_signal_6129, new_AGEMA_signal_6128, new_AGEMA_signal_6127, KeyExpansionOutput[114]}), .c ({new_AGEMA_signal_6465, new_AGEMA_signal_6464, new_AGEMA_signal_6463, RoundKeyOutput[114]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_115_U1 ( .s (new_AGEMA_signal_16141), .b ({new_AGEMA_signal_15753, new_AGEMA_signal_15749, new_AGEMA_signal_15745, new_AGEMA_signal_15741}), .a ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, new_AGEMA_signal_6124, KeyExpansionOutput[115]}), .c ({new_AGEMA_signal_6468, new_AGEMA_signal_6467, new_AGEMA_signal_6466, RoundKeyOutput[115]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_116_U1 ( .s (new_AGEMA_signal_16165), .b ({new_AGEMA_signal_15737, new_AGEMA_signal_15733, new_AGEMA_signal_15729, new_AGEMA_signal_15725}), .a ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, new_AGEMA_signal_6121, KeyExpansionOutput[116]}), .c ({new_AGEMA_signal_6471, new_AGEMA_signal_6470, new_AGEMA_signal_6469, RoundKeyOutput[116]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_117_U1 ( .s (new_AGEMA_signal_16165), .b ({new_AGEMA_signal_15721, new_AGEMA_signal_15717, new_AGEMA_signal_15713, new_AGEMA_signal_15709}), .a ({new_AGEMA_signal_6120, new_AGEMA_signal_6119, new_AGEMA_signal_6118, KeyExpansionOutput[117]}), .c ({new_AGEMA_signal_6474, new_AGEMA_signal_6473, new_AGEMA_signal_6472, RoundKeyOutput[117]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_118_U1 ( .s (new_AGEMA_signal_16165), .b ({new_AGEMA_signal_15705, new_AGEMA_signal_15701, new_AGEMA_signal_15697, new_AGEMA_signal_15693}), .a ({new_AGEMA_signal_6117, new_AGEMA_signal_6116, new_AGEMA_signal_6115, KeyExpansionOutput[118]}), .c ({new_AGEMA_signal_6477, new_AGEMA_signal_6476, new_AGEMA_signal_6475, RoundKeyOutput[118]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_119_U1 ( .s (new_AGEMA_signal_16165), .b ({new_AGEMA_signal_15689, new_AGEMA_signal_15685, new_AGEMA_signal_15681, new_AGEMA_signal_15677}), .a ({new_AGEMA_signal_6114, new_AGEMA_signal_6113, new_AGEMA_signal_6112, KeyExpansionOutput[119]}), .c ({new_AGEMA_signal_6480, new_AGEMA_signal_6479, new_AGEMA_signal_6478, RoundKeyOutput[119]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_120_U1 ( .s (new_AGEMA_signal_16165), .b ({new_AGEMA_signal_15625, new_AGEMA_signal_15621, new_AGEMA_signal_15617, new_AGEMA_signal_15613}), .a ({new_AGEMA_signal_6111, new_AGEMA_signal_6110, new_AGEMA_signal_6109, KeyExpansionOutput[120]}), .c ({new_AGEMA_signal_6483, new_AGEMA_signal_6482, new_AGEMA_signal_6481, RoundKeyOutput[120]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_121_U1 ( .s (new_AGEMA_signal_16165), .b ({new_AGEMA_signal_15609, new_AGEMA_signal_15605, new_AGEMA_signal_15601, new_AGEMA_signal_15597}), .a ({new_AGEMA_signal_6399, new_AGEMA_signal_6398, new_AGEMA_signal_6397, KeyExpansionOutput[121]}), .c ({new_AGEMA_signal_6903, new_AGEMA_signal_6902, new_AGEMA_signal_6901, RoundKeyOutput[121]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_122_U1 ( .s (new_AGEMA_signal_16165), .b ({new_AGEMA_signal_15593, new_AGEMA_signal_15589, new_AGEMA_signal_15585, new_AGEMA_signal_15581}), .a ({new_AGEMA_signal_6396, new_AGEMA_signal_6395, new_AGEMA_signal_6394, KeyExpansionOutput[122]}), .c ({new_AGEMA_signal_6906, new_AGEMA_signal_6905, new_AGEMA_signal_6904, RoundKeyOutput[122]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_123_U1 ( .s (new_AGEMA_signal_16165), .b ({new_AGEMA_signal_15577, new_AGEMA_signal_15573, new_AGEMA_signal_15569, new_AGEMA_signal_15565}), .a ({new_AGEMA_signal_6393, new_AGEMA_signal_6392, new_AGEMA_signal_6391, KeyExpansionOutput[123]}), .c ({new_AGEMA_signal_6909, new_AGEMA_signal_6908, new_AGEMA_signal_6907, RoundKeyOutput[123]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_124_U1 ( .s (new_AGEMA_signal_16165), .b ({new_AGEMA_signal_15561, new_AGEMA_signal_15557, new_AGEMA_signal_15553, new_AGEMA_signal_15549}), .a ({new_AGEMA_signal_6390, new_AGEMA_signal_6389, new_AGEMA_signal_6388, KeyExpansionOutput[124]}), .c ({new_AGEMA_signal_6912, new_AGEMA_signal_6911, new_AGEMA_signal_6910, RoundKeyOutput[124]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_125_U1 ( .s (new_AGEMA_signal_16165), .b ({new_AGEMA_signal_15545, new_AGEMA_signal_15541, new_AGEMA_signal_15537, new_AGEMA_signal_15533}), .a ({new_AGEMA_signal_6387, new_AGEMA_signal_6386, new_AGEMA_signal_6385, KeyExpansionOutput[125]}), .c ({new_AGEMA_signal_6915, new_AGEMA_signal_6914, new_AGEMA_signal_6913, RoundKeyOutput[125]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_126_U1 ( .s (new_AGEMA_signal_16165), .b ({new_AGEMA_signal_15529, new_AGEMA_signal_15525, new_AGEMA_signal_15521, new_AGEMA_signal_15517}), .a ({new_AGEMA_signal_6384, new_AGEMA_signal_6383, new_AGEMA_signal_6382, KeyExpansionOutput[126]}), .c ({new_AGEMA_signal_6918, new_AGEMA_signal_6917, new_AGEMA_signal_6916, RoundKeyOutput[126]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(1)) MuxKeyExpansion_mux_inst_127_U1 ( .s (new_AGEMA_signal_16165), .b ({new_AGEMA_signal_15513, new_AGEMA_signal_15509, new_AGEMA_signal_15505, new_AGEMA_signal_15501}), .a ({new_AGEMA_signal_6381, new_AGEMA_signal_6380, new_AGEMA_signal_6379, KeyExpansionOutput[127]}), .c ({new_AGEMA_signal_6921, new_AGEMA_signal_6920, new_AGEMA_signal_6919, RoundKeyOutput[127]}) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C (clk), .D (new_AGEMA_signal_10080), .Q (new_AGEMA_signal_10081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2260 ( .C (clk), .D (new_AGEMA_signal_10084), .Q (new_AGEMA_signal_10085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2264 ( .C (clk), .D (new_AGEMA_signal_10088), .Q (new_AGEMA_signal_10089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2268 ( .C (clk), .D (new_AGEMA_signal_10092), .Q (new_AGEMA_signal_10093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2272 ( .C (clk), .D (new_AGEMA_signal_10096), .Q (new_AGEMA_signal_10097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2276 ( .C (clk), .D (new_AGEMA_signal_10100), .Q (new_AGEMA_signal_10101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2280 ( .C (clk), .D (new_AGEMA_signal_10104), .Q (new_AGEMA_signal_10105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2284 ( .C (clk), .D (new_AGEMA_signal_10108), .Q (new_AGEMA_signal_10109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2288 ( .C (clk), .D (new_AGEMA_signal_10112), .Q (new_AGEMA_signal_10113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2292 ( .C (clk), .D (new_AGEMA_signal_10116), .Q (new_AGEMA_signal_10117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2296 ( .C (clk), .D (new_AGEMA_signal_10120), .Q (new_AGEMA_signal_10121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2300 ( .C (clk), .D (new_AGEMA_signal_10124), .Q (new_AGEMA_signal_10125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2304 ( .C (clk), .D (new_AGEMA_signal_10128), .Q (new_AGEMA_signal_10129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2308 ( .C (clk), .D (new_AGEMA_signal_10132), .Q (new_AGEMA_signal_10133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2312 ( .C (clk), .D (new_AGEMA_signal_10136), .Q (new_AGEMA_signal_10137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2316 ( .C (clk), .D (new_AGEMA_signal_10140), .Q (new_AGEMA_signal_10141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2320 ( .C (clk), .D (new_AGEMA_signal_10144), .Q (new_AGEMA_signal_10145) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2324 ( .C (clk), .D (new_AGEMA_signal_10148), .Q (new_AGEMA_signal_10149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2328 ( .C (clk), .D (new_AGEMA_signal_10152), .Q (new_AGEMA_signal_10153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2332 ( .C (clk), .D (new_AGEMA_signal_10156), .Q (new_AGEMA_signal_10157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2336 ( .C (clk), .D (new_AGEMA_signal_10160), .Q (new_AGEMA_signal_10161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2340 ( .C (clk), .D (new_AGEMA_signal_10164), .Q (new_AGEMA_signal_10165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2344 ( .C (clk), .D (new_AGEMA_signal_10168), .Q (new_AGEMA_signal_10169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2348 ( .C (clk), .D (new_AGEMA_signal_10172), .Q (new_AGEMA_signal_10173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2352 ( .C (clk), .D (new_AGEMA_signal_10176), .Q (new_AGEMA_signal_10177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2356 ( .C (clk), .D (new_AGEMA_signal_10180), .Q (new_AGEMA_signal_10181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2360 ( .C (clk), .D (new_AGEMA_signal_10184), .Q (new_AGEMA_signal_10185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2364 ( .C (clk), .D (new_AGEMA_signal_10188), .Q (new_AGEMA_signal_10189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2368 ( .C (clk), .D (new_AGEMA_signal_10192), .Q (new_AGEMA_signal_10193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2372 ( .C (clk), .D (new_AGEMA_signal_10196), .Q (new_AGEMA_signal_10197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2376 ( .C (clk), .D (new_AGEMA_signal_10200), .Q (new_AGEMA_signal_10201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2380 ( .C (clk), .D (new_AGEMA_signal_10204), .Q (new_AGEMA_signal_10205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2384 ( .C (clk), .D (new_AGEMA_signal_10208), .Q (new_AGEMA_signal_10209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2388 ( .C (clk), .D (new_AGEMA_signal_10212), .Q (new_AGEMA_signal_10213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2392 ( .C (clk), .D (new_AGEMA_signal_10216), .Q (new_AGEMA_signal_10217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2396 ( .C (clk), .D (new_AGEMA_signal_10220), .Q (new_AGEMA_signal_10221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2400 ( .C (clk), .D (new_AGEMA_signal_10224), .Q (new_AGEMA_signal_10225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2404 ( .C (clk), .D (new_AGEMA_signal_10228), .Q (new_AGEMA_signal_10229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2408 ( .C (clk), .D (new_AGEMA_signal_10232), .Q (new_AGEMA_signal_10233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2412 ( .C (clk), .D (new_AGEMA_signal_10236), .Q (new_AGEMA_signal_10237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2416 ( .C (clk), .D (new_AGEMA_signal_10240), .Q (new_AGEMA_signal_10241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2420 ( .C (clk), .D (new_AGEMA_signal_10244), .Q (new_AGEMA_signal_10245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2424 ( .C (clk), .D (new_AGEMA_signal_10248), .Q (new_AGEMA_signal_10249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2428 ( .C (clk), .D (new_AGEMA_signal_10252), .Q (new_AGEMA_signal_10253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2432 ( .C (clk), .D (new_AGEMA_signal_10256), .Q (new_AGEMA_signal_10257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2436 ( .C (clk), .D (new_AGEMA_signal_10260), .Q (new_AGEMA_signal_10261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2440 ( .C (clk), .D (new_AGEMA_signal_10264), .Q (new_AGEMA_signal_10265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2444 ( .C (clk), .D (new_AGEMA_signal_10268), .Q (new_AGEMA_signal_10269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2448 ( .C (clk), .D (new_AGEMA_signal_10272), .Q (new_AGEMA_signal_10273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2452 ( .C (clk), .D (new_AGEMA_signal_10276), .Q (new_AGEMA_signal_10277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2456 ( .C (clk), .D (new_AGEMA_signal_10280), .Q (new_AGEMA_signal_10281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2460 ( .C (clk), .D (new_AGEMA_signal_10284), .Q (new_AGEMA_signal_10285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2464 ( .C (clk), .D (new_AGEMA_signal_10288), .Q (new_AGEMA_signal_10289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2468 ( .C (clk), .D (new_AGEMA_signal_10292), .Q (new_AGEMA_signal_10293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2472 ( .C (clk), .D (new_AGEMA_signal_10296), .Q (new_AGEMA_signal_10297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2476 ( .C (clk), .D (new_AGEMA_signal_10300), .Q (new_AGEMA_signal_10301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2480 ( .C (clk), .D (new_AGEMA_signal_10304), .Q (new_AGEMA_signal_10305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2484 ( .C (clk), .D (new_AGEMA_signal_10308), .Q (new_AGEMA_signal_10309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2488 ( .C (clk), .D (new_AGEMA_signal_10312), .Q (new_AGEMA_signal_10313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2492 ( .C (clk), .D (new_AGEMA_signal_10316), .Q (new_AGEMA_signal_10317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2496 ( .C (clk), .D (new_AGEMA_signal_10320), .Q (new_AGEMA_signal_10321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2500 ( .C (clk), .D (new_AGEMA_signal_10324), .Q (new_AGEMA_signal_10325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2504 ( .C (clk), .D (new_AGEMA_signal_10328), .Q (new_AGEMA_signal_10329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2508 ( .C (clk), .D (new_AGEMA_signal_10332), .Q (new_AGEMA_signal_10333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2512 ( .C (clk), .D (new_AGEMA_signal_10336), .Q (new_AGEMA_signal_10337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2516 ( .C (clk), .D (new_AGEMA_signal_10340), .Q (new_AGEMA_signal_10341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2520 ( .C (clk), .D (new_AGEMA_signal_10344), .Q (new_AGEMA_signal_10345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2524 ( .C (clk), .D (new_AGEMA_signal_10348), .Q (new_AGEMA_signal_10349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2528 ( .C (clk), .D (new_AGEMA_signal_10352), .Q (new_AGEMA_signal_10353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2532 ( .C (clk), .D (new_AGEMA_signal_10356), .Q (new_AGEMA_signal_10357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2536 ( .C (clk), .D (new_AGEMA_signal_10360), .Q (new_AGEMA_signal_10361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2540 ( .C (clk), .D (new_AGEMA_signal_10364), .Q (new_AGEMA_signal_10365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2544 ( .C (clk), .D (new_AGEMA_signal_10368), .Q (new_AGEMA_signal_10369) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2548 ( .C (clk), .D (new_AGEMA_signal_10372), .Q (new_AGEMA_signal_10373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2552 ( .C (clk), .D (new_AGEMA_signal_10376), .Q (new_AGEMA_signal_10377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2556 ( .C (clk), .D (new_AGEMA_signal_10380), .Q (new_AGEMA_signal_10381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2560 ( .C (clk), .D (new_AGEMA_signal_10384), .Q (new_AGEMA_signal_10385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2564 ( .C (clk), .D (new_AGEMA_signal_10388), .Q (new_AGEMA_signal_10389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2568 ( .C (clk), .D (new_AGEMA_signal_10392), .Q (new_AGEMA_signal_10393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2572 ( .C (clk), .D (new_AGEMA_signal_10396), .Q (new_AGEMA_signal_10397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2576 ( .C (clk), .D (new_AGEMA_signal_10400), .Q (new_AGEMA_signal_10401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2580 ( .C (clk), .D (new_AGEMA_signal_10404), .Q (new_AGEMA_signal_10405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2584 ( .C (clk), .D (new_AGEMA_signal_10408), .Q (new_AGEMA_signal_10409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2588 ( .C (clk), .D (new_AGEMA_signal_10412), .Q (new_AGEMA_signal_10413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2592 ( .C (clk), .D (new_AGEMA_signal_10416), .Q (new_AGEMA_signal_10417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2596 ( .C (clk), .D (new_AGEMA_signal_10420), .Q (new_AGEMA_signal_10421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2600 ( .C (clk), .D (new_AGEMA_signal_10424), .Q (new_AGEMA_signal_10425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2604 ( .C (clk), .D (new_AGEMA_signal_10428), .Q (new_AGEMA_signal_10429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2608 ( .C (clk), .D (new_AGEMA_signal_10432), .Q (new_AGEMA_signal_10433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2612 ( .C (clk), .D (new_AGEMA_signal_10436), .Q (new_AGEMA_signal_10437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2616 ( .C (clk), .D (new_AGEMA_signal_10440), .Q (new_AGEMA_signal_10441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2620 ( .C (clk), .D (new_AGEMA_signal_10444), .Q (new_AGEMA_signal_10445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2624 ( .C (clk), .D (new_AGEMA_signal_10448), .Q (new_AGEMA_signal_10449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2628 ( .C (clk), .D (new_AGEMA_signal_10452), .Q (new_AGEMA_signal_10453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2632 ( .C (clk), .D (new_AGEMA_signal_10456), .Q (new_AGEMA_signal_10457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2636 ( .C (clk), .D (new_AGEMA_signal_10460), .Q (new_AGEMA_signal_10461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2640 ( .C (clk), .D (new_AGEMA_signal_10464), .Q (new_AGEMA_signal_10465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2644 ( .C (clk), .D (new_AGEMA_signal_10468), .Q (new_AGEMA_signal_10469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2648 ( .C (clk), .D (new_AGEMA_signal_10472), .Q (new_AGEMA_signal_10473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2652 ( .C (clk), .D (new_AGEMA_signal_10476), .Q (new_AGEMA_signal_10477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2656 ( .C (clk), .D (new_AGEMA_signal_10480), .Q (new_AGEMA_signal_10481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2660 ( .C (clk), .D (new_AGEMA_signal_10484), .Q (new_AGEMA_signal_10485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2664 ( .C (clk), .D (new_AGEMA_signal_10488), .Q (new_AGEMA_signal_10489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2668 ( .C (clk), .D (new_AGEMA_signal_10492), .Q (new_AGEMA_signal_10493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2672 ( .C (clk), .D (new_AGEMA_signal_10496), .Q (new_AGEMA_signal_10497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2676 ( .C (clk), .D (new_AGEMA_signal_10500), .Q (new_AGEMA_signal_10501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2680 ( .C (clk), .D (new_AGEMA_signal_10504), .Q (new_AGEMA_signal_10505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2684 ( .C (clk), .D (new_AGEMA_signal_10508), .Q (new_AGEMA_signal_10509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2688 ( .C (clk), .D (new_AGEMA_signal_10512), .Q (new_AGEMA_signal_10513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2692 ( .C (clk), .D (new_AGEMA_signal_10516), .Q (new_AGEMA_signal_10517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2696 ( .C (clk), .D (new_AGEMA_signal_10520), .Q (new_AGEMA_signal_10521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2700 ( .C (clk), .D (new_AGEMA_signal_10524), .Q (new_AGEMA_signal_10525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2704 ( .C (clk), .D (new_AGEMA_signal_10528), .Q (new_AGEMA_signal_10529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2708 ( .C (clk), .D (new_AGEMA_signal_10532), .Q (new_AGEMA_signal_10533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2712 ( .C (clk), .D (new_AGEMA_signal_10536), .Q (new_AGEMA_signal_10537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2716 ( .C (clk), .D (new_AGEMA_signal_10540), .Q (new_AGEMA_signal_10541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2720 ( .C (clk), .D (new_AGEMA_signal_10544), .Q (new_AGEMA_signal_10545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2724 ( .C (clk), .D (new_AGEMA_signal_10548), .Q (new_AGEMA_signal_10549) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2728 ( .C (clk), .D (new_AGEMA_signal_10552), .Q (new_AGEMA_signal_10553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2732 ( .C (clk), .D (new_AGEMA_signal_10556), .Q (new_AGEMA_signal_10557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2736 ( .C (clk), .D (new_AGEMA_signal_10560), .Q (new_AGEMA_signal_10561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2740 ( .C (clk), .D (new_AGEMA_signal_10564), .Q (new_AGEMA_signal_10565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2744 ( .C (clk), .D (new_AGEMA_signal_10568), .Q (new_AGEMA_signal_10569) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2748 ( .C (clk), .D (new_AGEMA_signal_10572), .Q (new_AGEMA_signal_10573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2752 ( .C (clk), .D (new_AGEMA_signal_10576), .Q (new_AGEMA_signal_10577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2756 ( .C (clk), .D (new_AGEMA_signal_10580), .Q (new_AGEMA_signal_10581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2760 ( .C (clk), .D (new_AGEMA_signal_10584), .Q (new_AGEMA_signal_10585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2764 ( .C (clk), .D (new_AGEMA_signal_10588), .Q (new_AGEMA_signal_10589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2768 ( .C (clk), .D (new_AGEMA_signal_10592), .Q (new_AGEMA_signal_10593) ) ;
    buf_clk new_AGEMA_reg_buffer_3636 ( .C (clk), .D (new_AGEMA_signal_11460), .Q (new_AGEMA_signal_11461) ) ;
    buf_clk new_AGEMA_reg_buffer_3640 ( .C (clk), .D (new_AGEMA_signal_11464), .Q (new_AGEMA_signal_11465) ) ;
    buf_clk new_AGEMA_reg_buffer_3644 ( .C (clk), .D (new_AGEMA_signal_11468), .Q (new_AGEMA_signal_11469) ) ;
    buf_clk new_AGEMA_reg_buffer_3648 ( .C (clk), .D (new_AGEMA_signal_11472), .Q (new_AGEMA_signal_11473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3652 ( .C (clk), .D (new_AGEMA_signal_11476), .Q (new_AGEMA_signal_11477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3656 ( .C (clk), .D (new_AGEMA_signal_11480), .Q (new_AGEMA_signal_11481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3660 ( .C (clk), .D (new_AGEMA_signal_11484), .Q (new_AGEMA_signal_11485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3664 ( .C (clk), .D (new_AGEMA_signal_11488), .Q (new_AGEMA_signal_11489) ) ;
    buf_clk new_AGEMA_reg_buffer_3668 ( .C (clk), .D (new_AGEMA_signal_11492), .Q (new_AGEMA_signal_11493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3672 ( .C (clk), .D (new_AGEMA_signal_11496), .Q (new_AGEMA_signal_11497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3676 ( .C (clk), .D (new_AGEMA_signal_11500), .Q (new_AGEMA_signal_11501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3680 ( .C (clk), .D (new_AGEMA_signal_11504), .Q (new_AGEMA_signal_11505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3684 ( .C (clk), .D (new_AGEMA_signal_11508), .Q (new_AGEMA_signal_11509) ) ;
    buf_clk new_AGEMA_reg_buffer_3688 ( .C (clk), .D (new_AGEMA_signal_11512), .Q (new_AGEMA_signal_11513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3692 ( .C (clk), .D (new_AGEMA_signal_11516), .Q (new_AGEMA_signal_11517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3696 ( .C (clk), .D (new_AGEMA_signal_11520), .Q (new_AGEMA_signal_11521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3700 ( .C (clk), .D (new_AGEMA_signal_11524), .Q (new_AGEMA_signal_11525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3704 ( .C (clk), .D (new_AGEMA_signal_11528), .Q (new_AGEMA_signal_11529) ) ;
    buf_clk new_AGEMA_reg_buffer_3708 ( .C (clk), .D (new_AGEMA_signal_11532), .Q (new_AGEMA_signal_11533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3712 ( .C (clk), .D (new_AGEMA_signal_11536), .Q (new_AGEMA_signal_11537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3716 ( .C (clk), .D (new_AGEMA_signal_11540), .Q (new_AGEMA_signal_11541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3720 ( .C (clk), .D (new_AGEMA_signal_11544), .Q (new_AGEMA_signal_11545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3724 ( .C (clk), .D (new_AGEMA_signal_11548), .Q (new_AGEMA_signal_11549) ) ;
    buf_clk new_AGEMA_reg_buffer_3728 ( .C (clk), .D (new_AGEMA_signal_11552), .Q (new_AGEMA_signal_11553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3732 ( .C (clk), .D (new_AGEMA_signal_11556), .Q (new_AGEMA_signal_11557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3736 ( .C (clk), .D (new_AGEMA_signal_11560), .Q (new_AGEMA_signal_11561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3740 ( .C (clk), .D (new_AGEMA_signal_11564), .Q (new_AGEMA_signal_11565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3744 ( .C (clk), .D (new_AGEMA_signal_11568), .Q (new_AGEMA_signal_11569) ) ;
    buf_clk new_AGEMA_reg_buffer_3748 ( .C (clk), .D (new_AGEMA_signal_11572), .Q (new_AGEMA_signal_11573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3752 ( .C (clk), .D (new_AGEMA_signal_11576), .Q (new_AGEMA_signal_11577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3756 ( .C (clk), .D (new_AGEMA_signal_11580), .Q (new_AGEMA_signal_11581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3760 ( .C (clk), .D (new_AGEMA_signal_11584), .Q (new_AGEMA_signal_11585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3764 ( .C (clk), .D (new_AGEMA_signal_11588), .Q (new_AGEMA_signal_11589) ) ;
    buf_clk new_AGEMA_reg_buffer_3768 ( .C (clk), .D (new_AGEMA_signal_11592), .Q (new_AGEMA_signal_11593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3772 ( .C (clk), .D (new_AGEMA_signal_11596), .Q (new_AGEMA_signal_11597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3776 ( .C (clk), .D (new_AGEMA_signal_11600), .Q (new_AGEMA_signal_11601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3780 ( .C (clk), .D (new_AGEMA_signal_11604), .Q (new_AGEMA_signal_11605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3784 ( .C (clk), .D (new_AGEMA_signal_11608), .Q (new_AGEMA_signal_11609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3788 ( .C (clk), .D (new_AGEMA_signal_11612), .Q (new_AGEMA_signal_11613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3792 ( .C (clk), .D (new_AGEMA_signal_11616), .Q (new_AGEMA_signal_11617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3796 ( .C (clk), .D (new_AGEMA_signal_11620), .Q (new_AGEMA_signal_11621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3800 ( .C (clk), .D (new_AGEMA_signal_11624), .Q (new_AGEMA_signal_11625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3804 ( .C (clk), .D (new_AGEMA_signal_11628), .Q (new_AGEMA_signal_11629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3808 ( .C (clk), .D (new_AGEMA_signal_11632), .Q (new_AGEMA_signal_11633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3812 ( .C (clk), .D (new_AGEMA_signal_11636), .Q (new_AGEMA_signal_11637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3816 ( .C (clk), .D (new_AGEMA_signal_11640), .Q (new_AGEMA_signal_11641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3820 ( .C (clk), .D (new_AGEMA_signal_11644), .Q (new_AGEMA_signal_11645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3824 ( .C (clk), .D (new_AGEMA_signal_11648), .Q (new_AGEMA_signal_11649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3828 ( .C (clk), .D (new_AGEMA_signal_11652), .Q (new_AGEMA_signal_11653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3832 ( .C (clk), .D (new_AGEMA_signal_11656), .Q (new_AGEMA_signal_11657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3836 ( .C (clk), .D (new_AGEMA_signal_11660), .Q (new_AGEMA_signal_11661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3840 ( .C (clk), .D (new_AGEMA_signal_11664), .Q (new_AGEMA_signal_11665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3844 ( .C (clk), .D (new_AGEMA_signal_11668), .Q (new_AGEMA_signal_11669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3848 ( .C (clk), .D (new_AGEMA_signal_11672), .Q (new_AGEMA_signal_11673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3852 ( .C (clk), .D (new_AGEMA_signal_11676), .Q (new_AGEMA_signal_11677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3856 ( .C (clk), .D (new_AGEMA_signal_11680), .Q (new_AGEMA_signal_11681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3860 ( .C (clk), .D (new_AGEMA_signal_11684), .Q (new_AGEMA_signal_11685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3864 ( .C (clk), .D (new_AGEMA_signal_11688), .Q (new_AGEMA_signal_11689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3868 ( .C (clk), .D (new_AGEMA_signal_11692), .Q (new_AGEMA_signal_11693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3872 ( .C (clk), .D (new_AGEMA_signal_11696), .Q (new_AGEMA_signal_11697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3876 ( .C (clk), .D (new_AGEMA_signal_11700), .Q (new_AGEMA_signal_11701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3880 ( .C (clk), .D (new_AGEMA_signal_11704), .Q (new_AGEMA_signal_11705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3884 ( .C (clk), .D (new_AGEMA_signal_11708), .Q (new_AGEMA_signal_11709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3888 ( .C (clk), .D (new_AGEMA_signal_11712), .Q (new_AGEMA_signal_11713) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3892 ( .C (clk), .D (new_AGEMA_signal_11716), .Q (new_AGEMA_signal_11717) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3896 ( .C (clk), .D (new_AGEMA_signal_11720), .Q (new_AGEMA_signal_11721) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3900 ( .C (clk), .D (new_AGEMA_signal_11724), .Q (new_AGEMA_signal_11725) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3904 ( .C (clk), .D (new_AGEMA_signal_11728), .Q (new_AGEMA_signal_11729) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3908 ( .C (clk), .D (new_AGEMA_signal_11732), .Q (new_AGEMA_signal_11733) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3912 ( .C (clk), .D (new_AGEMA_signal_11736), .Q (new_AGEMA_signal_11737) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3916 ( .C (clk), .D (new_AGEMA_signal_11740), .Q (new_AGEMA_signal_11741) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3920 ( .C (clk), .D (new_AGEMA_signal_11744), .Q (new_AGEMA_signal_11745) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3924 ( .C (clk), .D (new_AGEMA_signal_11748), .Q (new_AGEMA_signal_11749) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3928 ( .C (clk), .D (new_AGEMA_signal_11752), .Q (new_AGEMA_signal_11753) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3932 ( .C (clk), .D (new_AGEMA_signal_11756), .Q (new_AGEMA_signal_11757) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3936 ( .C (clk), .D (new_AGEMA_signal_11760), .Q (new_AGEMA_signal_11761) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3940 ( .C (clk), .D (new_AGEMA_signal_11764), .Q (new_AGEMA_signal_11765) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3944 ( .C (clk), .D (new_AGEMA_signal_11768), .Q (new_AGEMA_signal_11769) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3948 ( .C (clk), .D (new_AGEMA_signal_11772), .Q (new_AGEMA_signal_11773) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3952 ( .C (clk), .D (new_AGEMA_signal_11776), .Q (new_AGEMA_signal_11777) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3956 ( .C (clk), .D (new_AGEMA_signal_11780), .Q (new_AGEMA_signal_11781) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3960 ( .C (clk), .D (new_AGEMA_signal_11784), .Q (new_AGEMA_signal_11785) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3964 ( .C (clk), .D (new_AGEMA_signal_11788), .Q (new_AGEMA_signal_11789) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3968 ( .C (clk), .D (new_AGEMA_signal_11792), .Q (new_AGEMA_signal_11793) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3972 ( .C (clk), .D (new_AGEMA_signal_11796), .Q (new_AGEMA_signal_11797) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3976 ( .C (clk), .D (new_AGEMA_signal_11800), .Q (new_AGEMA_signal_11801) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3980 ( .C (clk), .D (new_AGEMA_signal_11804), .Q (new_AGEMA_signal_11805) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3984 ( .C (clk), .D (new_AGEMA_signal_11808), .Q (new_AGEMA_signal_11809) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3988 ( .C (clk), .D (new_AGEMA_signal_11812), .Q (new_AGEMA_signal_11813) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3992 ( .C (clk), .D (new_AGEMA_signal_11816), .Q (new_AGEMA_signal_11817) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3996 ( .C (clk), .D (new_AGEMA_signal_11820), .Q (new_AGEMA_signal_11821) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4000 ( .C (clk), .D (new_AGEMA_signal_11824), .Q (new_AGEMA_signal_11825) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4004 ( .C (clk), .D (new_AGEMA_signal_11828), .Q (new_AGEMA_signal_11829) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4008 ( .C (clk), .D (new_AGEMA_signal_11832), .Q (new_AGEMA_signal_11833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4012 ( .C (clk), .D (new_AGEMA_signal_11836), .Q (new_AGEMA_signal_11837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4016 ( .C (clk), .D (new_AGEMA_signal_11840), .Q (new_AGEMA_signal_11841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4020 ( .C (clk), .D (new_AGEMA_signal_11844), .Q (new_AGEMA_signal_11845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4024 ( .C (clk), .D (new_AGEMA_signal_11848), .Q (new_AGEMA_signal_11849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4028 ( .C (clk), .D (new_AGEMA_signal_11852), .Q (new_AGEMA_signal_11853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4032 ( .C (clk), .D (new_AGEMA_signal_11856), .Q (new_AGEMA_signal_11857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4036 ( .C (clk), .D (new_AGEMA_signal_11860), .Q (new_AGEMA_signal_11861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4040 ( .C (clk), .D (new_AGEMA_signal_11864), .Q (new_AGEMA_signal_11865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4044 ( .C (clk), .D (new_AGEMA_signal_11868), .Q (new_AGEMA_signal_11869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4048 ( .C (clk), .D (new_AGEMA_signal_11872), .Q (new_AGEMA_signal_11873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4052 ( .C (clk), .D (new_AGEMA_signal_11876), .Q (new_AGEMA_signal_11877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4056 ( .C (clk), .D (new_AGEMA_signal_11880), .Q (new_AGEMA_signal_11881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4060 ( .C (clk), .D (new_AGEMA_signal_11884), .Q (new_AGEMA_signal_11885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4064 ( .C (clk), .D (new_AGEMA_signal_11888), .Q (new_AGEMA_signal_11889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4068 ( .C (clk), .D (new_AGEMA_signal_11892), .Q (new_AGEMA_signal_11893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4072 ( .C (clk), .D (new_AGEMA_signal_11896), .Q (new_AGEMA_signal_11897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4076 ( .C (clk), .D (new_AGEMA_signal_11900), .Q (new_AGEMA_signal_11901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4080 ( .C (clk), .D (new_AGEMA_signal_11904), .Q (new_AGEMA_signal_11905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4084 ( .C (clk), .D (new_AGEMA_signal_11908), .Q (new_AGEMA_signal_11909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4088 ( .C (clk), .D (new_AGEMA_signal_11912), .Q (new_AGEMA_signal_11913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4092 ( .C (clk), .D (new_AGEMA_signal_11916), .Q (new_AGEMA_signal_11917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4096 ( .C (clk), .D (new_AGEMA_signal_11920), .Q (new_AGEMA_signal_11921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4100 ( .C (clk), .D (new_AGEMA_signal_11924), .Q (new_AGEMA_signal_11925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4104 ( .C (clk), .D (new_AGEMA_signal_11928), .Q (new_AGEMA_signal_11929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4108 ( .C (clk), .D (new_AGEMA_signal_11932), .Q (new_AGEMA_signal_11933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4112 ( .C (clk), .D (new_AGEMA_signal_11936), .Q (new_AGEMA_signal_11937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4116 ( .C (clk), .D (new_AGEMA_signal_11940), .Q (new_AGEMA_signal_11941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4120 ( .C (clk), .D (new_AGEMA_signal_11944), .Q (new_AGEMA_signal_11945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4124 ( .C (clk), .D (new_AGEMA_signal_11948), .Q (new_AGEMA_signal_11949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4128 ( .C (clk), .D (new_AGEMA_signal_11952), .Q (new_AGEMA_signal_11953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4132 ( .C (clk), .D (new_AGEMA_signal_11956), .Q (new_AGEMA_signal_11957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4136 ( .C (clk), .D (new_AGEMA_signal_11960), .Q (new_AGEMA_signal_11961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4140 ( .C (clk), .D (new_AGEMA_signal_11964), .Q (new_AGEMA_signal_11965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4144 ( .C (clk), .D (new_AGEMA_signal_11968), .Q (new_AGEMA_signal_11969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4148 ( .C (clk), .D (new_AGEMA_signal_11972), .Q (new_AGEMA_signal_11973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4152 ( .C (clk), .D (new_AGEMA_signal_11976), .Q (new_AGEMA_signal_11977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4156 ( .C (clk), .D (new_AGEMA_signal_11980), .Q (new_AGEMA_signal_11981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4160 ( .C (clk), .D (new_AGEMA_signal_11984), .Q (new_AGEMA_signal_11985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4164 ( .C (clk), .D (new_AGEMA_signal_11988), .Q (new_AGEMA_signal_11989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4168 ( .C (clk), .D (new_AGEMA_signal_11992), .Q (new_AGEMA_signal_11993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4172 ( .C (clk), .D (new_AGEMA_signal_11996), .Q (new_AGEMA_signal_11997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4176 ( .C (clk), .D (new_AGEMA_signal_12000), .Q (new_AGEMA_signal_12001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4180 ( .C (clk), .D (new_AGEMA_signal_12004), .Q (new_AGEMA_signal_12005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4184 ( .C (clk), .D (new_AGEMA_signal_12008), .Q (new_AGEMA_signal_12009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4188 ( .C (clk), .D (new_AGEMA_signal_12012), .Q (new_AGEMA_signal_12013) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4192 ( .C (clk), .D (new_AGEMA_signal_12016), .Q (new_AGEMA_signal_12017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4196 ( .C (clk), .D (new_AGEMA_signal_12020), .Q (new_AGEMA_signal_12021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4200 ( .C (clk), .D (new_AGEMA_signal_12024), .Q (new_AGEMA_signal_12025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4204 ( .C (clk), .D (new_AGEMA_signal_12028), .Q (new_AGEMA_signal_12029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4208 ( .C (clk), .D (new_AGEMA_signal_12032), .Q (new_AGEMA_signal_12033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4212 ( .C (clk), .D (new_AGEMA_signal_12036), .Q (new_AGEMA_signal_12037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4216 ( .C (clk), .D (new_AGEMA_signal_12040), .Q (new_AGEMA_signal_12041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4220 ( .C (clk), .D (new_AGEMA_signal_12044), .Q (new_AGEMA_signal_12045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4224 ( .C (clk), .D (new_AGEMA_signal_12048), .Q (new_AGEMA_signal_12049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4228 ( .C (clk), .D (new_AGEMA_signal_12052), .Q (new_AGEMA_signal_12053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4232 ( .C (clk), .D (new_AGEMA_signal_12056), .Q (new_AGEMA_signal_12057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4236 ( .C (clk), .D (new_AGEMA_signal_12060), .Q (new_AGEMA_signal_12061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4240 ( .C (clk), .D (new_AGEMA_signal_12064), .Q (new_AGEMA_signal_12065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4244 ( .C (clk), .D (new_AGEMA_signal_12068), .Q (new_AGEMA_signal_12069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4248 ( .C (clk), .D (new_AGEMA_signal_12072), .Q (new_AGEMA_signal_12073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4252 ( .C (clk), .D (new_AGEMA_signal_12076), .Q (new_AGEMA_signal_12077) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4256 ( .C (clk), .D (new_AGEMA_signal_12080), .Q (new_AGEMA_signal_12081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4260 ( .C (clk), .D (new_AGEMA_signal_12084), .Q (new_AGEMA_signal_12085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4264 ( .C (clk), .D (new_AGEMA_signal_12088), .Q (new_AGEMA_signal_12089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4268 ( .C (clk), .D (new_AGEMA_signal_12092), .Q (new_AGEMA_signal_12093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4272 ( .C (clk), .D (new_AGEMA_signal_12096), .Q (new_AGEMA_signal_12097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4276 ( .C (clk), .D (new_AGEMA_signal_12100), .Q (new_AGEMA_signal_12101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4280 ( .C (clk), .D (new_AGEMA_signal_12104), .Q (new_AGEMA_signal_12105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4284 ( .C (clk), .D (new_AGEMA_signal_12108), .Q (new_AGEMA_signal_12109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4288 ( .C (clk), .D (new_AGEMA_signal_12112), .Q (new_AGEMA_signal_12113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4292 ( .C (clk), .D (new_AGEMA_signal_12116), .Q (new_AGEMA_signal_12117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4296 ( .C (clk), .D (new_AGEMA_signal_12120), .Q (new_AGEMA_signal_12121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4300 ( .C (clk), .D (new_AGEMA_signal_12124), .Q (new_AGEMA_signal_12125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4304 ( .C (clk), .D (new_AGEMA_signal_12128), .Q (new_AGEMA_signal_12129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4308 ( .C (clk), .D (new_AGEMA_signal_12132), .Q (new_AGEMA_signal_12133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4312 ( .C (clk), .D (new_AGEMA_signal_12136), .Q (new_AGEMA_signal_12137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4316 ( .C (clk), .D (new_AGEMA_signal_12140), .Q (new_AGEMA_signal_12141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4320 ( .C (clk), .D (new_AGEMA_signal_12144), .Q (new_AGEMA_signal_12145) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4324 ( .C (clk), .D (new_AGEMA_signal_12148), .Q (new_AGEMA_signal_12149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4328 ( .C (clk), .D (new_AGEMA_signal_12152), .Q (new_AGEMA_signal_12153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4332 ( .C (clk), .D (new_AGEMA_signal_12156), .Q (new_AGEMA_signal_12157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4336 ( .C (clk), .D (new_AGEMA_signal_12160), .Q (new_AGEMA_signal_12161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4340 ( .C (clk), .D (new_AGEMA_signal_12164), .Q (new_AGEMA_signal_12165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4344 ( .C (clk), .D (new_AGEMA_signal_12168), .Q (new_AGEMA_signal_12169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4348 ( .C (clk), .D (new_AGEMA_signal_12172), .Q (new_AGEMA_signal_12173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4352 ( .C (clk), .D (new_AGEMA_signal_12176), .Q (new_AGEMA_signal_12177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4356 ( .C (clk), .D (new_AGEMA_signal_12180), .Q (new_AGEMA_signal_12181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4360 ( .C (clk), .D (new_AGEMA_signal_12184), .Q (new_AGEMA_signal_12185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4364 ( .C (clk), .D (new_AGEMA_signal_12188), .Q (new_AGEMA_signal_12189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4368 ( .C (clk), .D (new_AGEMA_signal_12192), .Q (new_AGEMA_signal_12193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4372 ( .C (clk), .D (new_AGEMA_signal_12196), .Q (new_AGEMA_signal_12197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4376 ( .C (clk), .D (new_AGEMA_signal_12200), .Q (new_AGEMA_signal_12201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4380 ( .C (clk), .D (new_AGEMA_signal_12204), .Q (new_AGEMA_signal_12205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4384 ( .C (clk), .D (new_AGEMA_signal_12208), .Q (new_AGEMA_signal_12209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4388 ( .C (clk), .D (new_AGEMA_signal_12212), .Q (new_AGEMA_signal_12213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4392 ( .C (clk), .D (new_AGEMA_signal_12216), .Q (new_AGEMA_signal_12217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4396 ( .C (clk), .D (new_AGEMA_signal_12220), .Q (new_AGEMA_signal_12221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4400 ( .C (clk), .D (new_AGEMA_signal_12224), .Q (new_AGEMA_signal_12225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4404 ( .C (clk), .D (new_AGEMA_signal_12228), .Q (new_AGEMA_signal_12229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4408 ( .C (clk), .D (new_AGEMA_signal_12232), .Q (new_AGEMA_signal_12233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4412 ( .C (clk), .D (new_AGEMA_signal_12236), .Q (new_AGEMA_signal_12237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4416 ( .C (clk), .D (new_AGEMA_signal_12240), .Q (new_AGEMA_signal_12241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4420 ( .C (clk), .D (new_AGEMA_signal_12244), .Q (new_AGEMA_signal_12245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4424 ( .C (clk), .D (new_AGEMA_signal_12248), .Q (new_AGEMA_signal_12249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4428 ( .C (clk), .D (new_AGEMA_signal_12252), .Q (new_AGEMA_signal_12253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4432 ( .C (clk), .D (new_AGEMA_signal_12256), .Q (new_AGEMA_signal_12257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4436 ( .C (clk), .D (new_AGEMA_signal_12260), .Q (new_AGEMA_signal_12261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4440 ( .C (clk), .D (new_AGEMA_signal_12264), .Q (new_AGEMA_signal_12265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4444 ( .C (clk), .D (new_AGEMA_signal_12268), .Q (new_AGEMA_signal_12269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4448 ( .C (clk), .D (new_AGEMA_signal_12272), .Q (new_AGEMA_signal_12273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4452 ( .C (clk), .D (new_AGEMA_signal_12276), .Q (new_AGEMA_signal_12277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4456 ( .C (clk), .D (new_AGEMA_signal_12280), .Q (new_AGEMA_signal_12281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4460 ( .C (clk), .D (new_AGEMA_signal_12284), .Q (new_AGEMA_signal_12285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4464 ( .C (clk), .D (new_AGEMA_signal_12288), .Q (new_AGEMA_signal_12289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4468 ( .C (clk), .D (new_AGEMA_signal_12292), .Q (new_AGEMA_signal_12293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4472 ( .C (clk), .D (new_AGEMA_signal_12296), .Q (new_AGEMA_signal_12297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4476 ( .C (clk), .D (new_AGEMA_signal_12300), .Q (new_AGEMA_signal_12301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4480 ( .C (clk), .D (new_AGEMA_signal_12304), .Q (new_AGEMA_signal_12305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4484 ( .C (clk), .D (new_AGEMA_signal_12308), .Q (new_AGEMA_signal_12309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4488 ( .C (clk), .D (new_AGEMA_signal_12312), .Q (new_AGEMA_signal_12313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4492 ( .C (clk), .D (new_AGEMA_signal_12316), .Q (new_AGEMA_signal_12317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4496 ( .C (clk), .D (new_AGEMA_signal_12320), .Q (new_AGEMA_signal_12321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4500 ( .C (clk), .D (new_AGEMA_signal_12324), .Q (new_AGEMA_signal_12325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4504 ( .C (clk), .D (new_AGEMA_signal_12328), .Q (new_AGEMA_signal_12329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4508 ( .C (clk), .D (new_AGEMA_signal_12332), .Q (new_AGEMA_signal_12333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4512 ( .C (clk), .D (new_AGEMA_signal_12336), .Q (new_AGEMA_signal_12337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4516 ( .C (clk), .D (new_AGEMA_signal_12340), .Q (new_AGEMA_signal_12341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4520 ( .C (clk), .D (new_AGEMA_signal_12344), .Q (new_AGEMA_signal_12345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4524 ( .C (clk), .D (new_AGEMA_signal_12348), .Q (new_AGEMA_signal_12349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4528 ( .C (clk), .D (new_AGEMA_signal_12352), .Q (new_AGEMA_signal_12353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4532 ( .C (clk), .D (new_AGEMA_signal_12356), .Q (new_AGEMA_signal_12357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4536 ( .C (clk), .D (new_AGEMA_signal_12360), .Q (new_AGEMA_signal_12361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4540 ( .C (clk), .D (new_AGEMA_signal_12364), .Q (new_AGEMA_signal_12365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4544 ( .C (clk), .D (new_AGEMA_signal_12368), .Q (new_AGEMA_signal_12369) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4548 ( .C (clk), .D (new_AGEMA_signal_12372), .Q (new_AGEMA_signal_12373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4552 ( .C (clk), .D (new_AGEMA_signal_12376), .Q (new_AGEMA_signal_12377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4556 ( .C (clk), .D (new_AGEMA_signal_12380), .Q (new_AGEMA_signal_12381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4560 ( .C (clk), .D (new_AGEMA_signal_12384), .Q (new_AGEMA_signal_12385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4564 ( .C (clk), .D (new_AGEMA_signal_12388), .Q (new_AGEMA_signal_12389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4568 ( .C (clk), .D (new_AGEMA_signal_12392), .Q (new_AGEMA_signal_12393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4572 ( .C (clk), .D (new_AGEMA_signal_12396), .Q (new_AGEMA_signal_12397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4576 ( .C (clk), .D (new_AGEMA_signal_12400), .Q (new_AGEMA_signal_12401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4580 ( .C (clk), .D (new_AGEMA_signal_12404), .Q (new_AGEMA_signal_12405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4584 ( .C (clk), .D (new_AGEMA_signal_12408), .Q (new_AGEMA_signal_12409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4588 ( .C (clk), .D (new_AGEMA_signal_12412), .Q (new_AGEMA_signal_12413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4592 ( .C (clk), .D (new_AGEMA_signal_12416), .Q (new_AGEMA_signal_12417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4596 ( .C (clk), .D (new_AGEMA_signal_12420), .Q (new_AGEMA_signal_12421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4600 ( .C (clk), .D (new_AGEMA_signal_12424), .Q (new_AGEMA_signal_12425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4604 ( .C (clk), .D (new_AGEMA_signal_12428), .Q (new_AGEMA_signal_12429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4608 ( .C (clk), .D (new_AGEMA_signal_12432), .Q (new_AGEMA_signal_12433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4612 ( .C (clk), .D (new_AGEMA_signal_12436), .Q (new_AGEMA_signal_12437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4616 ( .C (clk), .D (new_AGEMA_signal_12440), .Q (new_AGEMA_signal_12441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4620 ( .C (clk), .D (new_AGEMA_signal_12444), .Q (new_AGEMA_signal_12445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4624 ( .C (clk), .D (new_AGEMA_signal_12448), .Q (new_AGEMA_signal_12449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4628 ( .C (clk), .D (new_AGEMA_signal_12452), .Q (new_AGEMA_signal_12453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4632 ( .C (clk), .D (new_AGEMA_signal_12456), .Q (new_AGEMA_signal_12457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4636 ( .C (clk), .D (new_AGEMA_signal_12460), .Q (new_AGEMA_signal_12461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4640 ( .C (clk), .D (new_AGEMA_signal_12464), .Q (new_AGEMA_signal_12465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4644 ( .C (clk), .D (new_AGEMA_signal_12468), .Q (new_AGEMA_signal_12469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4648 ( .C (clk), .D (new_AGEMA_signal_12472), .Q (new_AGEMA_signal_12473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4652 ( .C (clk), .D (new_AGEMA_signal_12476), .Q (new_AGEMA_signal_12477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4656 ( .C (clk), .D (new_AGEMA_signal_12480), .Q (new_AGEMA_signal_12481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4660 ( .C (clk), .D (new_AGEMA_signal_12484), .Q (new_AGEMA_signal_12485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4664 ( .C (clk), .D (new_AGEMA_signal_12488), .Q (new_AGEMA_signal_12489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4668 ( .C (clk), .D (new_AGEMA_signal_12492), .Q (new_AGEMA_signal_12493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4672 ( .C (clk), .D (new_AGEMA_signal_12496), .Q (new_AGEMA_signal_12497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4676 ( .C (clk), .D (new_AGEMA_signal_12500), .Q (new_AGEMA_signal_12501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4680 ( .C (clk), .D (new_AGEMA_signal_12504), .Q (new_AGEMA_signal_12505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4684 ( .C (clk), .D (new_AGEMA_signal_12508), .Q (new_AGEMA_signal_12509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4688 ( .C (clk), .D (new_AGEMA_signal_12512), .Q (new_AGEMA_signal_12513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4692 ( .C (clk), .D (new_AGEMA_signal_12516), .Q (new_AGEMA_signal_12517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4696 ( .C (clk), .D (new_AGEMA_signal_12520), .Q (new_AGEMA_signal_12521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4700 ( .C (clk), .D (new_AGEMA_signal_12524), .Q (new_AGEMA_signal_12525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4704 ( .C (clk), .D (new_AGEMA_signal_12528), .Q (new_AGEMA_signal_12529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4708 ( .C (clk), .D (new_AGEMA_signal_12532), .Q (new_AGEMA_signal_12533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4712 ( .C (clk), .D (new_AGEMA_signal_12536), .Q (new_AGEMA_signal_12537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4716 ( .C (clk), .D (new_AGEMA_signal_12540), .Q (new_AGEMA_signal_12541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4720 ( .C (clk), .D (new_AGEMA_signal_12544), .Q (new_AGEMA_signal_12545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4724 ( .C (clk), .D (new_AGEMA_signal_12548), .Q (new_AGEMA_signal_12549) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4728 ( .C (clk), .D (new_AGEMA_signal_12552), .Q (new_AGEMA_signal_12553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4732 ( .C (clk), .D (new_AGEMA_signal_12556), .Q (new_AGEMA_signal_12557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4736 ( .C (clk), .D (new_AGEMA_signal_12560), .Q (new_AGEMA_signal_12561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4740 ( .C (clk), .D (new_AGEMA_signal_12564), .Q (new_AGEMA_signal_12565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4744 ( .C (clk), .D (new_AGEMA_signal_12568), .Q (new_AGEMA_signal_12569) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4748 ( .C (clk), .D (new_AGEMA_signal_12572), .Q (new_AGEMA_signal_12573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4752 ( .C (clk), .D (new_AGEMA_signal_12576), .Q (new_AGEMA_signal_12577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4756 ( .C (clk), .D (new_AGEMA_signal_12580), .Q (new_AGEMA_signal_12581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4760 ( .C (clk), .D (new_AGEMA_signal_12584), .Q (new_AGEMA_signal_12585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4764 ( .C (clk), .D (new_AGEMA_signal_12588), .Q (new_AGEMA_signal_12589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4768 ( .C (clk), .D (new_AGEMA_signal_12592), .Q (new_AGEMA_signal_12593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4772 ( .C (clk), .D (new_AGEMA_signal_12596), .Q (new_AGEMA_signal_12597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4776 ( .C (clk), .D (new_AGEMA_signal_12600), .Q (new_AGEMA_signal_12601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4780 ( .C (clk), .D (new_AGEMA_signal_12604), .Q (new_AGEMA_signal_12605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4784 ( .C (clk), .D (new_AGEMA_signal_12608), .Q (new_AGEMA_signal_12609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4788 ( .C (clk), .D (new_AGEMA_signal_12612), .Q (new_AGEMA_signal_12613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4792 ( .C (clk), .D (new_AGEMA_signal_12616), .Q (new_AGEMA_signal_12617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4796 ( .C (clk), .D (new_AGEMA_signal_12620), .Q (new_AGEMA_signal_12621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4800 ( .C (clk), .D (new_AGEMA_signal_12624), .Q (new_AGEMA_signal_12625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4804 ( .C (clk), .D (new_AGEMA_signal_12628), .Q (new_AGEMA_signal_12629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4808 ( .C (clk), .D (new_AGEMA_signal_12632), .Q (new_AGEMA_signal_12633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4812 ( .C (clk), .D (new_AGEMA_signal_12636), .Q (new_AGEMA_signal_12637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4816 ( .C (clk), .D (new_AGEMA_signal_12640), .Q (new_AGEMA_signal_12641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4820 ( .C (clk), .D (new_AGEMA_signal_12644), .Q (new_AGEMA_signal_12645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4824 ( .C (clk), .D (new_AGEMA_signal_12648), .Q (new_AGEMA_signal_12649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4828 ( .C (clk), .D (new_AGEMA_signal_12652), .Q (new_AGEMA_signal_12653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4832 ( .C (clk), .D (new_AGEMA_signal_12656), .Q (new_AGEMA_signal_12657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4836 ( .C (clk), .D (new_AGEMA_signal_12660), .Q (new_AGEMA_signal_12661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4840 ( .C (clk), .D (new_AGEMA_signal_12664), .Q (new_AGEMA_signal_12665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4844 ( .C (clk), .D (new_AGEMA_signal_12668), .Q (new_AGEMA_signal_12669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4848 ( .C (clk), .D (new_AGEMA_signal_12672), .Q (new_AGEMA_signal_12673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4852 ( .C (clk), .D (new_AGEMA_signal_12676), .Q (new_AGEMA_signal_12677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4856 ( .C (clk), .D (new_AGEMA_signal_12680), .Q (new_AGEMA_signal_12681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4860 ( .C (clk), .D (new_AGEMA_signal_12684), .Q (new_AGEMA_signal_12685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4864 ( .C (clk), .D (new_AGEMA_signal_12688), .Q (new_AGEMA_signal_12689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4868 ( .C (clk), .D (new_AGEMA_signal_12692), .Q (new_AGEMA_signal_12693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4872 ( .C (clk), .D (new_AGEMA_signal_12696), .Q (new_AGEMA_signal_12697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4876 ( .C (clk), .D (new_AGEMA_signal_12700), .Q (new_AGEMA_signal_12701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4880 ( .C (clk), .D (new_AGEMA_signal_12704), .Q (new_AGEMA_signal_12705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4884 ( .C (clk), .D (new_AGEMA_signal_12708), .Q (new_AGEMA_signal_12709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4888 ( .C (clk), .D (new_AGEMA_signal_12712), .Q (new_AGEMA_signal_12713) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4892 ( .C (clk), .D (new_AGEMA_signal_12716), .Q (new_AGEMA_signal_12717) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4896 ( .C (clk), .D (new_AGEMA_signal_12720), .Q (new_AGEMA_signal_12721) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4900 ( .C (clk), .D (new_AGEMA_signal_12724), .Q (new_AGEMA_signal_12725) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4904 ( .C (clk), .D (new_AGEMA_signal_12728), .Q (new_AGEMA_signal_12729) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4908 ( .C (clk), .D (new_AGEMA_signal_12732), .Q (new_AGEMA_signal_12733) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4912 ( .C (clk), .D (new_AGEMA_signal_12736), .Q (new_AGEMA_signal_12737) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4916 ( .C (clk), .D (new_AGEMA_signal_12740), .Q (new_AGEMA_signal_12741) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4920 ( .C (clk), .D (new_AGEMA_signal_12744), .Q (new_AGEMA_signal_12745) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4924 ( .C (clk), .D (new_AGEMA_signal_12748), .Q (new_AGEMA_signal_12749) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4928 ( .C (clk), .D (new_AGEMA_signal_12752), .Q (new_AGEMA_signal_12753) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4932 ( .C (clk), .D (new_AGEMA_signal_12756), .Q (new_AGEMA_signal_12757) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4936 ( .C (clk), .D (new_AGEMA_signal_12760), .Q (new_AGEMA_signal_12761) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4940 ( .C (clk), .D (new_AGEMA_signal_12764), .Q (new_AGEMA_signal_12765) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4944 ( .C (clk), .D (new_AGEMA_signal_12768), .Q (new_AGEMA_signal_12769) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4948 ( .C (clk), .D (new_AGEMA_signal_12772), .Q (new_AGEMA_signal_12773) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4952 ( .C (clk), .D (new_AGEMA_signal_12776), .Q (new_AGEMA_signal_12777) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4956 ( .C (clk), .D (new_AGEMA_signal_12780), .Q (new_AGEMA_signal_12781) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4960 ( .C (clk), .D (new_AGEMA_signal_12784), .Q (new_AGEMA_signal_12785) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4964 ( .C (clk), .D (new_AGEMA_signal_12788), .Q (new_AGEMA_signal_12789) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4968 ( .C (clk), .D (new_AGEMA_signal_12792), .Q (new_AGEMA_signal_12793) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4972 ( .C (clk), .D (new_AGEMA_signal_12796), .Q (new_AGEMA_signal_12797) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4976 ( .C (clk), .D (new_AGEMA_signal_12800), .Q (new_AGEMA_signal_12801) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4980 ( .C (clk), .D (new_AGEMA_signal_12804), .Q (new_AGEMA_signal_12805) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4984 ( .C (clk), .D (new_AGEMA_signal_12808), .Q (new_AGEMA_signal_12809) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4988 ( .C (clk), .D (new_AGEMA_signal_12812), .Q (new_AGEMA_signal_12813) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4992 ( .C (clk), .D (new_AGEMA_signal_12816), .Q (new_AGEMA_signal_12817) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4996 ( .C (clk), .D (new_AGEMA_signal_12820), .Q (new_AGEMA_signal_12821) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5000 ( .C (clk), .D (new_AGEMA_signal_12824), .Q (new_AGEMA_signal_12825) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5004 ( .C (clk), .D (new_AGEMA_signal_12828), .Q (new_AGEMA_signal_12829) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5008 ( .C (clk), .D (new_AGEMA_signal_12832), .Q (new_AGEMA_signal_12833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5012 ( .C (clk), .D (new_AGEMA_signal_12836), .Q (new_AGEMA_signal_12837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5016 ( .C (clk), .D (new_AGEMA_signal_12840), .Q (new_AGEMA_signal_12841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5020 ( .C (clk), .D (new_AGEMA_signal_12844), .Q (new_AGEMA_signal_12845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5024 ( .C (clk), .D (new_AGEMA_signal_12848), .Q (new_AGEMA_signal_12849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5028 ( .C (clk), .D (new_AGEMA_signal_12852), .Q (new_AGEMA_signal_12853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5032 ( .C (clk), .D (new_AGEMA_signal_12856), .Q (new_AGEMA_signal_12857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5036 ( .C (clk), .D (new_AGEMA_signal_12860), .Q (new_AGEMA_signal_12861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5040 ( .C (clk), .D (new_AGEMA_signal_12864), .Q (new_AGEMA_signal_12865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5044 ( .C (clk), .D (new_AGEMA_signal_12868), .Q (new_AGEMA_signal_12869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5048 ( .C (clk), .D (new_AGEMA_signal_12872), .Q (new_AGEMA_signal_12873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5052 ( .C (clk), .D (new_AGEMA_signal_12876), .Q (new_AGEMA_signal_12877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5056 ( .C (clk), .D (new_AGEMA_signal_12880), .Q (new_AGEMA_signal_12881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5060 ( .C (clk), .D (new_AGEMA_signal_12884), .Q (new_AGEMA_signal_12885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5064 ( .C (clk), .D (new_AGEMA_signal_12888), .Q (new_AGEMA_signal_12889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5068 ( .C (clk), .D (new_AGEMA_signal_12892), .Q (new_AGEMA_signal_12893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5072 ( .C (clk), .D (new_AGEMA_signal_12896), .Q (new_AGEMA_signal_12897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5076 ( .C (clk), .D (new_AGEMA_signal_12900), .Q (new_AGEMA_signal_12901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5080 ( .C (clk), .D (new_AGEMA_signal_12904), .Q (new_AGEMA_signal_12905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5084 ( .C (clk), .D (new_AGEMA_signal_12908), .Q (new_AGEMA_signal_12909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5088 ( .C (clk), .D (new_AGEMA_signal_12912), .Q (new_AGEMA_signal_12913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5092 ( .C (clk), .D (new_AGEMA_signal_12916), .Q (new_AGEMA_signal_12917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5096 ( .C (clk), .D (new_AGEMA_signal_12920), .Q (new_AGEMA_signal_12921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5100 ( .C (clk), .D (new_AGEMA_signal_12924), .Q (new_AGEMA_signal_12925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5104 ( .C (clk), .D (new_AGEMA_signal_12928), .Q (new_AGEMA_signal_12929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5108 ( .C (clk), .D (new_AGEMA_signal_12932), .Q (new_AGEMA_signal_12933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5112 ( .C (clk), .D (new_AGEMA_signal_12936), .Q (new_AGEMA_signal_12937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5116 ( .C (clk), .D (new_AGEMA_signal_12940), .Q (new_AGEMA_signal_12941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5120 ( .C (clk), .D (new_AGEMA_signal_12944), .Q (new_AGEMA_signal_12945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5124 ( .C (clk), .D (new_AGEMA_signal_12948), .Q (new_AGEMA_signal_12949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5128 ( .C (clk), .D (new_AGEMA_signal_12952), .Q (new_AGEMA_signal_12953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5132 ( .C (clk), .D (new_AGEMA_signal_12956), .Q (new_AGEMA_signal_12957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5136 ( .C (clk), .D (new_AGEMA_signal_12960), .Q (new_AGEMA_signal_12961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5140 ( .C (clk), .D (new_AGEMA_signal_12964), .Q (new_AGEMA_signal_12965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5144 ( .C (clk), .D (new_AGEMA_signal_12968), .Q (new_AGEMA_signal_12969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5148 ( .C (clk), .D (new_AGEMA_signal_12972), .Q (new_AGEMA_signal_12973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5152 ( .C (clk), .D (new_AGEMA_signal_12976), .Q (new_AGEMA_signal_12977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5156 ( .C (clk), .D (new_AGEMA_signal_12980), .Q (new_AGEMA_signal_12981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5160 ( .C (clk), .D (new_AGEMA_signal_12984), .Q (new_AGEMA_signal_12985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5164 ( .C (clk), .D (new_AGEMA_signal_12988), .Q (new_AGEMA_signal_12989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5168 ( .C (clk), .D (new_AGEMA_signal_12992), .Q (new_AGEMA_signal_12993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5172 ( .C (clk), .D (new_AGEMA_signal_12996), .Q (new_AGEMA_signal_12997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5176 ( .C (clk), .D (new_AGEMA_signal_13000), .Q (new_AGEMA_signal_13001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5180 ( .C (clk), .D (new_AGEMA_signal_13004), .Q (new_AGEMA_signal_13005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5184 ( .C (clk), .D (new_AGEMA_signal_13008), .Q (new_AGEMA_signal_13009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5188 ( .C (clk), .D (new_AGEMA_signal_13012), .Q (new_AGEMA_signal_13013) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5192 ( .C (clk), .D (new_AGEMA_signal_13016), .Q (new_AGEMA_signal_13017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5196 ( .C (clk), .D (new_AGEMA_signal_13020), .Q (new_AGEMA_signal_13021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5200 ( .C (clk), .D (new_AGEMA_signal_13024), .Q (new_AGEMA_signal_13025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5204 ( .C (clk), .D (new_AGEMA_signal_13028), .Q (new_AGEMA_signal_13029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5208 ( .C (clk), .D (new_AGEMA_signal_13032), .Q (new_AGEMA_signal_13033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5212 ( .C (clk), .D (new_AGEMA_signal_13036), .Q (new_AGEMA_signal_13037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5216 ( .C (clk), .D (new_AGEMA_signal_13040), .Q (new_AGEMA_signal_13041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5220 ( .C (clk), .D (new_AGEMA_signal_13044), .Q (new_AGEMA_signal_13045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5224 ( .C (clk), .D (new_AGEMA_signal_13048), .Q (new_AGEMA_signal_13049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5228 ( .C (clk), .D (new_AGEMA_signal_13052), .Q (new_AGEMA_signal_13053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5232 ( .C (clk), .D (new_AGEMA_signal_13056), .Q (new_AGEMA_signal_13057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5236 ( .C (clk), .D (new_AGEMA_signal_13060), .Q (new_AGEMA_signal_13061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5240 ( .C (clk), .D (new_AGEMA_signal_13064), .Q (new_AGEMA_signal_13065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5244 ( .C (clk), .D (new_AGEMA_signal_13068), .Q (new_AGEMA_signal_13069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5248 ( .C (clk), .D (new_AGEMA_signal_13072), .Q (new_AGEMA_signal_13073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5252 ( .C (clk), .D (new_AGEMA_signal_13076), .Q (new_AGEMA_signal_13077) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5256 ( .C (clk), .D (new_AGEMA_signal_13080), .Q (new_AGEMA_signal_13081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5260 ( .C (clk), .D (new_AGEMA_signal_13084), .Q (new_AGEMA_signal_13085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5264 ( .C (clk), .D (new_AGEMA_signal_13088), .Q (new_AGEMA_signal_13089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5268 ( .C (clk), .D (new_AGEMA_signal_13092), .Q (new_AGEMA_signal_13093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5272 ( .C (clk), .D (new_AGEMA_signal_13096), .Q (new_AGEMA_signal_13097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5276 ( .C (clk), .D (new_AGEMA_signal_13100), .Q (new_AGEMA_signal_13101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5280 ( .C (clk), .D (new_AGEMA_signal_13104), .Q (new_AGEMA_signal_13105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5284 ( .C (clk), .D (new_AGEMA_signal_13108), .Q (new_AGEMA_signal_13109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5288 ( .C (clk), .D (new_AGEMA_signal_13112), .Q (new_AGEMA_signal_13113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5292 ( .C (clk), .D (new_AGEMA_signal_13116), .Q (new_AGEMA_signal_13117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5296 ( .C (clk), .D (new_AGEMA_signal_13120), .Q (new_AGEMA_signal_13121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5300 ( .C (clk), .D (new_AGEMA_signal_13124), .Q (new_AGEMA_signal_13125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5304 ( .C (clk), .D (new_AGEMA_signal_13128), .Q (new_AGEMA_signal_13129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5308 ( .C (clk), .D (new_AGEMA_signal_13132), .Q (new_AGEMA_signal_13133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5312 ( .C (clk), .D (new_AGEMA_signal_13136), .Q (new_AGEMA_signal_13137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5316 ( .C (clk), .D (new_AGEMA_signal_13140), .Q (new_AGEMA_signal_13141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5320 ( .C (clk), .D (new_AGEMA_signal_13144), .Q (new_AGEMA_signal_13145) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5324 ( .C (clk), .D (new_AGEMA_signal_13148), .Q (new_AGEMA_signal_13149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5328 ( .C (clk), .D (new_AGEMA_signal_13152), .Q (new_AGEMA_signal_13153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5332 ( .C (clk), .D (new_AGEMA_signal_13156), .Q (new_AGEMA_signal_13157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5336 ( .C (clk), .D (new_AGEMA_signal_13160), .Q (new_AGEMA_signal_13161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5340 ( .C (clk), .D (new_AGEMA_signal_13164), .Q (new_AGEMA_signal_13165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5344 ( .C (clk), .D (new_AGEMA_signal_13168), .Q (new_AGEMA_signal_13169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5348 ( .C (clk), .D (new_AGEMA_signal_13172), .Q (new_AGEMA_signal_13173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5352 ( .C (clk), .D (new_AGEMA_signal_13176), .Q (new_AGEMA_signal_13177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5356 ( .C (clk), .D (new_AGEMA_signal_13180), .Q (new_AGEMA_signal_13181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5360 ( .C (clk), .D (new_AGEMA_signal_13184), .Q (new_AGEMA_signal_13185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5364 ( .C (clk), .D (new_AGEMA_signal_13188), .Q (new_AGEMA_signal_13189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5368 ( .C (clk), .D (new_AGEMA_signal_13192), .Q (new_AGEMA_signal_13193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5372 ( .C (clk), .D (new_AGEMA_signal_13196), .Q (new_AGEMA_signal_13197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5376 ( .C (clk), .D (new_AGEMA_signal_13200), .Q (new_AGEMA_signal_13201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5380 ( .C (clk), .D (new_AGEMA_signal_13204), .Q (new_AGEMA_signal_13205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5384 ( .C (clk), .D (new_AGEMA_signal_13208), .Q (new_AGEMA_signal_13209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5388 ( .C (clk), .D (new_AGEMA_signal_13212), .Q (new_AGEMA_signal_13213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5392 ( .C (clk), .D (new_AGEMA_signal_13216), .Q (new_AGEMA_signal_13217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5396 ( .C (clk), .D (new_AGEMA_signal_13220), .Q (new_AGEMA_signal_13221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5400 ( .C (clk), .D (new_AGEMA_signal_13224), .Q (new_AGEMA_signal_13225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5404 ( .C (clk), .D (new_AGEMA_signal_13228), .Q (new_AGEMA_signal_13229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5408 ( .C (clk), .D (new_AGEMA_signal_13232), .Q (new_AGEMA_signal_13233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5412 ( .C (clk), .D (new_AGEMA_signal_13236), .Q (new_AGEMA_signal_13237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5416 ( .C (clk), .D (new_AGEMA_signal_13240), .Q (new_AGEMA_signal_13241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5420 ( .C (clk), .D (new_AGEMA_signal_13244), .Q (new_AGEMA_signal_13245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5424 ( .C (clk), .D (new_AGEMA_signal_13248), .Q (new_AGEMA_signal_13249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5428 ( .C (clk), .D (new_AGEMA_signal_13252), .Q (new_AGEMA_signal_13253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5432 ( .C (clk), .D (new_AGEMA_signal_13256), .Q (new_AGEMA_signal_13257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5436 ( .C (clk), .D (new_AGEMA_signal_13260), .Q (new_AGEMA_signal_13261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5440 ( .C (clk), .D (new_AGEMA_signal_13264), .Q (new_AGEMA_signal_13265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5444 ( .C (clk), .D (new_AGEMA_signal_13268), .Q (new_AGEMA_signal_13269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5448 ( .C (clk), .D (new_AGEMA_signal_13272), .Q (new_AGEMA_signal_13273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5452 ( .C (clk), .D (new_AGEMA_signal_13276), .Q (new_AGEMA_signal_13277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5456 ( .C (clk), .D (new_AGEMA_signal_13280), .Q (new_AGEMA_signal_13281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5460 ( .C (clk), .D (new_AGEMA_signal_13284), .Q (new_AGEMA_signal_13285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5464 ( .C (clk), .D (new_AGEMA_signal_13288), .Q (new_AGEMA_signal_13289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5468 ( .C (clk), .D (new_AGEMA_signal_13292), .Q (new_AGEMA_signal_13293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5472 ( .C (clk), .D (new_AGEMA_signal_13296), .Q (new_AGEMA_signal_13297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5476 ( .C (clk), .D (new_AGEMA_signal_13300), .Q (new_AGEMA_signal_13301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5480 ( .C (clk), .D (new_AGEMA_signal_13304), .Q (new_AGEMA_signal_13305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5484 ( .C (clk), .D (new_AGEMA_signal_13308), .Q (new_AGEMA_signal_13309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5488 ( .C (clk), .D (new_AGEMA_signal_13312), .Q (new_AGEMA_signal_13313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5492 ( .C (clk), .D (new_AGEMA_signal_13316), .Q (new_AGEMA_signal_13317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5496 ( .C (clk), .D (new_AGEMA_signal_13320), .Q (new_AGEMA_signal_13321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5500 ( .C (clk), .D (new_AGEMA_signal_13324), .Q (new_AGEMA_signal_13325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5504 ( .C (clk), .D (new_AGEMA_signal_13328), .Q (new_AGEMA_signal_13329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5508 ( .C (clk), .D (new_AGEMA_signal_13332), .Q (new_AGEMA_signal_13333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5512 ( .C (clk), .D (new_AGEMA_signal_13336), .Q (new_AGEMA_signal_13337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5516 ( .C (clk), .D (new_AGEMA_signal_13340), .Q (new_AGEMA_signal_13341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5520 ( .C (clk), .D (new_AGEMA_signal_13344), .Q (new_AGEMA_signal_13345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5524 ( .C (clk), .D (new_AGEMA_signal_13348), .Q (new_AGEMA_signal_13349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5528 ( .C (clk), .D (new_AGEMA_signal_13352), .Q (new_AGEMA_signal_13353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5532 ( .C (clk), .D (new_AGEMA_signal_13356), .Q (new_AGEMA_signal_13357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5536 ( .C (clk), .D (new_AGEMA_signal_13360), .Q (new_AGEMA_signal_13361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5540 ( .C (clk), .D (new_AGEMA_signal_13364), .Q (new_AGEMA_signal_13365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5544 ( .C (clk), .D (new_AGEMA_signal_13368), .Q (new_AGEMA_signal_13369) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5548 ( .C (clk), .D (new_AGEMA_signal_13372), .Q (new_AGEMA_signal_13373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5552 ( .C (clk), .D (new_AGEMA_signal_13376), .Q (new_AGEMA_signal_13377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5556 ( .C (clk), .D (new_AGEMA_signal_13380), .Q (new_AGEMA_signal_13381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5560 ( .C (clk), .D (new_AGEMA_signal_13384), .Q (new_AGEMA_signal_13385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5564 ( .C (clk), .D (new_AGEMA_signal_13388), .Q (new_AGEMA_signal_13389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5568 ( .C (clk), .D (new_AGEMA_signal_13392), .Q (new_AGEMA_signal_13393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5572 ( .C (clk), .D (new_AGEMA_signal_13396), .Q (new_AGEMA_signal_13397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5576 ( .C (clk), .D (new_AGEMA_signal_13400), .Q (new_AGEMA_signal_13401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5580 ( .C (clk), .D (new_AGEMA_signal_13404), .Q (new_AGEMA_signal_13405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5584 ( .C (clk), .D (new_AGEMA_signal_13408), .Q (new_AGEMA_signal_13409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5588 ( .C (clk), .D (new_AGEMA_signal_13412), .Q (new_AGEMA_signal_13413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5592 ( .C (clk), .D (new_AGEMA_signal_13416), .Q (new_AGEMA_signal_13417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5596 ( .C (clk), .D (new_AGEMA_signal_13420), .Q (new_AGEMA_signal_13421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5600 ( .C (clk), .D (new_AGEMA_signal_13424), .Q (new_AGEMA_signal_13425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5604 ( .C (clk), .D (new_AGEMA_signal_13428), .Q (new_AGEMA_signal_13429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5608 ( .C (clk), .D (new_AGEMA_signal_13432), .Q (new_AGEMA_signal_13433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5612 ( .C (clk), .D (new_AGEMA_signal_13436), .Q (new_AGEMA_signal_13437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5616 ( .C (clk), .D (new_AGEMA_signal_13440), .Q (new_AGEMA_signal_13441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5620 ( .C (clk), .D (new_AGEMA_signal_13444), .Q (new_AGEMA_signal_13445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5624 ( .C (clk), .D (new_AGEMA_signal_13448), .Q (new_AGEMA_signal_13449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5628 ( .C (clk), .D (new_AGEMA_signal_13452), .Q (new_AGEMA_signal_13453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5632 ( .C (clk), .D (new_AGEMA_signal_13456), .Q (new_AGEMA_signal_13457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5636 ( .C (clk), .D (new_AGEMA_signal_13460), .Q (new_AGEMA_signal_13461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5640 ( .C (clk), .D (new_AGEMA_signal_13464), .Q (new_AGEMA_signal_13465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5644 ( .C (clk), .D (new_AGEMA_signal_13468), .Q (new_AGEMA_signal_13469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5648 ( .C (clk), .D (new_AGEMA_signal_13472), .Q (new_AGEMA_signal_13473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5652 ( .C (clk), .D (new_AGEMA_signal_13476), .Q (new_AGEMA_signal_13477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5656 ( .C (clk), .D (new_AGEMA_signal_13480), .Q (new_AGEMA_signal_13481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5660 ( .C (clk), .D (new_AGEMA_signal_13484), .Q (new_AGEMA_signal_13485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5664 ( .C (clk), .D (new_AGEMA_signal_13488), .Q (new_AGEMA_signal_13489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5668 ( .C (clk), .D (new_AGEMA_signal_13492), .Q (new_AGEMA_signal_13493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5672 ( .C (clk), .D (new_AGEMA_signal_13496), .Q (new_AGEMA_signal_13497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5676 ( .C (clk), .D (new_AGEMA_signal_13500), .Q (new_AGEMA_signal_13501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5680 ( .C (clk), .D (new_AGEMA_signal_13504), .Q (new_AGEMA_signal_13505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5684 ( .C (clk), .D (new_AGEMA_signal_13508), .Q (new_AGEMA_signal_13509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5688 ( .C (clk), .D (new_AGEMA_signal_13512), .Q (new_AGEMA_signal_13513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5692 ( .C (clk), .D (new_AGEMA_signal_13516), .Q (new_AGEMA_signal_13517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5696 ( .C (clk), .D (new_AGEMA_signal_13520), .Q (new_AGEMA_signal_13521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5700 ( .C (clk), .D (new_AGEMA_signal_13524), .Q (new_AGEMA_signal_13525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5704 ( .C (clk), .D (new_AGEMA_signal_13528), .Q (new_AGEMA_signal_13529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5708 ( .C (clk), .D (new_AGEMA_signal_13532), .Q (new_AGEMA_signal_13533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5712 ( .C (clk), .D (new_AGEMA_signal_13536), .Q (new_AGEMA_signal_13537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5716 ( .C (clk), .D (new_AGEMA_signal_13540), .Q (new_AGEMA_signal_13541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5720 ( .C (clk), .D (new_AGEMA_signal_13544), .Q (new_AGEMA_signal_13545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5724 ( .C (clk), .D (new_AGEMA_signal_13548), .Q (new_AGEMA_signal_13549) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5728 ( .C (clk), .D (new_AGEMA_signal_13552), .Q (new_AGEMA_signal_13553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5732 ( .C (clk), .D (new_AGEMA_signal_13556), .Q (new_AGEMA_signal_13557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5736 ( .C (clk), .D (new_AGEMA_signal_13560), .Q (new_AGEMA_signal_13561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5740 ( .C (clk), .D (new_AGEMA_signal_13564), .Q (new_AGEMA_signal_13565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5744 ( .C (clk), .D (new_AGEMA_signal_13568), .Q (new_AGEMA_signal_13569) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5748 ( .C (clk), .D (new_AGEMA_signal_13572), .Q (new_AGEMA_signal_13573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5752 ( .C (clk), .D (new_AGEMA_signal_13576), .Q (new_AGEMA_signal_13577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5756 ( .C (clk), .D (new_AGEMA_signal_13580), .Q (new_AGEMA_signal_13581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5760 ( .C (clk), .D (new_AGEMA_signal_13584), .Q (new_AGEMA_signal_13585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5764 ( .C (clk), .D (new_AGEMA_signal_13588), .Q (new_AGEMA_signal_13589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5768 ( .C (clk), .D (new_AGEMA_signal_13592), .Q (new_AGEMA_signal_13593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5772 ( .C (clk), .D (new_AGEMA_signal_13596), .Q (new_AGEMA_signal_13597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5776 ( .C (clk), .D (new_AGEMA_signal_13600), .Q (new_AGEMA_signal_13601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5780 ( .C (clk), .D (new_AGEMA_signal_13604), .Q (new_AGEMA_signal_13605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5784 ( .C (clk), .D (new_AGEMA_signal_13608), .Q (new_AGEMA_signal_13609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5788 ( .C (clk), .D (new_AGEMA_signal_13612), .Q (new_AGEMA_signal_13613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5792 ( .C (clk), .D (new_AGEMA_signal_13616), .Q (new_AGEMA_signal_13617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5796 ( .C (clk), .D (new_AGEMA_signal_13620), .Q (new_AGEMA_signal_13621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5800 ( .C (clk), .D (new_AGEMA_signal_13624), .Q (new_AGEMA_signal_13625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5804 ( .C (clk), .D (new_AGEMA_signal_13628), .Q (new_AGEMA_signal_13629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5808 ( .C (clk), .D (new_AGEMA_signal_13632), .Q (new_AGEMA_signal_13633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5812 ( .C (clk), .D (new_AGEMA_signal_13636), .Q (new_AGEMA_signal_13637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5816 ( .C (clk), .D (new_AGEMA_signal_13640), .Q (new_AGEMA_signal_13641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5820 ( .C (clk), .D (new_AGEMA_signal_13644), .Q (new_AGEMA_signal_13645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5824 ( .C (clk), .D (new_AGEMA_signal_13648), .Q (new_AGEMA_signal_13649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5828 ( .C (clk), .D (new_AGEMA_signal_13652), .Q (new_AGEMA_signal_13653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5832 ( .C (clk), .D (new_AGEMA_signal_13656), .Q (new_AGEMA_signal_13657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5836 ( .C (clk), .D (new_AGEMA_signal_13660), .Q (new_AGEMA_signal_13661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5840 ( .C (clk), .D (new_AGEMA_signal_13664), .Q (new_AGEMA_signal_13665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5844 ( .C (clk), .D (new_AGEMA_signal_13668), .Q (new_AGEMA_signal_13669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5848 ( .C (clk), .D (new_AGEMA_signal_13672), .Q (new_AGEMA_signal_13673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5852 ( .C (clk), .D (new_AGEMA_signal_13676), .Q (new_AGEMA_signal_13677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5856 ( .C (clk), .D (new_AGEMA_signal_13680), .Q (new_AGEMA_signal_13681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5860 ( .C (clk), .D (new_AGEMA_signal_13684), .Q (new_AGEMA_signal_13685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5864 ( .C (clk), .D (new_AGEMA_signal_13688), .Q (new_AGEMA_signal_13689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5868 ( .C (clk), .D (new_AGEMA_signal_13692), .Q (new_AGEMA_signal_13693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5872 ( .C (clk), .D (new_AGEMA_signal_13696), .Q (new_AGEMA_signal_13697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5876 ( .C (clk), .D (new_AGEMA_signal_13700), .Q (new_AGEMA_signal_13701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5880 ( .C (clk), .D (new_AGEMA_signal_13704), .Q (new_AGEMA_signal_13705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5884 ( .C (clk), .D (new_AGEMA_signal_13708), .Q (new_AGEMA_signal_13709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5888 ( .C (clk), .D (new_AGEMA_signal_13712), .Q (new_AGEMA_signal_13713) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5892 ( .C (clk), .D (new_AGEMA_signal_13716), .Q (new_AGEMA_signal_13717) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5896 ( .C (clk), .D (new_AGEMA_signal_13720), .Q (new_AGEMA_signal_13721) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5900 ( .C (clk), .D (new_AGEMA_signal_13724), .Q (new_AGEMA_signal_13725) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5904 ( .C (clk), .D (new_AGEMA_signal_13728), .Q (new_AGEMA_signal_13729) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5908 ( .C (clk), .D (new_AGEMA_signal_13732), .Q (new_AGEMA_signal_13733) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5912 ( .C (clk), .D (new_AGEMA_signal_13736), .Q (new_AGEMA_signal_13737) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5916 ( .C (clk), .D (new_AGEMA_signal_13740), .Q (new_AGEMA_signal_13741) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5920 ( .C (clk), .D (new_AGEMA_signal_13744), .Q (new_AGEMA_signal_13745) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5924 ( .C (clk), .D (new_AGEMA_signal_13748), .Q (new_AGEMA_signal_13749) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5928 ( .C (clk), .D (new_AGEMA_signal_13752), .Q (new_AGEMA_signal_13753) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5932 ( .C (clk), .D (new_AGEMA_signal_13756), .Q (new_AGEMA_signal_13757) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5936 ( .C (clk), .D (new_AGEMA_signal_13760), .Q (new_AGEMA_signal_13761) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5940 ( .C (clk), .D (new_AGEMA_signal_13764), .Q (new_AGEMA_signal_13765) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5944 ( .C (clk), .D (new_AGEMA_signal_13768), .Q (new_AGEMA_signal_13769) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5948 ( .C (clk), .D (new_AGEMA_signal_13772), .Q (new_AGEMA_signal_13773) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5952 ( .C (clk), .D (new_AGEMA_signal_13776), .Q (new_AGEMA_signal_13777) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5956 ( .C (clk), .D (new_AGEMA_signal_13780), .Q (new_AGEMA_signal_13781) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5960 ( .C (clk), .D (new_AGEMA_signal_13784), .Q (new_AGEMA_signal_13785) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5964 ( .C (clk), .D (new_AGEMA_signal_13788), .Q (new_AGEMA_signal_13789) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5968 ( .C (clk), .D (new_AGEMA_signal_13792), .Q (new_AGEMA_signal_13793) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5972 ( .C (clk), .D (new_AGEMA_signal_13796), .Q (new_AGEMA_signal_13797) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5976 ( .C (clk), .D (new_AGEMA_signal_13800), .Q (new_AGEMA_signal_13801) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5980 ( .C (clk), .D (new_AGEMA_signal_13804), .Q (new_AGEMA_signal_13805) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5984 ( .C (clk), .D (new_AGEMA_signal_13808), .Q (new_AGEMA_signal_13809) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5988 ( .C (clk), .D (new_AGEMA_signal_13812), .Q (new_AGEMA_signal_13813) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5992 ( .C (clk), .D (new_AGEMA_signal_13816), .Q (new_AGEMA_signal_13817) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5996 ( .C (clk), .D (new_AGEMA_signal_13820), .Q (new_AGEMA_signal_13821) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6000 ( .C (clk), .D (new_AGEMA_signal_13824), .Q (new_AGEMA_signal_13825) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6004 ( .C (clk), .D (new_AGEMA_signal_13828), .Q (new_AGEMA_signal_13829) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6008 ( .C (clk), .D (new_AGEMA_signal_13832), .Q (new_AGEMA_signal_13833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6012 ( .C (clk), .D (new_AGEMA_signal_13836), .Q (new_AGEMA_signal_13837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6016 ( .C (clk), .D (new_AGEMA_signal_13840), .Q (new_AGEMA_signal_13841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6020 ( .C (clk), .D (new_AGEMA_signal_13844), .Q (new_AGEMA_signal_13845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6024 ( .C (clk), .D (new_AGEMA_signal_13848), .Q (new_AGEMA_signal_13849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6028 ( .C (clk), .D (new_AGEMA_signal_13852), .Q (new_AGEMA_signal_13853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6032 ( .C (clk), .D (new_AGEMA_signal_13856), .Q (new_AGEMA_signal_13857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6036 ( .C (clk), .D (new_AGEMA_signal_13860), .Q (new_AGEMA_signal_13861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6040 ( .C (clk), .D (new_AGEMA_signal_13864), .Q (new_AGEMA_signal_13865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6044 ( .C (clk), .D (new_AGEMA_signal_13868), .Q (new_AGEMA_signal_13869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6048 ( .C (clk), .D (new_AGEMA_signal_13872), .Q (new_AGEMA_signal_13873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6052 ( .C (clk), .D (new_AGEMA_signal_13876), .Q (new_AGEMA_signal_13877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6056 ( .C (clk), .D (new_AGEMA_signal_13880), .Q (new_AGEMA_signal_13881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6060 ( .C (clk), .D (new_AGEMA_signal_13884), .Q (new_AGEMA_signal_13885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6064 ( .C (clk), .D (new_AGEMA_signal_13888), .Q (new_AGEMA_signal_13889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6068 ( .C (clk), .D (new_AGEMA_signal_13892), .Q (new_AGEMA_signal_13893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6072 ( .C (clk), .D (new_AGEMA_signal_13896), .Q (new_AGEMA_signal_13897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6076 ( .C (clk), .D (new_AGEMA_signal_13900), .Q (new_AGEMA_signal_13901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6080 ( .C (clk), .D (new_AGEMA_signal_13904), .Q (new_AGEMA_signal_13905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6084 ( .C (clk), .D (new_AGEMA_signal_13908), .Q (new_AGEMA_signal_13909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6088 ( .C (clk), .D (new_AGEMA_signal_13912), .Q (new_AGEMA_signal_13913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6092 ( .C (clk), .D (new_AGEMA_signal_13916), .Q (new_AGEMA_signal_13917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6096 ( .C (clk), .D (new_AGEMA_signal_13920), .Q (new_AGEMA_signal_13921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6100 ( .C (clk), .D (new_AGEMA_signal_13924), .Q (new_AGEMA_signal_13925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6104 ( .C (clk), .D (new_AGEMA_signal_13928), .Q (new_AGEMA_signal_13929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6108 ( .C (clk), .D (new_AGEMA_signal_13932), .Q (new_AGEMA_signal_13933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6112 ( .C (clk), .D (new_AGEMA_signal_13936), .Q (new_AGEMA_signal_13937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6116 ( .C (clk), .D (new_AGEMA_signal_13940), .Q (new_AGEMA_signal_13941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6120 ( .C (clk), .D (new_AGEMA_signal_13944), .Q (new_AGEMA_signal_13945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6124 ( .C (clk), .D (new_AGEMA_signal_13948), .Q (new_AGEMA_signal_13949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6128 ( .C (clk), .D (new_AGEMA_signal_13952), .Q (new_AGEMA_signal_13953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6132 ( .C (clk), .D (new_AGEMA_signal_13956), .Q (new_AGEMA_signal_13957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6136 ( .C (clk), .D (new_AGEMA_signal_13960), .Q (new_AGEMA_signal_13961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6140 ( .C (clk), .D (new_AGEMA_signal_13964), .Q (new_AGEMA_signal_13965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6144 ( .C (clk), .D (new_AGEMA_signal_13968), .Q (new_AGEMA_signal_13969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6148 ( .C (clk), .D (new_AGEMA_signal_13972), .Q (new_AGEMA_signal_13973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6152 ( .C (clk), .D (new_AGEMA_signal_13976), .Q (new_AGEMA_signal_13977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6156 ( .C (clk), .D (new_AGEMA_signal_13980), .Q (new_AGEMA_signal_13981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6160 ( .C (clk), .D (new_AGEMA_signal_13984), .Q (new_AGEMA_signal_13985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6164 ( .C (clk), .D (new_AGEMA_signal_13988), .Q (new_AGEMA_signal_13989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6168 ( .C (clk), .D (new_AGEMA_signal_13992), .Q (new_AGEMA_signal_13993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6172 ( .C (clk), .D (new_AGEMA_signal_13996), .Q (new_AGEMA_signal_13997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6176 ( .C (clk), .D (new_AGEMA_signal_14000), .Q (new_AGEMA_signal_14001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6180 ( .C (clk), .D (new_AGEMA_signal_14004), .Q (new_AGEMA_signal_14005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6184 ( .C (clk), .D (new_AGEMA_signal_14008), .Q (new_AGEMA_signal_14009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6188 ( .C (clk), .D (new_AGEMA_signal_14012), .Q (new_AGEMA_signal_14013) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6192 ( .C (clk), .D (new_AGEMA_signal_14016), .Q (new_AGEMA_signal_14017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6196 ( .C (clk), .D (new_AGEMA_signal_14020), .Q (new_AGEMA_signal_14021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6200 ( .C (clk), .D (new_AGEMA_signal_14024), .Q (new_AGEMA_signal_14025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6204 ( .C (clk), .D (new_AGEMA_signal_14028), .Q (new_AGEMA_signal_14029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6208 ( .C (clk), .D (new_AGEMA_signal_14032), .Q (new_AGEMA_signal_14033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6212 ( .C (clk), .D (new_AGEMA_signal_14036), .Q (new_AGEMA_signal_14037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6216 ( .C (clk), .D (new_AGEMA_signal_14040), .Q (new_AGEMA_signal_14041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6220 ( .C (clk), .D (new_AGEMA_signal_14044), .Q (new_AGEMA_signal_14045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6224 ( .C (clk), .D (new_AGEMA_signal_14048), .Q (new_AGEMA_signal_14049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6228 ( .C (clk), .D (new_AGEMA_signal_14052), .Q (new_AGEMA_signal_14053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6232 ( .C (clk), .D (new_AGEMA_signal_14056), .Q (new_AGEMA_signal_14057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6236 ( .C (clk), .D (new_AGEMA_signal_14060), .Q (new_AGEMA_signal_14061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6240 ( .C (clk), .D (new_AGEMA_signal_14064), .Q (new_AGEMA_signal_14065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6244 ( .C (clk), .D (new_AGEMA_signal_14068), .Q (new_AGEMA_signal_14069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6248 ( .C (clk), .D (new_AGEMA_signal_14072), .Q (new_AGEMA_signal_14073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6252 ( .C (clk), .D (new_AGEMA_signal_14076), .Q (new_AGEMA_signal_14077) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6256 ( .C (clk), .D (new_AGEMA_signal_14080), .Q (new_AGEMA_signal_14081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6260 ( .C (clk), .D (new_AGEMA_signal_14084), .Q (new_AGEMA_signal_14085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6264 ( .C (clk), .D (new_AGEMA_signal_14088), .Q (new_AGEMA_signal_14089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6268 ( .C (clk), .D (new_AGEMA_signal_14092), .Q (new_AGEMA_signal_14093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6272 ( .C (clk), .D (new_AGEMA_signal_14096), .Q (new_AGEMA_signal_14097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6276 ( .C (clk), .D (new_AGEMA_signal_14100), .Q (new_AGEMA_signal_14101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6280 ( .C (clk), .D (new_AGEMA_signal_14104), .Q (new_AGEMA_signal_14105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6284 ( .C (clk), .D (new_AGEMA_signal_14108), .Q (new_AGEMA_signal_14109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6288 ( .C (clk), .D (new_AGEMA_signal_14112), .Q (new_AGEMA_signal_14113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6292 ( .C (clk), .D (new_AGEMA_signal_14116), .Q (new_AGEMA_signal_14117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6296 ( .C (clk), .D (new_AGEMA_signal_14120), .Q (new_AGEMA_signal_14121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6300 ( .C (clk), .D (new_AGEMA_signal_14124), .Q (new_AGEMA_signal_14125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6304 ( .C (clk), .D (new_AGEMA_signal_14128), .Q (new_AGEMA_signal_14129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6308 ( .C (clk), .D (new_AGEMA_signal_14132), .Q (new_AGEMA_signal_14133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6312 ( .C (clk), .D (new_AGEMA_signal_14136), .Q (new_AGEMA_signal_14137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6316 ( .C (clk), .D (new_AGEMA_signal_14140), .Q (new_AGEMA_signal_14141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6320 ( .C (clk), .D (new_AGEMA_signal_14144), .Q (new_AGEMA_signal_14145) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6324 ( .C (clk), .D (new_AGEMA_signal_14148), .Q (new_AGEMA_signal_14149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6328 ( .C (clk), .D (new_AGEMA_signal_14152), .Q (new_AGEMA_signal_14153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6332 ( .C (clk), .D (new_AGEMA_signal_14156), .Q (new_AGEMA_signal_14157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6336 ( .C (clk), .D (new_AGEMA_signal_14160), .Q (new_AGEMA_signal_14161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6340 ( .C (clk), .D (new_AGEMA_signal_14164), .Q (new_AGEMA_signal_14165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6344 ( .C (clk), .D (new_AGEMA_signal_14168), .Q (new_AGEMA_signal_14169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6348 ( .C (clk), .D (new_AGEMA_signal_14172), .Q (new_AGEMA_signal_14173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6352 ( .C (clk), .D (new_AGEMA_signal_14176), .Q (new_AGEMA_signal_14177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6356 ( .C (clk), .D (new_AGEMA_signal_14180), .Q (new_AGEMA_signal_14181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6360 ( .C (clk), .D (new_AGEMA_signal_14184), .Q (new_AGEMA_signal_14185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6364 ( .C (clk), .D (new_AGEMA_signal_14188), .Q (new_AGEMA_signal_14189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6368 ( .C (clk), .D (new_AGEMA_signal_14192), .Q (new_AGEMA_signal_14193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6372 ( .C (clk), .D (new_AGEMA_signal_14196), .Q (new_AGEMA_signal_14197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6376 ( .C (clk), .D (new_AGEMA_signal_14200), .Q (new_AGEMA_signal_14201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6380 ( .C (clk), .D (new_AGEMA_signal_14204), .Q (new_AGEMA_signal_14205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6384 ( .C (clk), .D (new_AGEMA_signal_14208), .Q (new_AGEMA_signal_14209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6388 ( .C (clk), .D (new_AGEMA_signal_14212), .Q (new_AGEMA_signal_14213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6392 ( .C (clk), .D (new_AGEMA_signal_14216), .Q (new_AGEMA_signal_14217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6396 ( .C (clk), .D (new_AGEMA_signal_14220), .Q (new_AGEMA_signal_14221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6400 ( .C (clk), .D (new_AGEMA_signal_14224), .Q (new_AGEMA_signal_14225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6404 ( .C (clk), .D (new_AGEMA_signal_14228), .Q (new_AGEMA_signal_14229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6408 ( .C (clk), .D (new_AGEMA_signal_14232), .Q (new_AGEMA_signal_14233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6412 ( .C (clk), .D (new_AGEMA_signal_14236), .Q (new_AGEMA_signal_14237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6416 ( .C (clk), .D (new_AGEMA_signal_14240), .Q (new_AGEMA_signal_14241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6420 ( .C (clk), .D (new_AGEMA_signal_14244), .Q (new_AGEMA_signal_14245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6424 ( .C (clk), .D (new_AGEMA_signal_14248), .Q (new_AGEMA_signal_14249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6428 ( .C (clk), .D (new_AGEMA_signal_14252), .Q (new_AGEMA_signal_14253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6432 ( .C (clk), .D (new_AGEMA_signal_14256), .Q (new_AGEMA_signal_14257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6436 ( .C (clk), .D (new_AGEMA_signal_14260), .Q (new_AGEMA_signal_14261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6440 ( .C (clk), .D (new_AGEMA_signal_14264), .Q (new_AGEMA_signal_14265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6444 ( .C (clk), .D (new_AGEMA_signal_14268), .Q (new_AGEMA_signal_14269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6448 ( .C (clk), .D (new_AGEMA_signal_14272), .Q (new_AGEMA_signal_14273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6452 ( .C (clk), .D (new_AGEMA_signal_14276), .Q (new_AGEMA_signal_14277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6456 ( .C (clk), .D (new_AGEMA_signal_14280), .Q (new_AGEMA_signal_14281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6460 ( .C (clk), .D (new_AGEMA_signal_14284), .Q (new_AGEMA_signal_14285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6464 ( .C (clk), .D (new_AGEMA_signal_14288), .Q (new_AGEMA_signal_14289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6468 ( .C (clk), .D (new_AGEMA_signal_14292), .Q (new_AGEMA_signal_14293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6472 ( .C (clk), .D (new_AGEMA_signal_14296), .Q (new_AGEMA_signal_14297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6476 ( .C (clk), .D (new_AGEMA_signal_14300), .Q (new_AGEMA_signal_14301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6480 ( .C (clk), .D (new_AGEMA_signal_14304), .Q (new_AGEMA_signal_14305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6484 ( .C (clk), .D (new_AGEMA_signal_14308), .Q (new_AGEMA_signal_14309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6488 ( .C (clk), .D (new_AGEMA_signal_14312), .Q (new_AGEMA_signal_14313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6492 ( .C (clk), .D (new_AGEMA_signal_14316), .Q (new_AGEMA_signal_14317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6496 ( .C (clk), .D (new_AGEMA_signal_14320), .Q (new_AGEMA_signal_14321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6500 ( .C (clk), .D (new_AGEMA_signal_14324), .Q (new_AGEMA_signal_14325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6504 ( .C (clk), .D (new_AGEMA_signal_14328), .Q (new_AGEMA_signal_14329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6508 ( .C (clk), .D (new_AGEMA_signal_14332), .Q (new_AGEMA_signal_14333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6512 ( .C (clk), .D (new_AGEMA_signal_14336), .Q (new_AGEMA_signal_14337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6516 ( .C (clk), .D (new_AGEMA_signal_14340), .Q (new_AGEMA_signal_14341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6520 ( .C (clk), .D (new_AGEMA_signal_14344), .Q (new_AGEMA_signal_14345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6524 ( .C (clk), .D (new_AGEMA_signal_14348), .Q (new_AGEMA_signal_14349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6528 ( .C (clk), .D (new_AGEMA_signal_14352), .Q (new_AGEMA_signal_14353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6532 ( .C (clk), .D (new_AGEMA_signal_14356), .Q (new_AGEMA_signal_14357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6536 ( .C (clk), .D (new_AGEMA_signal_14360), .Q (new_AGEMA_signal_14361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6540 ( .C (clk), .D (new_AGEMA_signal_14364), .Q (new_AGEMA_signal_14365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6544 ( .C (clk), .D (new_AGEMA_signal_14368), .Q (new_AGEMA_signal_14369) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6548 ( .C (clk), .D (new_AGEMA_signal_14372), .Q (new_AGEMA_signal_14373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6552 ( .C (clk), .D (new_AGEMA_signal_14376), .Q (new_AGEMA_signal_14377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6556 ( .C (clk), .D (new_AGEMA_signal_14380), .Q (new_AGEMA_signal_14381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6560 ( .C (clk), .D (new_AGEMA_signal_14384), .Q (new_AGEMA_signal_14385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6564 ( .C (clk), .D (new_AGEMA_signal_14388), .Q (new_AGEMA_signal_14389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6568 ( .C (clk), .D (new_AGEMA_signal_14392), .Q (new_AGEMA_signal_14393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6572 ( .C (clk), .D (new_AGEMA_signal_14396), .Q (new_AGEMA_signal_14397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6576 ( .C (clk), .D (new_AGEMA_signal_14400), .Q (new_AGEMA_signal_14401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6580 ( .C (clk), .D (new_AGEMA_signal_14404), .Q (new_AGEMA_signal_14405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6584 ( .C (clk), .D (new_AGEMA_signal_14408), .Q (new_AGEMA_signal_14409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6588 ( .C (clk), .D (new_AGEMA_signal_14412), .Q (new_AGEMA_signal_14413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6592 ( .C (clk), .D (new_AGEMA_signal_14416), .Q (new_AGEMA_signal_14417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6596 ( .C (clk), .D (new_AGEMA_signal_14420), .Q (new_AGEMA_signal_14421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6600 ( .C (clk), .D (new_AGEMA_signal_14424), .Q (new_AGEMA_signal_14425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6604 ( .C (clk), .D (new_AGEMA_signal_14428), .Q (new_AGEMA_signal_14429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6608 ( .C (clk), .D (new_AGEMA_signal_14432), .Q (new_AGEMA_signal_14433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6612 ( .C (clk), .D (new_AGEMA_signal_14436), .Q (new_AGEMA_signal_14437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6616 ( .C (clk), .D (new_AGEMA_signal_14440), .Q (new_AGEMA_signal_14441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6620 ( .C (clk), .D (new_AGEMA_signal_14444), .Q (new_AGEMA_signal_14445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6624 ( .C (clk), .D (new_AGEMA_signal_14448), .Q (new_AGEMA_signal_14449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6628 ( .C (clk), .D (new_AGEMA_signal_14452), .Q (new_AGEMA_signal_14453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6632 ( .C (clk), .D (new_AGEMA_signal_14456), .Q (new_AGEMA_signal_14457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6636 ( .C (clk), .D (new_AGEMA_signal_14460), .Q (new_AGEMA_signal_14461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6640 ( .C (clk), .D (new_AGEMA_signal_14464), .Q (new_AGEMA_signal_14465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6644 ( .C (clk), .D (new_AGEMA_signal_14468), .Q (new_AGEMA_signal_14469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6648 ( .C (clk), .D (new_AGEMA_signal_14472), .Q (new_AGEMA_signal_14473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6652 ( .C (clk), .D (new_AGEMA_signal_14476), .Q (new_AGEMA_signal_14477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6656 ( .C (clk), .D (new_AGEMA_signal_14480), .Q (new_AGEMA_signal_14481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6660 ( .C (clk), .D (new_AGEMA_signal_14484), .Q (new_AGEMA_signal_14485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6664 ( .C (clk), .D (new_AGEMA_signal_14488), .Q (new_AGEMA_signal_14489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6668 ( .C (clk), .D (new_AGEMA_signal_14492), .Q (new_AGEMA_signal_14493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6672 ( .C (clk), .D (new_AGEMA_signal_14496), .Q (new_AGEMA_signal_14497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6676 ( .C (clk), .D (new_AGEMA_signal_14500), .Q (new_AGEMA_signal_14501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6680 ( .C (clk), .D (new_AGEMA_signal_14504), .Q (new_AGEMA_signal_14505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6684 ( .C (clk), .D (new_AGEMA_signal_14508), .Q (new_AGEMA_signal_14509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6688 ( .C (clk), .D (new_AGEMA_signal_14512), .Q (new_AGEMA_signal_14513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6692 ( .C (clk), .D (new_AGEMA_signal_14516), .Q (new_AGEMA_signal_14517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6696 ( .C (clk), .D (new_AGEMA_signal_14520), .Q (new_AGEMA_signal_14521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6700 ( .C (clk), .D (new_AGEMA_signal_14524), .Q (new_AGEMA_signal_14525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6704 ( .C (clk), .D (new_AGEMA_signal_14528), .Q (new_AGEMA_signal_14529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6708 ( .C (clk), .D (new_AGEMA_signal_14532), .Q (new_AGEMA_signal_14533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6712 ( .C (clk), .D (new_AGEMA_signal_14536), .Q (new_AGEMA_signal_14537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6716 ( .C (clk), .D (new_AGEMA_signal_14540), .Q (new_AGEMA_signal_14541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6720 ( .C (clk), .D (new_AGEMA_signal_14544), .Q (new_AGEMA_signal_14545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6724 ( .C (clk), .D (new_AGEMA_signal_14548), .Q (new_AGEMA_signal_14549) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6728 ( .C (clk), .D (new_AGEMA_signal_14552), .Q (new_AGEMA_signal_14553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6732 ( .C (clk), .D (new_AGEMA_signal_14556), .Q (new_AGEMA_signal_14557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6736 ( .C (clk), .D (new_AGEMA_signal_14560), .Q (new_AGEMA_signal_14561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6740 ( .C (clk), .D (new_AGEMA_signal_14564), .Q (new_AGEMA_signal_14565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6744 ( .C (clk), .D (new_AGEMA_signal_14568), .Q (new_AGEMA_signal_14569) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6748 ( .C (clk), .D (new_AGEMA_signal_14572), .Q (new_AGEMA_signal_14573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6752 ( .C (clk), .D (new_AGEMA_signal_14576), .Q (new_AGEMA_signal_14577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6756 ( .C (clk), .D (new_AGEMA_signal_14580), .Q (new_AGEMA_signal_14581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6760 ( .C (clk), .D (new_AGEMA_signal_14584), .Q (new_AGEMA_signal_14585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6764 ( .C (clk), .D (new_AGEMA_signal_14588), .Q (new_AGEMA_signal_14589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6768 ( .C (clk), .D (new_AGEMA_signal_14592), .Q (new_AGEMA_signal_14593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6772 ( .C (clk), .D (new_AGEMA_signal_14596), .Q (new_AGEMA_signal_14597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6776 ( .C (clk), .D (new_AGEMA_signal_14600), .Q (new_AGEMA_signal_14601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6780 ( .C (clk), .D (new_AGEMA_signal_14604), .Q (new_AGEMA_signal_14605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6784 ( .C (clk), .D (new_AGEMA_signal_14608), .Q (new_AGEMA_signal_14609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6788 ( .C (clk), .D (new_AGEMA_signal_14612), .Q (new_AGEMA_signal_14613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6792 ( .C (clk), .D (new_AGEMA_signal_14616), .Q (new_AGEMA_signal_14617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6796 ( .C (clk), .D (new_AGEMA_signal_14620), .Q (new_AGEMA_signal_14621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6800 ( .C (clk), .D (new_AGEMA_signal_14624), .Q (new_AGEMA_signal_14625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6804 ( .C (clk), .D (new_AGEMA_signal_14628), .Q (new_AGEMA_signal_14629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6808 ( .C (clk), .D (new_AGEMA_signal_14632), .Q (new_AGEMA_signal_14633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6812 ( .C (clk), .D (new_AGEMA_signal_14636), .Q (new_AGEMA_signal_14637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6816 ( .C (clk), .D (new_AGEMA_signal_14640), .Q (new_AGEMA_signal_14641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6820 ( .C (clk), .D (new_AGEMA_signal_14644), .Q (new_AGEMA_signal_14645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6824 ( .C (clk), .D (new_AGEMA_signal_14648), .Q (new_AGEMA_signal_14649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6828 ( .C (clk), .D (new_AGEMA_signal_14652), .Q (new_AGEMA_signal_14653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6832 ( .C (clk), .D (new_AGEMA_signal_14656), .Q (new_AGEMA_signal_14657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6836 ( .C (clk), .D (new_AGEMA_signal_14660), .Q (new_AGEMA_signal_14661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6840 ( .C (clk), .D (new_AGEMA_signal_14664), .Q (new_AGEMA_signal_14665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6844 ( .C (clk), .D (new_AGEMA_signal_14668), .Q (new_AGEMA_signal_14669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6848 ( .C (clk), .D (new_AGEMA_signal_14672), .Q (new_AGEMA_signal_14673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6852 ( .C (clk), .D (new_AGEMA_signal_14676), .Q (new_AGEMA_signal_14677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6856 ( .C (clk), .D (new_AGEMA_signal_14680), .Q (new_AGEMA_signal_14681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6860 ( .C (clk), .D (new_AGEMA_signal_14684), .Q (new_AGEMA_signal_14685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6864 ( .C (clk), .D (new_AGEMA_signal_14688), .Q (new_AGEMA_signal_14689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6868 ( .C (clk), .D (new_AGEMA_signal_14692), .Q (new_AGEMA_signal_14693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6872 ( .C (clk), .D (new_AGEMA_signal_14696), .Q (new_AGEMA_signal_14697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6876 ( .C (clk), .D (new_AGEMA_signal_14700), .Q (new_AGEMA_signal_14701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6880 ( .C (clk), .D (new_AGEMA_signal_14704), .Q (new_AGEMA_signal_14705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6884 ( .C (clk), .D (new_AGEMA_signal_14708), .Q (new_AGEMA_signal_14709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6888 ( .C (clk), .D (new_AGEMA_signal_14712), .Q (new_AGEMA_signal_14713) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6892 ( .C (clk), .D (new_AGEMA_signal_14716), .Q (new_AGEMA_signal_14717) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6896 ( .C (clk), .D (new_AGEMA_signal_14720), .Q (new_AGEMA_signal_14721) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6900 ( .C (clk), .D (new_AGEMA_signal_14724), .Q (new_AGEMA_signal_14725) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6904 ( .C (clk), .D (new_AGEMA_signal_14728), .Q (new_AGEMA_signal_14729) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6908 ( .C (clk), .D (new_AGEMA_signal_14732), .Q (new_AGEMA_signal_14733) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6912 ( .C (clk), .D (new_AGEMA_signal_14736), .Q (new_AGEMA_signal_14737) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6916 ( .C (clk), .D (new_AGEMA_signal_14740), .Q (new_AGEMA_signal_14741) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6920 ( .C (clk), .D (new_AGEMA_signal_14744), .Q (new_AGEMA_signal_14745) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6924 ( .C (clk), .D (new_AGEMA_signal_14748), .Q (new_AGEMA_signal_14749) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6928 ( .C (clk), .D (new_AGEMA_signal_14752), .Q (new_AGEMA_signal_14753) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6932 ( .C (clk), .D (new_AGEMA_signal_14756), .Q (new_AGEMA_signal_14757) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6936 ( .C (clk), .D (new_AGEMA_signal_14760), .Q (new_AGEMA_signal_14761) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6940 ( .C (clk), .D (new_AGEMA_signal_14764), .Q (new_AGEMA_signal_14765) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6944 ( .C (clk), .D (new_AGEMA_signal_14768), .Q (new_AGEMA_signal_14769) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6948 ( .C (clk), .D (new_AGEMA_signal_14772), .Q (new_AGEMA_signal_14773) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6952 ( .C (clk), .D (new_AGEMA_signal_14776), .Q (new_AGEMA_signal_14777) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6956 ( .C (clk), .D (new_AGEMA_signal_14780), .Q (new_AGEMA_signal_14781) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6960 ( .C (clk), .D (new_AGEMA_signal_14784), .Q (new_AGEMA_signal_14785) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6964 ( .C (clk), .D (new_AGEMA_signal_14788), .Q (new_AGEMA_signal_14789) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6968 ( .C (clk), .D (new_AGEMA_signal_14792), .Q (new_AGEMA_signal_14793) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6972 ( .C (clk), .D (new_AGEMA_signal_14796), .Q (new_AGEMA_signal_14797) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6976 ( .C (clk), .D (new_AGEMA_signal_14800), .Q (new_AGEMA_signal_14801) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6980 ( .C (clk), .D (new_AGEMA_signal_14804), .Q (new_AGEMA_signal_14805) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6984 ( .C (clk), .D (new_AGEMA_signal_14808), .Q (new_AGEMA_signal_14809) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6988 ( .C (clk), .D (new_AGEMA_signal_14812), .Q (new_AGEMA_signal_14813) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6992 ( .C (clk), .D (new_AGEMA_signal_14816), .Q (new_AGEMA_signal_14817) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6996 ( .C (clk), .D (new_AGEMA_signal_14820), .Q (new_AGEMA_signal_14821) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7000 ( .C (clk), .D (new_AGEMA_signal_14824), .Q (new_AGEMA_signal_14825) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7004 ( .C (clk), .D (new_AGEMA_signal_14828), .Q (new_AGEMA_signal_14829) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7008 ( .C (clk), .D (new_AGEMA_signal_14832), .Q (new_AGEMA_signal_14833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7012 ( .C (clk), .D (new_AGEMA_signal_14836), .Q (new_AGEMA_signal_14837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7016 ( .C (clk), .D (new_AGEMA_signal_14840), .Q (new_AGEMA_signal_14841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7020 ( .C (clk), .D (new_AGEMA_signal_14844), .Q (new_AGEMA_signal_14845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7024 ( .C (clk), .D (new_AGEMA_signal_14848), .Q (new_AGEMA_signal_14849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7028 ( .C (clk), .D (new_AGEMA_signal_14852), .Q (new_AGEMA_signal_14853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7032 ( .C (clk), .D (new_AGEMA_signal_14856), .Q (new_AGEMA_signal_14857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7036 ( .C (clk), .D (new_AGEMA_signal_14860), .Q (new_AGEMA_signal_14861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7040 ( .C (clk), .D (new_AGEMA_signal_14864), .Q (new_AGEMA_signal_14865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7044 ( .C (clk), .D (new_AGEMA_signal_14868), .Q (new_AGEMA_signal_14869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7048 ( .C (clk), .D (new_AGEMA_signal_14872), .Q (new_AGEMA_signal_14873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7052 ( .C (clk), .D (new_AGEMA_signal_14876), .Q (new_AGEMA_signal_14877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7056 ( .C (clk), .D (new_AGEMA_signal_14880), .Q (new_AGEMA_signal_14881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7060 ( .C (clk), .D (new_AGEMA_signal_14884), .Q (new_AGEMA_signal_14885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7064 ( .C (clk), .D (new_AGEMA_signal_14888), .Q (new_AGEMA_signal_14889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7068 ( .C (clk), .D (new_AGEMA_signal_14892), .Q (new_AGEMA_signal_14893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7072 ( .C (clk), .D (new_AGEMA_signal_14896), .Q (new_AGEMA_signal_14897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7076 ( .C (clk), .D (new_AGEMA_signal_14900), .Q (new_AGEMA_signal_14901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7080 ( .C (clk), .D (new_AGEMA_signal_14904), .Q (new_AGEMA_signal_14905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7084 ( .C (clk), .D (new_AGEMA_signal_14908), .Q (new_AGEMA_signal_14909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7088 ( .C (clk), .D (new_AGEMA_signal_14912), .Q (new_AGEMA_signal_14913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7092 ( .C (clk), .D (new_AGEMA_signal_14916), .Q (new_AGEMA_signal_14917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7096 ( .C (clk), .D (new_AGEMA_signal_14920), .Q (new_AGEMA_signal_14921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7100 ( .C (clk), .D (new_AGEMA_signal_14924), .Q (new_AGEMA_signal_14925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7104 ( .C (clk), .D (new_AGEMA_signal_14928), .Q (new_AGEMA_signal_14929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7108 ( .C (clk), .D (new_AGEMA_signal_14932), .Q (new_AGEMA_signal_14933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7112 ( .C (clk), .D (new_AGEMA_signal_14936), .Q (new_AGEMA_signal_14937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7116 ( .C (clk), .D (new_AGEMA_signal_14940), .Q (new_AGEMA_signal_14941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7120 ( .C (clk), .D (new_AGEMA_signal_14944), .Q (new_AGEMA_signal_14945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7124 ( .C (clk), .D (new_AGEMA_signal_14948), .Q (new_AGEMA_signal_14949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7128 ( .C (clk), .D (new_AGEMA_signal_14952), .Q (new_AGEMA_signal_14953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7132 ( .C (clk), .D (new_AGEMA_signal_14956), .Q (new_AGEMA_signal_14957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7136 ( .C (clk), .D (new_AGEMA_signal_14960), .Q (new_AGEMA_signal_14961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7140 ( .C (clk), .D (new_AGEMA_signal_14964), .Q (new_AGEMA_signal_14965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7144 ( .C (clk), .D (new_AGEMA_signal_14968), .Q (new_AGEMA_signal_14969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7148 ( .C (clk), .D (new_AGEMA_signal_14972), .Q (new_AGEMA_signal_14973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7152 ( .C (clk), .D (new_AGEMA_signal_14976), .Q (new_AGEMA_signal_14977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7156 ( .C (clk), .D (new_AGEMA_signal_14980), .Q (new_AGEMA_signal_14981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7160 ( .C (clk), .D (new_AGEMA_signal_14984), .Q (new_AGEMA_signal_14985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7164 ( .C (clk), .D (new_AGEMA_signal_14988), .Q (new_AGEMA_signal_14989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7168 ( .C (clk), .D (new_AGEMA_signal_14992), .Q (new_AGEMA_signal_14993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7172 ( .C (clk), .D (new_AGEMA_signal_14996), .Q (new_AGEMA_signal_14997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7176 ( .C (clk), .D (new_AGEMA_signal_15000), .Q (new_AGEMA_signal_15001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7180 ( .C (clk), .D (new_AGEMA_signal_15004), .Q (new_AGEMA_signal_15005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7184 ( .C (clk), .D (new_AGEMA_signal_15008), .Q (new_AGEMA_signal_15009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7188 ( .C (clk), .D (new_AGEMA_signal_15012), .Q (new_AGEMA_signal_15013) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7192 ( .C (clk), .D (new_AGEMA_signal_15016), .Q (new_AGEMA_signal_15017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7196 ( .C (clk), .D (new_AGEMA_signal_15020), .Q (new_AGEMA_signal_15021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7200 ( .C (clk), .D (new_AGEMA_signal_15024), .Q (new_AGEMA_signal_15025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7204 ( .C (clk), .D (new_AGEMA_signal_15028), .Q (new_AGEMA_signal_15029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7208 ( .C (clk), .D (new_AGEMA_signal_15032), .Q (new_AGEMA_signal_15033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7212 ( .C (clk), .D (new_AGEMA_signal_15036), .Q (new_AGEMA_signal_15037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7216 ( .C (clk), .D (new_AGEMA_signal_15040), .Q (new_AGEMA_signal_15041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7220 ( .C (clk), .D (new_AGEMA_signal_15044), .Q (new_AGEMA_signal_15045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7224 ( .C (clk), .D (new_AGEMA_signal_15048), .Q (new_AGEMA_signal_15049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7228 ( .C (clk), .D (new_AGEMA_signal_15052), .Q (new_AGEMA_signal_15053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7232 ( .C (clk), .D (new_AGEMA_signal_15056), .Q (new_AGEMA_signal_15057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7236 ( .C (clk), .D (new_AGEMA_signal_15060), .Q (new_AGEMA_signal_15061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7240 ( .C (clk), .D (new_AGEMA_signal_15064), .Q (new_AGEMA_signal_15065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7244 ( .C (clk), .D (new_AGEMA_signal_15068), .Q (new_AGEMA_signal_15069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7248 ( .C (clk), .D (new_AGEMA_signal_15072), .Q (new_AGEMA_signal_15073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7252 ( .C (clk), .D (new_AGEMA_signal_15076), .Q (new_AGEMA_signal_15077) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7256 ( .C (clk), .D (new_AGEMA_signal_15080), .Q (new_AGEMA_signal_15081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7260 ( .C (clk), .D (new_AGEMA_signal_15084), .Q (new_AGEMA_signal_15085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7264 ( .C (clk), .D (new_AGEMA_signal_15088), .Q (new_AGEMA_signal_15089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7268 ( .C (clk), .D (new_AGEMA_signal_15092), .Q (new_AGEMA_signal_15093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7272 ( .C (clk), .D (new_AGEMA_signal_15096), .Q (new_AGEMA_signal_15097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7276 ( .C (clk), .D (new_AGEMA_signal_15100), .Q (new_AGEMA_signal_15101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7280 ( .C (clk), .D (new_AGEMA_signal_15104), .Q (new_AGEMA_signal_15105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7284 ( .C (clk), .D (new_AGEMA_signal_15108), .Q (new_AGEMA_signal_15109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7288 ( .C (clk), .D (new_AGEMA_signal_15112), .Q (new_AGEMA_signal_15113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7292 ( .C (clk), .D (new_AGEMA_signal_15116), .Q (new_AGEMA_signal_15117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7296 ( .C (clk), .D (new_AGEMA_signal_15120), .Q (new_AGEMA_signal_15121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7300 ( .C (clk), .D (new_AGEMA_signal_15124), .Q (new_AGEMA_signal_15125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7304 ( .C (clk), .D (new_AGEMA_signal_15128), .Q (new_AGEMA_signal_15129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7308 ( .C (clk), .D (new_AGEMA_signal_15132), .Q (new_AGEMA_signal_15133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7312 ( .C (clk), .D (new_AGEMA_signal_15136), .Q (new_AGEMA_signal_15137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7316 ( .C (clk), .D (new_AGEMA_signal_15140), .Q (new_AGEMA_signal_15141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7320 ( .C (clk), .D (new_AGEMA_signal_15144), .Q (new_AGEMA_signal_15145) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7324 ( .C (clk), .D (new_AGEMA_signal_15148), .Q (new_AGEMA_signal_15149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7328 ( .C (clk), .D (new_AGEMA_signal_15152), .Q (new_AGEMA_signal_15153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7332 ( .C (clk), .D (new_AGEMA_signal_15156), .Q (new_AGEMA_signal_15157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7336 ( .C (clk), .D (new_AGEMA_signal_15160), .Q (new_AGEMA_signal_15161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7340 ( .C (clk), .D (new_AGEMA_signal_15164), .Q (new_AGEMA_signal_15165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7344 ( .C (clk), .D (new_AGEMA_signal_15168), .Q (new_AGEMA_signal_15169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7348 ( .C (clk), .D (new_AGEMA_signal_15172), .Q (new_AGEMA_signal_15173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7352 ( .C (clk), .D (new_AGEMA_signal_15176), .Q (new_AGEMA_signal_15177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7356 ( .C (clk), .D (new_AGEMA_signal_15180), .Q (new_AGEMA_signal_15181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7360 ( .C (clk), .D (new_AGEMA_signal_15184), .Q (new_AGEMA_signal_15185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7364 ( .C (clk), .D (new_AGEMA_signal_15188), .Q (new_AGEMA_signal_15189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7368 ( .C (clk), .D (new_AGEMA_signal_15192), .Q (new_AGEMA_signal_15193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7372 ( .C (clk), .D (new_AGEMA_signal_15196), .Q (new_AGEMA_signal_15197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7376 ( .C (clk), .D (new_AGEMA_signal_15200), .Q (new_AGEMA_signal_15201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7380 ( .C (clk), .D (new_AGEMA_signal_15204), .Q (new_AGEMA_signal_15205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7384 ( .C (clk), .D (new_AGEMA_signal_15208), .Q (new_AGEMA_signal_15209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7388 ( .C (clk), .D (new_AGEMA_signal_15212), .Q (new_AGEMA_signal_15213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7392 ( .C (clk), .D (new_AGEMA_signal_15216), .Q (new_AGEMA_signal_15217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7396 ( .C (clk), .D (new_AGEMA_signal_15220), .Q (new_AGEMA_signal_15221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7400 ( .C (clk), .D (new_AGEMA_signal_15224), .Q (new_AGEMA_signal_15225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7404 ( .C (clk), .D (new_AGEMA_signal_15228), .Q (new_AGEMA_signal_15229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7408 ( .C (clk), .D (new_AGEMA_signal_15232), .Q (new_AGEMA_signal_15233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7412 ( .C (clk), .D (new_AGEMA_signal_15236), .Q (new_AGEMA_signal_15237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7416 ( .C (clk), .D (new_AGEMA_signal_15240), .Q (new_AGEMA_signal_15241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7420 ( .C (clk), .D (new_AGEMA_signal_15244), .Q (new_AGEMA_signal_15245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7424 ( .C (clk), .D (new_AGEMA_signal_15248), .Q (new_AGEMA_signal_15249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7428 ( .C (clk), .D (new_AGEMA_signal_15252), .Q (new_AGEMA_signal_15253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7432 ( .C (clk), .D (new_AGEMA_signal_15256), .Q (new_AGEMA_signal_15257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7436 ( .C (clk), .D (new_AGEMA_signal_15260), .Q (new_AGEMA_signal_15261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7440 ( .C (clk), .D (new_AGEMA_signal_15264), .Q (new_AGEMA_signal_15265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7444 ( .C (clk), .D (new_AGEMA_signal_15268), .Q (new_AGEMA_signal_15269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7448 ( .C (clk), .D (new_AGEMA_signal_15272), .Q (new_AGEMA_signal_15273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7452 ( .C (clk), .D (new_AGEMA_signal_15276), .Q (new_AGEMA_signal_15277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7456 ( .C (clk), .D (new_AGEMA_signal_15280), .Q (new_AGEMA_signal_15281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7460 ( .C (clk), .D (new_AGEMA_signal_15284), .Q (new_AGEMA_signal_15285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7464 ( .C (clk), .D (new_AGEMA_signal_15288), .Q (new_AGEMA_signal_15289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7468 ( .C (clk), .D (new_AGEMA_signal_15292), .Q (new_AGEMA_signal_15293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7472 ( .C (clk), .D (new_AGEMA_signal_15296), .Q (new_AGEMA_signal_15297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7476 ( .C (clk), .D (new_AGEMA_signal_15300), .Q (new_AGEMA_signal_15301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7480 ( .C (clk), .D (new_AGEMA_signal_15304), .Q (new_AGEMA_signal_15305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7484 ( .C (clk), .D (new_AGEMA_signal_15308), .Q (new_AGEMA_signal_15309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7488 ( .C (clk), .D (new_AGEMA_signal_15312), .Q (new_AGEMA_signal_15313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7492 ( .C (clk), .D (new_AGEMA_signal_15316), .Q (new_AGEMA_signal_15317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7496 ( .C (clk), .D (new_AGEMA_signal_15320), .Q (new_AGEMA_signal_15321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7500 ( .C (clk), .D (new_AGEMA_signal_15324), .Q (new_AGEMA_signal_15325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7504 ( .C (clk), .D (new_AGEMA_signal_15328), .Q (new_AGEMA_signal_15329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7508 ( .C (clk), .D (new_AGEMA_signal_15332), .Q (new_AGEMA_signal_15333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7512 ( .C (clk), .D (new_AGEMA_signal_15336), .Q (new_AGEMA_signal_15337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7516 ( .C (clk), .D (new_AGEMA_signal_15340), .Q (new_AGEMA_signal_15341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7520 ( .C (clk), .D (new_AGEMA_signal_15344), .Q (new_AGEMA_signal_15345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7524 ( .C (clk), .D (new_AGEMA_signal_15348), .Q (new_AGEMA_signal_15349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7528 ( .C (clk), .D (new_AGEMA_signal_15352), .Q (new_AGEMA_signal_15353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7532 ( .C (clk), .D (new_AGEMA_signal_15356), .Q (new_AGEMA_signal_15357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7536 ( .C (clk), .D (new_AGEMA_signal_15360), .Q (new_AGEMA_signal_15361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7540 ( .C (clk), .D (new_AGEMA_signal_15364), .Q (new_AGEMA_signal_15365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7544 ( .C (clk), .D (new_AGEMA_signal_15368), .Q (new_AGEMA_signal_15369) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7548 ( .C (clk), .D (new_AGEMA_signal_15372), .Q (new_AGEMA_signal_15373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7552 ( .C (clk), .D (new_AGEMA_signal_15376), .Q (new_AGEMA_signal_15377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7556 ( .C (clk), .D (new_AGEMA_signal_15380), .Q (new_AGEMA_signal_15381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7560 ( .C (clk), .D (new_AGEMA_signal_15384), .Q (new_AGEMA_signal_15385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7564 ( .C (clk), .D (new_AGEMA_signal_15388), .Q (new_AGEMA_signal_15389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7568 ( .C (clk), .D (new_AGEMA_signal_15392), .Q (new_AGEMA_signal_15393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7572 ( .C (clk), .D (new_AGEMA_signal_15396), .Q (new_AGEMA_signal_15397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7576 ( .C (clk), .D (new_AGEMA_signal_15400), .Q (new_AGEMA_signal_15401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7580 ( .C (clk), .D (new_AGEMA_signal_15404), .Q (new_AGEMA_signal_15405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7584 ( .C (clk), .D (new_AGEMA_signal_15408), .Q (new_AGEMA_signal_15409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7588 ( .C (clk), .D (new_AGEMA_signal_15412), .Q (new_AGEMA_signal_15413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7592 ( .C (clk), .D (new_AGEMA_signal_15416), .Q (new_AGEMA_signal_15417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7596 ( .C (clk), .D (new_AGEMA_signal_15420), .Q (new_AGEMA_signal_15421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7600 ( .C (clk), .D (new_AGEMA_signal_15424), .Q (new_AGEMA_signal_15425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7604 ( .C (clk), .D (new_AGEMA_signal_15428), .Q (new_AGEMA_signal_15429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7608 ( .C (clk), .D (new_AGEMA_signal_15432), .Q (new_AGEMA_signal_15433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7612 ( .C (clk), .D (new_AGEMA_signal_15436), .Q (new_AGEMA_signal_15437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7616 ( .C (clk), .D (new_AGEMA_signal_15440), .Q (new_AGEMA_signal_15441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7620 ( .C (clk), .D (new_AGEMA_signal_15444), .Q (new_AGEMA_signal_15445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7624 ( .C (clk), .D (new_AGEMA_signal_15448), .Q (new_AGEMA_signal_15449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7628 ( .C (clk), .D (new_AGEMA_signal_15452), .Q (new_AGEMA_signal_15453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7632 ( .C (clk), .D (new_AGEMA_signal_15456), .Q (new_AGEMA_signal_15457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7636 ( .C (clk), .D (new_AGEMA_signal_15460), .Q (new_AGEMA_signal_15461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7640 ( .C (clk), .D (new_AGEMA_signal_15464), .Q (new_AGEMA_signal_15465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7644 ( .C (clk), .D (new_AGEMA_signal_15468), .Q (new_AGEMA_signal_15469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7648 ( .C (clk), .D (new_AGEMA_signal_15472), .Q (new_AGEMA_signal_15473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7652 ( .C (clk), .D (new_AGEMA_signal_15476), .Q (new_AGEMA_signal_15477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7656 ( .C (clk), .D (new_AGEMA_signal_15480), .Q (new_AGEMA_signal_15481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7660 ( .C (clk), .D (new_AGEMA_signal_15484), .Q (new_AGEMA_signal_15485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7664 ( .C (clk), .D (new_AGEMA_signal_15488), .Q (new_AGEMA_signal_15489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7668 ( .C (clk), .D (new_AGEMA_signal_15492), .Q (new_AGEMA_signal_15493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7672 ( .C (clk), .D (new_AGEMA_signal_15496), .Q (new_AGEMA_signal_15497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7676 ( .C (clk), .D (new_AGEMA_signal_15500), .Q (new_AGEMA_signal_15501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7680 ( .C (clk), .D (new_AGEMA_signal_15504), .Q (new_AGEMA_signal_15505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7684 ( .C (clk), .D (new_AGEMA_signal_15508), .Q (new_AGEMA_signal_15509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7688 ( .C (clk), .D (new_AGEMA_signal_15512), .Q (new_AGEMA_signal_15513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7692 ( .C (clk), .D (new_AGEMA_signal_15516), .Q (new_AGEMA_signal_15517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7696 ( .C (clk), .D (new_AGEMA_signal_15520), .Q (new_AGEMA_signal_15521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7700 ( .C (clk), .D (new_AGEMA_signal_15524), .Q (new_AGEMA_signal_15525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7704 ( .C (clk), .D (new_AGEMA_signal_15528), .Q (new_AGEMA_signal_15529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7708 ( .C (clk), .D (new_AGEMA_signal_15532), .Q (new_AGEMA_signal_15533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7712 ( .C (clk), .D (new_AGEMA_signal_15536), .Q (new_AGEMA_signal_15537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7716 ( .C (clk), .D (new_AGEMA_signal_15540), .Q (new_AGEMA_signal_15541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7720 ( .C (clk), .D (new_AGEMA_signal_15544), .Q (new_AGEMA_signal_15545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7724 ( .C (clk), .D (new_AGEMA_signal_15548), .Q (new_AGEMA_signal_15549) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7728 ( .C (clk), .D (new_AGEMA_signal_15552), .Q (new_AGEMA_signal_15553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7732 ( .C (clk), .D (new_AGEMA_signal_15556), .Q (new_AGEMA_signal_15557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7736 ( .C (clk), .D (new_AGEMA_signal_15560), .Q (new_AGEMA_signal_15561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7740 ( .C (clk), .D (new_AGEMA_signal_15564), .Q (new_AGEMA_signal_15565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7744 ( .C (clk), .D (new_AGEMA_signal_15568), .Q (new_AGEMA_signal_15569) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7748 ( .C (clk), .D (new_AGEMA_signal_15572), .Q (new_AGEMA_signal_15573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7752 ( .C (clk), .D (new_AGEMA_signal_15576), .Q (new_AGEMA_signal_15577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7756 ( .C (clk), .D (new_AGEMA_signal_15580), .Q (new_AGEMA_signal_15581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7760 ( .C (clk), .D (new_AGEMA_signal_15584), .Q (new_AGEMA_signal_15585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7764 ( .C (clk), .D (new_AGEMA_signal_15588), .Q (new_AGEMA_signal_15589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7768 ( .C (clk), .D (new_AGEMA_signal_15592), .Q (new_AGEMA_signal_15593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7772 ( .C (clk), .D (new_AGEMA_signal_15596), .Q (new_AGEMA_signal_15597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7776 ( .C (clk), .D (new_AGEMA_signal_15600), .Q (new_AGEMA_signal_15601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7780 ( .C (clk), .D (new_AGEMA_signal_15604), .Q (new_AGEMA_signal_15605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7784 ( .C (clk), .D (new_AGEMA_signal_15608), .Q (new_AGEMA_signal_15609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7788 ( .C (clk), .D (new_AGEMA_signal_15612), .Q (new_AGEMA_signal_15613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7792 ( .C (clk), .D (new_AGEMA_signal_15616), .Q (new_AGEMA_signal_15617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7796 ( .C (clk), .D (new_AGEMA_signal_15620), .Q (new_AGEMA_signal_15621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7800 ( .C (clk), .D (new_AGEMA_signal_15624), .Q (new_AGEMA_signal_15625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7804 ( .C (clk), .D (new_AGEMA_signal_15628), .Q (new_AGEMA_signal_15629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7808 ( .C (clk), .D (new_AGEMA_signal_15632), .Q (new_AGEMA_signal_15633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7812 ( .C (clk), .D (new_AGEMA_signal_15636), .Q (new_AGEMA_signal_15637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7816 ( .C (clk), .D (new_AGEMA_signal_15640), .Q (new_AGEMA_signal_15641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7820 ( .C (clk), .D (new_AGEMA_signal_15644), .Q (new_AGEMA_signal_15645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7824 ( .C (clk), .D (new_AGEMA_signal_15648), .Q (new_AGEMA_signal_15649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7828 ( .C (clk), .D (new_AGEMA_signal_15652), .Q (new_AGEMA_signal_15653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7832 ( .C (clk), .D (new_AGEMA_signal_15656), .Q (new_AGEMA_signal_15657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7836 ( .C (clk), .D (new_AGEMA_signal_15660), .Q (new_AGEMA_signal_15661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7840 ( .C (clk), .D (new_AGEMA_signal_15664), .Q (new_AGEMA_signal_15665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7844 ( .C (clk), .D (new_AGEMA_signal_15668), .Q (new_AGEMA_signal_15669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7848 ( .C (clk), .D (new_AGEMA_signal_15672), .Q (new_AGEMA_signal_15673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7852 ( .C (clk), .D (new_AGEMA_signal_15676), .Q (new_AGEMA_signal_15677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7856 ( .C (clk), .D (new_AGEMA_signal_15680), .Q (new_AGEMA_signal_15681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7860 ( .C (clk), .D (new_AGEMA_signal_15684), .Q (new_AGEMA_signal_15685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7864 ( .C (clk), .D (new_AGEMA_signal_15688), .Q (new_AGEMA_signal_15689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7868 ( .C (clk), .D (new_AGEMA_signal_15692), .Q (new_AGEMA_signal_15693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7872 ( .C (clk), .D (new_AGEMA_signal_15696), .Q (new_AGEMA_signal_15697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7876 ( .C (clk), .D (new_AGEMA_signal_15700), .Q (new_AGEMA_signal_15701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7880 ( .C (clk), .D (new_AGEMA_signal_15704), .Q (new_AGEMA_signal_15705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7884 ( .C (clk), .D (new_AGEMA_signal_15708), .Q (new_AGEMA_signal_15709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7888 ( .C (clk), .D (new_AGEMA_signal_15712), .Q (new_AGEMA_signal_15713) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7892 ( .C (clk), .D (new_AGEMA_signal_15716), .Q (new_AGEMA_signal_15717) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7896 ( .C (clk), .D (new_AGEMA_signal_15720), .Q (new_AGEMA_signal_15721) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7900 ( .C (clk), .D (new_AGEMA_signal_15724), .Q (new_AGEMA_signal_15725) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7904 ( .C (clk), .D (new_AGEMA_signal_15728), .Q (new_AGEMA_signal_15729) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7908 ( .C (clk), .D (new_AGEMA_signal_15732), .Q (new_AGEMA_signal_15733) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7912 ( .C (clk), .D (new_AGEMA_signal_15736), .Q (new_AGEMA_signal_15737) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7916 ( .C (clk), .D (new_AGEMA_signal_15740), .Q (new_AGEMA_signal_15741) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7920 ( .C (clk), .D (new_AGEMA_signal_15744), .Q (new_AGEMA_signal_15745) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7924 ( .C (clk), .D (new_AGEMA_signal_15748), .Q (new_AGEMA_signal_15749) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7928 ( .C (clk), .D (new_AGEMA_signal_15752), .Q (new_AGEMA_signal_15753) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7932 ( .C (clk), .D (new_AGEMA_signal_15756), .Q (new_AGEMA_signal_15757) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7936 ( .C (clk), .D (new_AGEMA_signal_15760), .Q (new_AGEMA_signal_15761) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7940 ( .C (clk), .D (new_AGEMA_signal_15764), .Q (new_AGEMA_signal_15765) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7944 ( .C (clk), .D (new_AGEMA_signal_15768), .Q (new_AGEMA_signal_15769) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7948 ( .C (clk), .D (new_AGEMA_signal_15772), .Q (new_AGEMA_signal_15773) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7952 ( .C (clk), .D (new_AGEMA_signal_15776), .Q (new_AGEMA_signal_15777) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7956 ( .C (clk), .D (new_AGEMA_signal_15780), .Q (new_AGEMA_signal_15781) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7960 ( .C (clk), .D (new_AGEMA_signal_15784), .Q (new_AGEMA_signal_15785) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7964 ( .C (clk), .D (new_AGEMA_signal_15788), .Q (new_AGEMA_signal_15789) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7968 ( .C (clk), .D (new_AGEMA_signal_15792), .Q (new_AGEMA_signal_15793) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7972 ( .C (clk), .D (new_AGEMA_signal_15796), .Q (new_AGEMA_signal_15797) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7976 ( .C (clk), .D (new_AGEMA_signal_15800), .Q (new_AGEMA_signal_15801) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7980 ( .C (clk), .D (new_AGEMA_signal_15804), .Q (new_AGEMA_signal_15805) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7984 ( .C (clk), .D (new_AGEMA_signal_15808), .Q (new_AGEMA_signal_15809) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7988 ( .C (clk), .D (new_AGEMA_signal_15812), .Q (new_AGEMA_signal_15813) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7992 ( .C (clk), .D (new_AGEMA_signal_15816), .Q (new_AGEMA_signal_15817) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7996 ( .C (clk), .D (new_AGEMA_signal_15820), .Q (new_AGEMA_signal_15821) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8000 ( .C (clk), .D (new_AGEMA_signal_15824), .Q (new_AGEMA_signal_15825) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8004 ( .C (clk), .D (new_AGEMA_signal_15828), .Q (new_AGEMA_signal_15829) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8008 ( .C (clk), .D (new_AGEMA_signal_15832), .Q (new_AGEMA_signal_15833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8012 ( .C (clk), .D (new_AGEMA_signal_15836), .Q (new_AGEMA_signal_15837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8016 ( .C (clk), .D (new_AGEMA_signal_15840), .Q (new_AGEMA_signal_15841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8020 ( .C (clk), .D (new_AGEMA_signal_15844), .Q (new_AGEMA_signal_15845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8024 ( .C (clk), .D (new_AGEMA_signal_15848), .Q (new_AGEMA_signal_15849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8028 ( .C (clk), .D (new_AGEMA_signal_15852), .Q (new_AGEMA_signal_15853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8032 ( .C (clk), .D (new_AGEMA_signal_15856), .Q (new_AGEMA_signal_15857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8036 ( .C (clk), .D (new_AGEMA_signal_15860), .Q (new_AGEMA_signal_15861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8040 ( .C (clk), .D (new_AGEMA_signal_15864), .Q (new_AGEMA_signal_15865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8044 ( .C (clk), .D (new_AGEMA_signal_15868), .Q (new_AGEMA_signal_15869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8048 ( .C (clk), .D (new_AGEMA_signal_15872), .Q (new_AGEMA_signal_15873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8052 ( .C (clk), .D (new_AGEMA_signal_15876), .Q (new_AGEMA_signal_15877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8056 ( .C (clk), .D (new_AGEMA_signal_15880), .Q (new_AGEMA_signal_15881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8060 ( .C (clk), .D (new_AGEMA_signal_15884), .Q (new_AGEMA_signal_15885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8064 ( .C (clk), .D (new_AGEMA_signal_15888), .Q (new_AGEMA_signal_15889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8068 ( .C (clk), .D (new_AGEMA_signal_15892), .Q (new_AGEMA_signal_15893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8072 ( .C (clk), .D (new_AGEMA_signal_15896), .Q (new_AGEMA_signal_15897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8076 ( .C (clk), .D (new_AGEMA_signal_15900), .Q (new_AGEMA_signal_15901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8080 ( .C (clk), .D (new_AGEMA_signal_15904), .Q (new_AGEMA_signal_15905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8084 ( .C (clk), .D (new_AGEMA_signal_15908), .Q (new_AGEMA_signal_15909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8088 ( .C (clk), .D (new_AGEMA_signal_15912), .Q (new_AGEMA_signal_15913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8092 ( .C (clk), .D (new_AGEMA_signal_15916), .Q (new_AGEMA_signal_15917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8096 ( .C (clk), .D (new_AGEMA_signal_15920), .Q (new_AGEMA_signal_15921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8100 ( .C (clk), .D (new_AGEMA_signal_15924), .Q (new_AGEMA_signal_15925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8104 ( .C (clk), .D (new_AGEMA_signal_15928), .Q (new_AGEMA_signal_15929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8108 ( .C (clk), .D (new_AGEMA_signal_15932), .Q (new_AGEMA_signal_15933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8112 ( .C (clk), .D (new_AGEMA_signal_15936), .Q (new_AGEMA_signal_15937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8116 ( .C (clk), .D (new_AGEMA_signal_15940), .Q (new_AGEMA_signal_15941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8120 ( .C (clk), .D (new_AGEMA_signal_15944), .Q (new_AGEMA_signal_15945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8124 ( .C (clk), .D (new_AGEMA_signal_15948), .Q (new_AGEMA_signal_15949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8128 ( .C (clk), .D (new_AGEMA_signal_15952), .Q (new_AGEMA_signal_15953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8132 ( .C (clk), .D (new_AGEMA_signal_15956), .Q (new_AGEMA_signal_15957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8136 ( .C (clk), .D (new_AGEMA_signal_15960), .Q (new_AGEMA_signal_15961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8140 ( .C (clk), .D (new_AGEMA_signal_15964), .Q (new_AGEMA_signal_15965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8144 ( .C (clk), .D (new_AGEMA_signal_15968), .Q (new_AGEMA_signal_15969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8148 ( .C (clk), .D (new_AGEMA_signal_15972), .Q (new_AGEMA_signal_15973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8152 ( .C (clk), .D (new_AGEMA_signal_15976), .Q (new_AGEMA_signal_15977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8156 ( .C (clk), .D (new_AGEMA_signal_15980), .Q (new_AGEMA_signal_15981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8160 ( .C (clk), .D (new_AGEMA_signal_15984), .Q (new_AGEMA_signal_15985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8164 ( .C (clk), .D (new_AGEMA_signal_15988), .Q (new_AGEMA_signal_15989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8168 ( .C (clk), .D (new_AGEMA_signal_15992), .Q (new_AGEMA_signal_15993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8172 ( .C (clk), .D (new_AGEMA_signal_15996), .Q (new_AGEMA_signal_15997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8176 ( .C (clk), .D (new_AGEMA_signal_16000), .Q (new_AGEMA_signal_16001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8180 ( .C (clk), .D (new_AGEMA_signal_16004), .Q (new_AGEMA_signal_16005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8184 ( .C (clk), .D (new_AGEMA_signal_16008), .Q (new_AGEMA_signal_16009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8188 ( .C (clk), .D (new_AGEMA_signal_16012), .Q (new_AGEMA_signal_16013) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8192 ( .C (clk), .D (new_AGEMA_signal_16016), .Q (new_AGEMA_signal_16017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8196 ( .C (clk), .D (new_AGEMA_signal_16020), .Q (new_AGEMA_signal_16021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8200 ( .C (clk), .D (new_AGEMA_signal_16024), .Q (new_AGEMA_signal_16025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8204 ( .C (clk), .D (new_AGEMA_signal_16028), .Q (new_AGEMA_signal_16029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8208 ( .C (clk), .D (new_AGEMA_signal_16032), .Q (new_AGEMA_signal_16033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8212 ( .C (clk), .D (new_AGEMA_signal_16036), .Q (new_AGEMA_signal_16037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8216 ( .C (clk), .D (new_AGEMA_signal_16040), .Q (new_AGEMA_signal_16041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8220 ( .C (clk), .D (new_AGEMA_signal_16044), .Q (new_AGEMA_signal_16045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8224 ( .C (clk), .D (new_AGEMA_signal_16048), .Q (new_AGEMA_signal_16049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8228 ( .C (clk), .D (new_AGEMA_signal_16052), .Q (new_AGEMA_signal_16053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8232 ( .C (clk), .D (new_AGEMA_signal_16056), .Q (new_AGEMA_signal_16057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8236 ( .C (clk), .D (new_AGEMA_signal_16060), .Q (new_AGEMA_signal_16061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8240 ( .C (clk), .D (new_AGEMA_signal_16064), .Q (new_AGEMA_signal_16065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8244 ( .C (clk), .D (new_AGEMA_signal_16068), .Q (new_AGEMA_signal_16069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8248 ( .C (clk), .D (new_AGEMA_signal_16072), .Q (new_AGEMA_signal_16073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8252 ( .C (clk), .D (new_AGEMA_signal_16076), .Q (new_AGEMA_signal_16077) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8256 ( .C (clk), .D (new_AGEMA_signal_16080), .Q (new_AGEMA_signal_16081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8260 ( .C (clk), .D (new_AGEMA_signal_16084), .Q (new_AGEMA_signal_16085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8264 ( .C (clk), .D (new_AGEMA_signal_16088), .Q (new_AGEMA_signal_16089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8268 ( .C (clk), .D (new_AGEMA_signal_16092), .Q (new_AGEMA_signal_16093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8272 ( .C (clk), .D (new_AGEMA_signal_16096), .Q (new_AGEMA_signal_16097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8276 ( .C (clk), .D (new_AGEMA_signal_16100), .Q (new_AGEMA_signal_16101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8280 ( .C (clk), .D (new_AGEMA_signal_16104), .Q (new_AGEMA_signal_16105) ) ;
    buf_clk new_AGEMA_reg_buffer_8284 ( .C (clk), .D (new_AGEMA_signal_16108), .Q (new_AGEMA_signal_16109) ) ;
    buf_clk new_AGEMA_reg_buffer_8288 ( .C (clk), .D (new_AGEMA_signal_16112), .Q (new_AGEMA_signal_16113) ) ;
    buf_clk new_AGEMA_reg_buffer_8292 ( .C (clk), .D (new_AGEMA_signal_16116), .Q (new_AGEMA_signal_16117) ) ;
    buf_clk new_AGEMA_reg_buffer_8296 ( .C (clk), .D (new_AGEMA_signal_16120), .Q (new_AGEMA_signal_16121) ) ;
    buf_clk new_AGEMA_reg_buffer_8300 ( .C (clk), .D (new_AGEMA_signal_16124), .Q (new_AGEMA_signal_16125) ) ;
    buf_clk new_AGEMA_reg_buffer_8304 ( .C (clk), .D (new_AGEMA_signal_16128), .Q (new_AGEMA_signal_16129) ) ;
    buf_clk new_AGEMA_reg_buffer_8308 ( .C (clk), .D (new_AGEMA_signal_16132), .Q (new_AGEMA_signal_16133) ) ;
    buf_clk new_AGEMA_reg_buffer_8312 ( .C (clk), .D (new_AGEMA_signal_16136), .Q (new_AGEMA_signal_16137) ) ;
    buf_clk new_AGEMA_reg_buffer_8316 ( .C (clk), .D (new_AGEMA_signal_16140), .Q (new_AGEMA_signal_16141) ) ;
    buf_clk new_AGEMA_reg_buffer_8320 ( .C (clk), .D (new_AGEMA_signal_16144), .Q (new_AGEMA_signal_16145) ) ;
    buf_clk new_AGEMA_reg_buffer_8324 ( .C (clk), .D (new_AGEMA_signal_16148), .Q (new_AGEMA_signal_16149) ) ;
    buf_clk new_AGEMA_reg_buffer_8328 ( .C (clk), .D (new_AGEMA_signal_16152), .Q (new_AGEMA_signal_16153) ) ;
    buf_clk new_AGEMA_reg_buffer_8332 ( .C (clk), .D (new_AGEMA_signal_16156), .Q (new_AGEMA_signal_16157) ) ;
    buf_clk new_AGEMA_reg_buffer_8336 ( .C (clk), .D (new_AGEMA_signal_16160), .Q (new_AGEMA_signal_16161) ) ;
    buf_clk new_AGEMA_reg_buffer_8340 ( .C (clk), .D (new_AGEMA_signal_16164), .Q (new_AGEMA_signal_16165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8344 ( .C (clk), .D (new_AGEMA_signal_16168), .Q (new_AGEMA_signal_16169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8348 ( .C (clk), .D (new_AGEMA_signal_16172), .Q (new_AGEMA_signal_16173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8352 ( .C (clk), .D (new_AGEMA_signal_16176), .Q (new_AGEMA_signal_16177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8356 ( .C (clk), .D (new_AGEMA_signal_16180), .Q (new_AGEMA_signal_16181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8360 ( .C (clk), .D (new_AGEMA_signal_16184), .Q (new_AGEMA_signal_16185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8364 ( .C (clk), .D (new_AGEMA_signal_16188), .Q (new_AGEMA_signal_16189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8368 ( .C (clk), .D (new_AGEMA_signal_16192), .Q (new_AGEMA_signal_16193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8372 ( .C (clk), .D (new_AGEMA_signal_16196), .Q (new_AGEMA_signal_16197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8376 ( .C (clk), .D (new_AGEMA_signal_16200), .Q (new_AGEMA_signal_16201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8380 ( .C (clk), .D (new_AGEMA_signal_16204), .Q (new_AGEMA_signal_16205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8384 ( .C (clk), .D (new_AGEMA_signal_16208), .Q (new_AGEMA_signal_16209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8388 ( .C (clk), .D (new_AGEMA_signal_16212), .Q (new_AGEMA_signal_16213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8392 ( .C (clk), .D (new_AGEMA_signal_16216), .Q (new_AGEMA_signal_16217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8396 ( .C (clk), .D (new_AGEMA_signal_16220), .Q (new_AGEMA_signal_16221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8400 ( .C (clk), .D (new_AGEMA_signal_16224), .Q (new_AGEMA_signal_16225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8404 ( .C (clk), .D (new_AGEMA_signal_16228), .Q (new_AGEMA_signal_16229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8408 ( .C (clk), .D (new_AGEMA_signal_16232), .Q (new_AGEMA_signal_16233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8412 ( .C (clk), .D (new_AGEMA_signal_16236), .Q (new_AGEMA_signal_16237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8416 ( .C (clk), .D (new_AGEMA_signal_16240), .Q (new_AGEMA_signal_16241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8420 ( .C (clk), .D (new_AGEMA_signal_16244), .Q (new_AGEMA_signal_16245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8424 ( .C (clk), .D (new_AGEMA_signal_16248), .Q (new_AGEMA_signal_16249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8428 ( .C (clk), .D (new_AGEMA_signal_16252), .Q (new_AGEMA_signal_16253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8432 ( .C (clk), .D (new_AGEMA_signal_16256), .Q (new_AGEMA_signal_16257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8436 ( .C (clk), .D (new_AGEMA_signal_16260), .Q (new_AGEMA_signal_16261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8440 ( .C (clk), .D (new_AGEMA_signal_16264), .Q (new_AGEMA_signal_16265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8444 ( .C (clk), .D (new_AGEMA_signal_16268), .Q (new_AGEMA_signal_16269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8448 ( .C (clk), .D (new_AGEMA_signal_16272), .Q (new_AGEMA_signal_16273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8452 ( .C (clk), .D (new_AGEMA_signal_16276), .Q (new_AGEMA_signal_16277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8456 ( .C (clk), .D (new_AGEMA_signal_16280), .Q (new_AGEMA_signal_16281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8460 ( .C (clk), .D (new_AGEMA_signal_16284), .Q (new_AGEMA_signal_16285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8464 ( .C (clk), .D (new_AGEMA_signal_16288), .Q (new_AGEMA_signal_16289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8468 ( .C (clk), .D (new_AGEMA_signal_16292), .Q (new_AGEMA_signal_16293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8472 ( .C (clk), .D (new_AGEMA_signal_16296), .Q (new_AGEMA_signal_16297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8476 ( .C (clk), .D (new_AGEMA_signal_16300), .Q (new_AGEMA_signal_16301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8480 ( .C (clk), .D (new_AGEMA_signal_16304), .Q (new_AGEMA_signal_16305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8484 ( .C (clk), .D (new_AGEMA_signal_16308), .Q (new_AGEMA_signal_16309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8488 ( .C (clk), .D (new_AGEMA_signal_16312), .Q (new_AGEMA_signal_16313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8492 ( .C (clk), .D (new_AGEMA_signal_16316), .Q (new_AGEMA_signal_16317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8496 ( .C (clk), .D (new_AGEMA_signal_16320), .Q (new_AGEMA_signal_16321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8500 ( .C (clk), .D (new_AGEMA_signal_16324), .Q (new_AGEMA_signal_16325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8504 ( .C (clk), .D (new_AGEMA_signal_16328), .Q (new_AGEMA_signal_16329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8508 ( .C (clk), .D (new_AGEMA_signal_16332), .Q (new_AGEMA_signal_16333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8512 ( .C (clk), .D (new_AGEMA_signal_16336), .Q (new_AGEMA_signal_16337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8516 ( .C (clk), .D (new_AGEMA_signal_16340), .Q (new_AGEMA_signal_16341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8520 ( .C (clk), .D (new_AGEMA_signal_16344), .Q (new_AGEMA_signal_16345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8524 ( .C (clk), .D (new_AGEMA_signal_16348), .Q (new_AGEMA_signal_16349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8528 ( .C (clk), .D (new_AGEMA_signal_16352), .Q (new_AGEMA_signal_16353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8532 ( .C (clk), .D (new_AGEMA_signal_16356), .Q (new_AGEMA_signal_16357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8536 ( .C (clk), .D (new_AGEMA_signal_16360), .Q (new_AGEMA_signal_16361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8540 ( .C (clk), .D (new_AGEMA_signal_16364), .Q (new_AGEMA_signal_16365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8544 ( .C (clk), .D (new_AGEMA_signal_16368), .Q (new_AGEMA_signal_16369) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8548 ( .C (clk), .D (new_AGEMA_signal_16372), .Q (new_AGEMA_signal_16373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8552 ( .C (clk), .D (new_AGEMA_signal_16376), .Q (new_AGEMA_signal_16377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8556 ( .C (clk), .D (new_AGEMA_signal_16380), .Q (new_AGEMA_signal_16381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8560 ( .C (clk), .D (new_AGEMA_signal_16384), .Q (new_AGEMA_signal_16385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8564 ( .C (clk), .D (new_AGEMA_signal_16388), .Q (new_AGEMA_signal_16389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8568 ( .C (clk), .D (new_AGEMA_signal_16392), .Q (new_AGEMA_signal_16393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8572 ( .C (clk), .D (new_AGEMA_signal_16396), .Q (new_AGEMA_signal_16397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8576 ( .C (clk), .D (new_AGEMA_signal_16400), .Q (new_AGEMA_signal_16401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8580 ( .C (clk), .D (new_AGEMA_signal_16404), .Q (new_AGEMA_signal_16405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8584 ( .C (clk), .D (new_AGEMA_signal_16408), .Q (new_AGEMA_signal_16409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8588 ( .C (clk), .D (new_AGEMA_signal_16412), .Q (new_AGEMA_signal_16413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8592 ( .C (clk), .D (new_AGEMA_signal_16416), .Q (new_AGEMA_signal_16417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8596 ( .C (clk), .D (new_AGEMA_signal_16420), .Q (new_AGEMA_signal_16421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8600 ( .C (clk), .D (new_AGEMA_signal_16424), .Q (new_AGEMA_signal_16425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8604 ( .C (clk), .D (new_AGEMA_signal_16428), .Q (new_AGEMA_signal_16429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8608 ( .C (clk), .D (new_AGEMA_signal_16432), .Q (new_AGEMA_signal_16433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8612 ( .C (clk), .D (new_AGEMA_signal_16436), .Q (new_AGEMA_signal_16437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8616 ( .C (clk), .D (new_AGEMA_signal_16440), .Q (new_AGEMA_signal_16441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8620 ( .C (clk), .D (new_AGEMA_signal_16444), .Q (new_AGEMA_signal_16445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8624 ( .C (clk), .D (new_AGEMA_signal_16448), .Q (new_AGEMA_signal_16449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8628 ( .C (clk), .D (new_AGEMA_signal_16452), .Q (new_AGEMA_signal_16453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8632 ( .C (clk), .D (new_AGEMA_signal_16456), .Q (new_AGEMA_signal_16457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8636 ( .C (clk), .D (new_AGEMA_signal_16460), .Q (new_AGEMA_signal_16461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8640 ( .C (clk), .D (new_AGEMA_signal_16464), .Q (new_AGEMA_signal_16465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8644 ( .C (clk), .D (new_AGEMA_signal_16468), .Q (new_AGEMA_signal_16469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8648 ( .C (clk), .D (new_AGEMA_signal_16472), .Q (new_AGEMA_signal_16473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8652 ( .C (clk), .D (new_AGEMA_signal_16476), .Q (new_AGEMA_signal_16477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8656 ( .C (clk), .D (new_AGEMA_signal_16480), .Q (new_AGEMA_signal_16481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8660 ( .C (clk), .D (new_AGEMA_signal_16484), .Q (new_AGEMA_signal_16485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8664 ( .C (clk), .D (new_AGEMA_signal_16488), .Q (new_AGEMA_signal_16489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8668 ( .C (clk), .D (new_AGEMA_signal_16492), .Q (new_AGEMA_signal_16493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8672 ( .C (clk), .D (new_AGEMA_signal_16496), .Q (new_AGEMA_signal_16497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8676 ( .C (clk), .D (new_AGEMA_signal_16500), .Q (new_AGEMA_signal_16501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8680 ( .C (clk), .D (new_AGEMA_signal_16504), .Q (new_AGEMA_signal_16505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8684 ( .C (clk), .D (new_AGEMA_signal_16508), .Q (new_AGEMA_signal_16509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8688 ( .C (clk), .D (new_AGEMA_signal_16512), .Q (new_AGEMA_signal_16513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8692 ( .C (clk), .D (new_AGEMA_signal_16516), .Q (new_AGEMA_signal_16517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8696 ( .C (clk), .D (new_AGEMA_signal_16520), .Q (new_AGEMA_signal_16521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8700 ( .C (clk), .D (new_AGEMA_signal_16524), .Q (new_AGEMA_signal_16525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8704 ( .C (clk), .D (new_AGEMA_signal_16528), .Q (new_AGEMA_signal_16529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8708 ( .C (clk), .D (new_AGEMA_signal_16532), .Q (new_AGEMA_signal_16533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8712 ( .C (clk), .D (new_AGEMA_signal_16536), .Q (new_AGEMA_signal_16537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8716 ( .C (clk), .D (new_AGEMA_signal_16540), .Q (new_AGEMA_signal_16541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8720 ( .C (clk), .D (new_AGEMA_signal_16544), .Q (new_AGEMA_signal_16545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8724 ( .C (clk), .D (new_AGEMA_signal_16548), .Q (new_AGEMA_signal_16549) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8728 ( .C (clk), .D (new_AGEMA_signal_16552), .Q (new_AGEMA_signal_16553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8732 ( .C (clk), .D (new_AGEMA_signal_16556), .Q (new_AGEMA_signal_16557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8736 ( .C (clk), .D (new_AGEMA_signal_16560), .Q (new_AGEMA_signal_16561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8740 ( .C (clk), .D (new_AGEMA_signal_16564), .Q (new_AGEMA_signal_16565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8744 ( .C (clk), .D (new_AGEMA_signal_16568), .Q (new_AGEMA_signal_16569) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8748 ( .C (clk), .D (new_AGEMA_signal_16572), .Q (new_AGEMA_signal_16573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8752 ( .C (clk), .D (new_AGEMA_signal_16576), .Q (new_AGEMA_signal_16577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8756 ( .C (clk), .D (new_AGEMA_signal_16580), .Q (new_AGEMA_signal_16581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8760 ( .C (clk), .D (new_AGEMA_signal_16584), .Q (new_AGEMA_signal_16585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8764 ( .C (clk), .D (new_AGEMA_signal_16588), .Q (new_AGEMA_signal_16589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8768 ( .C (clk), .D (new_AGEMA_signal_16592), .Q (new_AGEMA_signal_16593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8772 ( .C (clk), .D (new_AGEMA_signal_16596), .Q (new_AGEMA_signal_16597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8776 ( .C (clk), .D (new_AGEMA_signal_16600), .Q (new_AGEMA_signal_16601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8780 ( .C (clk), .D (new_AGEMA_signal_16604), .Q (new_AGEMA_signal_16605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8784 ( .C (clk), .D (new_AGEMA_signal_16608), .Q (new_AGEMA_signal_16609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8788 ( .C (clk), .D (new_AGEMA_signal_16612), .Q (new_AGEMA_signal_16613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8792 ( .C (clk), .D (new_AGEMA_signal_16616), .Q (new_AGEMA_signal_16617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8796 ( .C (clk), .D (new_AGEMA_signal_16620), .Q (new_AGEMA_signal_16621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8800 ( .C (clk), .D (new_AGEMA_signal_16624), .Q (new_AGEMA_signal_16625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8804 ( .C (clk), .D (new_AGEMA_signal_16628), .Q (new_AGEMA_signal_16629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8808 ( .C (clk), .D (new_AGEMA_signal_16632), .Q (new_AGEMA_signal_16633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8812 ( .C (clk), .D (new_AGEMA_signal_16636), .Q (new_AGEMA_signal_16637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8816 ( .C (clk), .D (new_AGEMA_signal_16640), .Q (new_AGEMA_signal_16641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8820 ( .C (clk), .D (new_AGEMA_signal_16644), .Q (new_AGEMA_signal_16645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8824 ( .C (clk), .D (new_AGEMA_signal_16648), .Q (new_AGEMA_signal_16649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8828 ( .C (clk), .D (new_AGEMA_signal_16652), .Q (new_AGEMA_signal_16653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8832 ( .C (clk), .D (new_AGEMA_signal_16656), .Q (new_AGEMA_signal_16657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8836 ( .C (clk), .D (new_AGEMA_signal_16660), .Q (new_AGEMA_signal_16661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8840 ( .C (clk), .D (new_AGEMA_signal_16664), .Q (new_AGEMA_signal_16665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8844 ( .C (clk), .D (new_AGEMA_signal_16668), .Q (new_AGEMA_signal_16669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8848 ( .C (clk), .D (new_AGEMA_signal_16672), .Q (new_AGEMA_signal_16673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8852 ( .C (clk), .D (new_AGEMA_signal_16676), .Q (new_AGEMA_signal_16677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8856 ( .C (clk), .D (new_AGEMA_signal_16680), .Q (new_AGEMA_signal_16681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8860 ( .C (clk), .D (new_AGEMA_signal_16684), .Q (new_AGEMA_signal_16685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8864 ( .C (clk), .D (new_AGEMA_signal_16688), .Q (new_AGEMA_signal_16689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8868 ( .C (clk), .D (new_AGEMA_signal_16692), .Q (new_AGEMA_signal_16693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8872 ( .C (clk), .D (new_AGEMA_signal_16696), .Q (new_AGEMA_signal_16697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8876 ( .C (clk), .D (new_AGEMA_signal_16700), .Q (new_AGEMA_signal_16701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8880 ( .C (clk), .D (new_AGEMA_signal_16704), .Q (new_AGEMA_signal_16705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8884 ( .C (clk), .D (new_AGEMA_signal_16708), .Q (new_AGEMA_signal_16709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8888 ( .C (clk), .D (new_AGEMA_signal_16712), .Q (new_AGEMA_signal_16713) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8892 ( .C (clk), .D (new_AGEMA_signal_16716), .Q (new_AGEMA_signal_16717) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8896 ( .C (clk), .D (new_AGEMA_signal_16720), .Q (new_AGEMA_signal_16721) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8900 ( .C (clk), .D (new_AGEMA_signal_16724), .Q (new_AGEMA_signal_16725) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8904 ( .C (clk), .D (new_AGEMA_signal_16728), .Q (new_AGEMA_signal_16729) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8908 ( .C (clk), .D (new_AGEMA_signal_16732), .Q (new_AGEMA_signal_16733) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8912 ( .C (clk), .D (new_AGEMA_signal_16736), .Q (new_AGEMA_signal_16737) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8916 ( .C (clk), .D (new_AGEMA_signal_16740), .Q (new_AGEMA_signal_16741) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8920 ( .C (clk), .D (new_AGEMA_signal_16744), .Q (new_AGEMA_signal_16745) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8924 ( .C (clk), .D (new_AGEMA_signal_16748), .Q (new_AGEMA_signal_16749) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8928 ( .C (clk), .D (new_AGEMA_signal_16752), .Q (new_AGEMA_signal_16753) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8932 ( .C (clk), .D (new_AGEMA_signal_16756), .Q (new_AGEMA_signal_16757) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8936 ( .C (clk), .D (new_AGEMA_signal_16760), .Q (new_AGEMA_signal_16761) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8940 ( .C (clk), .D (new_AGEMA_signal_16764), .Q (new_AGEMA_signal_16765) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8944 ( .C (clk), .D (new_AGEMA_signal_16768), .Q (new_AGEMA_signal_16769) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8948 ( .C (clk), .D (new_AGEMA_signal_16772), .Q (new_AGEMA_signal_16773) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8952 ( .C (clk), .D (new_AGEMA_signal_16776), .Q (new_AGEMA_signal_16777) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8956 ( .C (clk), .D (new_AGEMA_signal_16780), .Q (new_AGEMA_signal_16781) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8960 ( .C (clk), .D (new_AGEMA_signal_16784), .Q (new_AGEMA_signal_16785) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8964 ( .C (clk), .D (new_AGEMA_signal_16788), .Q (new_AGEMA_signal_16789) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8968 ( .C (clk), .D (new_AGEMA_signal_16792), .Q (new_AGEMA_signal_16793) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8972 ( .C (clk), .D (new_AGEMA_signal_16796), .Q (new_AGEMA_signal_16797) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8976 ( .C (clk), .D (new_AGEMA_signal_16800), .Q (new_AGEMA_signal_16801) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8980 ( .C (clk), .D (new_AGEMA_signal_16804), .Q (new_AGEMA_signal_16805) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8984 ( .C (clk), .D (new_AGEMA_signal_16808), .Q (new_AGEMA_signal_16809) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8988 ( .C (clk), .D (new_AGEMA_signal_16812), .Q (new_AGEMA_signal_16813) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8992 ( .C (clk), .D (new_AGEMA_signal_16816), .Q (new_AGEMA_signal_16817) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_8996 ( .C (clk), .D (new_AGEMA_signal_16820), .Q (new_AGEMA_signal_16821) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9000 ( .C (clk), .D (new_AGEMA_signal_16824), .Q (new_AGEMA_signal_16825) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9004 ( .C (clk), .D (new_AGEMA_signal_16828), .Q (new_AGEMA_signal_16829) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9008 ( .C (clk), .D (new_AGEMA_signal_16832), .Q (new_AGEMA_signal_16833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9012 ( .C (clk), .D (new_AGEMA_signal_16836), .Q (new_AGEMA_signal_16837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9016 ( .C (clk), .D (new_AGEMA_signal_16840), .Q (new_AGEMA_signal_16841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9020 ( .C (clk), .D (new_AGEMA_signal_16844), .Q (new_AGEMA_signal_16845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9024 ( .C (clk), .D (new_AGEMA_signal_16848), .Q (new_AGEMA_signal_16849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9028 ( .C (clk), .D (new_AGEMA_signal_16852), .Q (new_AGEMA_signal_16853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9032 ( .C (clk), .D (new_AGEMA_signal_16856), .Q (new_AGEMA_signal_16857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9036 ( .C (clk), .D (new_AGEMA_signal_16860), .Q (new_AGEMA_signal_16861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9040 ( .C (clk), .D (new_AGEMA_signal_16864), .Q (new_AGEMA_signal_16865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9044 ( .C (clk), .D (new_AGEMA_signal_16868), .Q (new_AGEMA_signal_16869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9048 ( .C (clk), .D (new_AGEMA_signal_16872), .Q (new_AGEMA_signal_16873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9052 ( .C (clk), .D (new_AGEMA_signal_16876), .Q (new_AGEMA_signal_16877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9056 ( .C (clk), .D (new_AGEMA_signal_16880), .Q (new_AGEMA_signal_16881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9060 ( .C (clk), .D (new_AGEMA_signal_16884), .Q (new_AGEMA_signal_16885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9064 ( .C (clk), .D (new_AGEMA_signal_16888), .Q (new_AGEMA_signal_16889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9068 ( .C (clk), .D (new_AGEMA_signal_16892), .Q (new_AGEMA_signal_16893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9072 ( .C (clk), .D (new_AGEMA_signal_16896), .Q (new_AGEMA_signal_16897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9076 ( .C (clk), .D (new_AGEMA_signal_16900), .Q (new_AGEMA_signal_16901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9080 ( .C (clk), .D (new_AGEMA_signal_16904), .Q (new_AGEMA_signal_16905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9084 ( .C (clk), .D (new_AGEMA_signal_16908), .Q (new_AGEMA_signal_16909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9088 ( .C (clk), .D (new_AGEMA_signal_16912), .Q (new_AGEMA_signal_16913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9092 ( .C (clk), .D (new_AGEMA_signal_16916), .Q (new_AGEMA_signal_16917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9096 ( .C (clk), .D (new_AGEMA_signal_16920), .Q (new_AGEMA_signal_16921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9100 ( .C (clk), .D (new_AGEMA_signal_16924), .Q (new_AGEMA_signal_16925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9104 ( .C (clk), .D (new_AGEMA_signal_16928), .Q (new_AGEMA_signal_16929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9108 ( .C (clk), .D (new_AGEMA_signal_16932), .Q (new_AGEMA_signal_16933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9112 ( .C (clk), .D (new_AGEMA_signal_16936), .Q (new_AGEMA_signal_16937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9116 ( .C (clk), .D (new_AGEMA_signal_16940), .Q (new_AGEMA_signal_16941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9120 ( .C (clk), .D (new_AGEMA_signal_16944), .Q (new_AGEMA_signal_16945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9124 ( .C (clk), .D (new_AGEMA_signal_16948), .Q (new_AGEMA_signal_16949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9128 ( .C (clk), .D (new_AGEMA_signal_16952), .Q (new_AGEMA_signal_16953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9132 ( .C (clk), .D (new_AGEMA_signal_16956), .Q (new_AGEMA_signal_16957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9136 ( .C (clk), .D (new_AGEMA_signal_16960), .Q (new_AGEMA_signal_16961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9140 ( .C (clk), .D (new_AGEMA_signal_16964), .Q (new_AGEMA_signal_16965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9144 ( .C (clk), .D (new_AGEMA_signal_16968), .Q (new_AGEMA_signal_16969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9148 ( .C (clk), .D (new_AGEMA_signal_16972), .Q (new_AGEMA_signal_16973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9152 ( .C (clk), .D (new_AGEMA_signal_16976), .Q (new_AGEMA_signal_16977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9156 ( .C (clk), .D (new_AGEMA_signal_16980), .Q (new_AGEMA_signal_16981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9160 ( .C (clk), .D (new_AGEMA_signal_16984), .Q (new_AGEMA_signal_16985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9164 ( .C (clk), .D (new_AGEMA_signal_16988), .Q (new_AGEMA_signal_16989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9168 ( .C (clk), .D (new_AGEMA_signal_16992), .Q (new_AGEMA_signal_16993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9172 ( .C (clk), .D (new_AGEMA_signal_16996), .Q (new_AGEMA_signal_16997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9176 ( .C (clk), .D (new_AGEMA_signal_17000), .Q (new_AGEMA_signal_17001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9180 ( .C (clk), .D (new_AGEMA_signal_17004), .Q (new_AGEMA_signal_17005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9184 ( .C (clk), .D (new_AGEMA_signal_17008), .Q (new_AGEMA_signal_17009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9188 ( .C (clk), .D (new_AGEMA_signal_17012), .Q (new_AGEMA_signal_17013) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9192 ( .C (clk), .D (new_AGEMA_signal_17016), .Q (new_AGEMA_signal_17017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9196 ( .C (clk), .D (new_AGEMA_signal_17020), .Q (new_AGEMA_signal_17021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9200 ( .C (clk), .D (new_AGEMA_signal_17024), .Q (new_AGEMA_signal_17025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9204 ( .C (clk), .D (new_AGEMA_signal_17028), .Q (new_AGEMA_signal_17029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9208 ( .C (clk), .D (new_AGEMA_signal_17032), .Q (new_AGEMA_signal_17033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9212 ( .C (clk), .D (new_AGEMA_signal_17036), .Q (new_AGEMA_signal_17037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9216 ( .C (clk), .D (new_AGEMA_signal_17040), .Q (new_AGEMA_signal_17041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9220 ( .C (clk), .D (new_AGEMA_signal_17044), .Q (new_AGEMA_signal_17045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9224 ( .C (clk), .D (new_AGEMA_signal_17048), .Q (new_AGEMA_signal_17049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9228 ( .C (clk), .D (new_AGEMA_signal_17052), .Q (new_AGEMA_signal_17053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9232 ( .C (clk), .D (new_AGEMA_signal_17056), .Q (new_AGEMA_signal_17057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9236 ( .C (clk), .D (new_AGEMA_signal_17060), .Q (new_AGEMA_signal_17061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9240 ( .C (clk), .D (new_AGEMA_signal_17064), .Q (new_AGEMA_signal_17065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9244 ( .C (clk), .D (new_AGEMA_signal_17068), .Q (new_AGEMA_signal_17069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9248 ( .C (clk), .D (new_AGEMA_signal_17072), .Q (new_AGEMA_signal_17073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9252 ( .C (clk), .D (new_AGEMA_signal_17076), .Q (new_AGEMA_signal_17077) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9256 ( .C (clk), .D (new_AGEMA_signal_17080), .Q (new_AGEMA_signal_17081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9260 ( .C (clk), .D (new_AGEMA_signal_17084), .Q (new_AGEMA_signal_17085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9264 ( .C (clk), .D (new_AGEMA_signal_17088), .Q (new_AGEMA_signal_17089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9268 ( .C (clk), .D (new_AGEMA_signal_17092), .Q (new_AGEMA_signal_17093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9272 ( .C (clk), .D (new_AGEMA_signal_17096), .Q (new_AGEMA_signal_17097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9276 ( .C (clk), .D (new_AGEMA_signal_17100), .Q (new_AGEMA_signal_17101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9280 ( .C (clk), .D (new_AGEMA_signal_17104), .Q (new_AGEMA_signal_17105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9284 ( .C (clk), .D (new_AGEMA_signal_17108), .Q (new_AGEMA_signal_17109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9288 ( .C (clk), .D (new_AGEMA_signal_17112), .Q (new_AGEMA_signal_17113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9292 ( .C (clk), .D (new_AGEMA_signal_17116), .Q (new_AGEMA_signal_17117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9296 ( .C (clk), .D (new_AGEMA_signal_17120), .Q (new_AGEMA_signal_17121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9300 ( .C (clk), .D (new_AGEMA_signal_17124), .Q (new_AGEMA_signal_17125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9304 ( .C (clk), .D (new_AGEMA_signal_17128), .Q (new_AGEMA_signal_17129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9308 ( .C (clk), .D (new_AGEMA_signal_17132), .Q (new_AGEMA_signal_17133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9312 ( .C (clk), .D (new_AGEMA_signal_17136), .Q (new_AGEMA_signal_17137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9316 ( .C (clk), .D (new_AGEMA_signal_17140), .Q (new_AGEMA_signal_17141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9320 ( .C (clk), .D (new_AGEMA_signal_17144), .Q (new_AGEMA_signal_17145) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9324 ( .C (clk), .D (new_AGEMA_signal_17148), .Q (new_AGEMA_signal_17149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9328 ( .C (clk), .D (new_AGEMA_signal_17152), .Q (new_AGEMA_signal_17153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9332 ( .C (clk), .D (new_AGEMA_signal_17156), .Q (new_AGEMA_signal_17157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9336 ( .C (clk), .D (new_AGEMA_signal_17160), .Q (new_AGEMA_signal_17161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9340 ( .C (clk), .D (new_AGEMA_signal_17164), .Q (new_AGEMA_signal_17165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9344 ( .C (clk), .D (new_AGEMA_signal_17168), .Q (new_AGEMA_signal_17169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9348 ( .C (clk), .D (new_AGEMA_signal_17172), .Q (new_AGEMA_signal_17173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9352 ( .C (clk), .D (new_AGEMA_signal_17176), .Q (new_AGEMA_signal_17177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9356 ( .C (clk), .D (new_AGEMA_signal_17180), .Q (new_AGEMA_signal_17181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9360 ( .C (clk), .D (new_AGEMA_signal_17184), .Q (new_AGEMA_signal_17185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9364 ( .C (clk), .D (new_AGEMA_signal_17188), .Q (new_AGEMA_signal_17189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9368 ( .C (clk), .D (new_AGEMA_signal_17192), .Q (new_AGEMA_signal_17193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9372 ( .C (clk), .D (new_AGEMA_signal_17196), .Q (new_AGEMA_signal_17197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9376 ( .C (clk), .D (new_AGEMA_signal_17200), .Q (new_AGEMA_signal_17201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9380 ( .C (clk), .D (new_AGEMA_signal_17204), .Q (new_AGEMA_signal_17205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9384 ( .C (clk), .D (new_AGEMA_signal_17208), .Q (new_AGEMA_signal_17209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9388 ( .C (clk), .D (new_AGEMA_signal_17212), .Q (new_AGEMA_signal_17213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9392 ( .C (clk), .D (new_AGEMA_signal_17216), .Q (new_AGEMA_signal_17217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9396 ( .C (clk), .D (new_AGEMA_signal_17220), .Q (new_AGEMA_signal_17221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9400 ( .C (clk), .D (new_AGEMA_signal_17224), .Q (new_AGEMA_signal_17225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9404 ( .C (clk), .D (new_AGEMA_signal_17228), .Q (new_AGEMA_signal_17229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9408 ( .C (clk), .D (new_AGEMA_signal_17232), .Q (new_AGEMA_signal_17233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9412 ( .C (clk), .D (new_AGEMA_signal_17236), .Q (new_AGEMA_signal_17237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9416 ( .C (clk), .D (new_AGEMA_signal_17240), .Q (new_AGEMA_signal_17241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9420 ( .C (clk), .D (new_AGEMA_signal_17244), .Q (new_AGEMA_signal_17245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9424 ( .C (clk), .D (new_AGEMA_signal_17248), .Q (new_AGEMA_signal_17249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9428 ( .C (clk), .D (new_AGEMA_signal_17252), .Q (new_AGEMA_signal_17253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9432 ( .C (clk), .D (new_AGEMA_signal_17256), .Q (new_AGEMA_signal_17257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9436 ( .C (clk), .D (new_AGEMA_signal_17260), .Q (new_AGEMA_signal_17261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9440 ( .C (clk), .D (new_AGEMA_signal_17264), .Q (new_AGEMA_signal_17265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9444 ( .C (clk), .D (new_AGEMA_signal_17268), .Q (new_AGEMA_signal_17269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9448 ( .C (clk), .D (new_AGEMA_signal_17272), .Q (new_AGEMA_signal_17273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9452 ( .C (clk), .D (new_AGEMA_signal_17276), .Q (new_AGEMA_signal_17277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9456 ( .C (clk), .D (new_AGEMA_signal_17280), .Q (new_AGEMA_signal_17281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9460 ( .C (clk), .D (new_AGEMA_signal_17284), .Q (new_AGEMA_signal_17285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9464 ( .C (clk), .D (new_AGEMA_signal_17288), .Q (new_AGEMA_signal_17289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9468 ( .C (clk), .D (new_AGEMA_signal_17292), .Q (new_AGEMA_signal_17293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9472 ( .C (clk), .D (new_AGEMA_signal_17296), .Q (new_AGEMA_signal_17297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9476 ( .C (clk), .D (new_AGEMA_signal_17300), .Q (new_AGEMA_signal_17301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9480 ( .C (clk), .D (new_AGEMA_signal_17304), .Q (new_AGEMA_signal_17305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9484 ( .C (clk), .D (new_AGEMA_signal_17308), .Q (new_AGEMA_signal_17309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9488 ( .C (clk), .D (new_AGEMA_signal_17312), .Q (new_AGEMA_signal_17313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9492 ( .C (clk), .D (new_AGEMA_signal_17316), .Q (new_AGEMA_signal_17317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9496 ( .C (clk), .D (new_AGEMA_signal_17320), .Q (new_AGEMA_signal_17321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9500 ( .C (clk), .D (new_AGEMA_signal_17324), .Q (new_AGEMA_signal_17325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9504 ( .C (clk), .D (new_AGEMA_signal_17328), .Q (new_AGEMA_signal_17329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9508 ( .C (clk), .D (new_AGEMA_signal_17332), .Q (new_AGEMA_signal_17333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9512 ( .C (clk), .D (new_AGEMA_signal_17336), .Q (new_AGEMA_signal_17337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9516 ( .C (clk), .D (new_AGEMA_signal_17340), .Q (new_AGEMA_signal_17341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9520 ( .C (clk), .D (new_AGEMA_signal_17344), .Q (new_AGEMA_signal_17345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9524 ( .C (clk), .D (new_AGEMA_signal_17348), .Q (new_AGEMA_signal_17349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9528 ( .C (clk), .D (new_AGEMA_signal_17352), .Q (new_AGEMA_signal_17353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9532 ( .C (clk), .D (new_AGEMA_signal_17356), .Q (new_AGEMA_signal_17357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9536 ( .C (clk), .D (new_AGEMA_signal_17360), .Q (new_AGEMA_signal_17361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9540 ( .C (clk), .D (new_AGEMA_signal_17364), .Q (new_AGEMA_signal_17365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9544 ( .C (clk), .D (new_AGEMA_signal_17368), .Q (new_AGEMA_signal_17369) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9548 ( .C (clk), .D (new_AGEMA_signal_17372), .Q (new_AGEMA_signal_17373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9552 ( .C (clk), .D (new_AGEMA_signal_17376), .Q (new_AGEMA_signal_17377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9556 ( .C (clk), .D (new_AGEMA_signal_17380), .Q (new_AGEMA_signal_17381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9560 ( .C (clk), .D (new_AGEMA_signal_17384), .Q (new_AGEMA_signal_17385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9564 ( .C (clk), .D (new_AGEMA_signal_17388), .Q (new_AGEMA_signal_17389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9568 ( .C (clk), .D (new_AGEMA_signal_17392), .Q (new_AGEMA_signal_17393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9572 ( .C (clk), .D (new_AGEMA_signal_17396), .Q (new_AGEMA_signal_17397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9576 ( .C (clk), .D (new_AGEMA_signal_17400), .Q (new_AGEMA_signal_17401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9580 ( .C (clk), .D (new_AGEMA_signal_17404), .Q (new_AGEMA_signal_17405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9584 ( .C (clk), .D (new_AGEMA_signal_17408), .Q (new_AGEMA_signal_17409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9588 ( .C (clk), .D (new_AGEMA_signal_17412), .Q (new_AGEMA_signal_17413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9592 ( .C (clk), .D (new_AGEMA_signal_17416), .Q (new_AGEMA_signal_17417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9596 ( .C (clk), .D (new_AGEMA_signal_17420), .Q (new_AGEMA_signal_17421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9600 ( .C (clk), .D (new_AGEMA_signal_17424), .Q (new_AGEMA_signal_17425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9604 ( .C (clk), .D (new_AGEMA_signal_17428), .Q (new_AGEMA_signal_17429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9608 ( .C (clk), .D (new_AGEMA_signal_17432), .Q (new_AGEMA_signal_17433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9612 ( .C (clk), .D (new_AGEMA_signal_17436), .Q (new_AGEMA_signal_17437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9616 ( .C (clk), .D (new_AGEMA_signal_17440), .Q (new_AGEMA_signal_17441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9620 ( .C (clk), .D (new_AGEMA_signal_17444), .Q (new_AGEMA_signal_17445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9624 ( .C (clk), .D (new_AGEMA_signal_17448), .Q (new_AGEMA_signal_17449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9628 ( .C (clk), .D (new_AGEMA_signal_17452), .Q (new_AGEMA_signal_17453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9632 ( .C (clk), .D (new_AGEMA_signal_17456), .Q (new_AGEMA_signal_17457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9636 ( .C (clk), .D (new_AGEMA_signal_17460), .Q (new_AGEMA_signal_17461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9640 ( .C (clk), .D (new_AGEMA_signal_17464), .Q (new_AGEMA_signal_17465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9644 ( .C (clk), .D (new_AGEMA_signal_17468), .Q (new_AGEMA_signal_17469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9648 ( .C (clk), .D (new_AGEMA_signal_17472), .Q (new_AGEMA_signal_17473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9652 ( .C (clk), .D (new_AGEMA_signal_17476), .Q (new_AGEMA_signal_17477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9656 ( .C (clk), .D (new_AGEMA_signal_17480), .Q (new_AGEMA_signal_17481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9660 ( .C (clk), .D (new_AGEMA_signal_17484), .Q (new_AGEMA_signal_17485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9664 ( .C (clk), .D (new_AGEMA_signal_17488), .Q (new_AGEMA_signal_17489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9668 ( .C (clk), .D (new_AGEMA_signal_17492), .Q (new_AGEMA_signal_17493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9672 ( .C (clk), .D (new_AGEMA_signal_17496), .Q (new_AGEMA_signal_17497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9676 ( .C (clk), .D (new_AGEMA_signal_17500), .Q (new_AGEMA_signal_17501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9680 ( .C (clk), .D (new_AGEMA_signal_17504), .Q (new_AGEMA_signal_17505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9684 ( .C (clk), .D (new_AGEMA_signal_17508), .Q (new_AGEMA_signal_17509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9688 ( .C (clk), .D (new_AGEMA_signal_17512), .Q (new_AGEMA_signal_17513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9692 ( .C (clk), .D (new_AGEMA_signal_17516), .Q (new_AGEMA_signal_17517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9696 ( .C (clk), .D (new_AGEMA_signal_17520), .Q (new_AGEMA_signal_17521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9700 ( .C (clk), .D (new_AGEMA_signal_17524), .Q (new_AGEMA_signal_17525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9704 ( .C (clk), .D (new_AGEMA_signal_17528), .Q (new_AGEMA_signal_17529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9708 ( .C (clk), .D (new_AGEMA_signal_17532), .Q (new_AGEMA_signal_17533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9712 ( .C (clk), .D (new_AGEMA_signal_17536), .Q (new_AGEMA_signal_17537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9716 ( .C (clk), .D (new_AGEMA_signal_17540), .Q (new_AGEMA_signal_17541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9720 ( .C (clk), .D (new_AGEMA_signal_17544), .Q (new_AGEMA_signal_17545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9724 ( .C (clk), .D (new_AGEMA_signal_17548), .Q (new_AGEMA_signal_17549) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9728 ( .C (clk), .D (new_AGEMA_signal_17552), .Q (new_AGEMA_signal_17553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9732 ( .C (clk), .D (new_AGEMA_signal_17556), .Q (new_AGEMA_signal_17557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9736 ( .C (clk), .D (new_AGEMA_signal_17560), .Q (new_AGEMA_signal_17561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9740 ( .C (clk), .D (new_AGEMA_signal_17564), .Q (new_AGEMA_signal_17565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9744 ( .C (clk), .D (new_AGEMA_signal_17568), .Q (new_AGEMA_signal_17569) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9748 ( .C (clk), .D (new_AGEMA_signal_17572), .Q (new_AGEMA_signal_17573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9752 ( .C (clk), .D (new_AGEMA_signal_17576), .Q (new_AGEMA_signal_17577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9756 ( .C (clk), .D (new_AGEMA_signal_17580), .Q (new_AGEMA_signal_17581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9760 ( .C (clk), .D (new_AGEMA_signal_17584), .Q (new_AGEMA_signal_17585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9764 ( .C (clk), .D (new_AGEMA_signal_17588), .Q (new_AGEMA_signal_17589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9768 ( .C (clk), .D (new_AGEMA_signal_17592), .Q (new_AGEMA_signal_17593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9772 ( .C (clk), .D (new_AGEMA_signal_17596), .Q (new_AGEMA_signal_17597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9776 ( .C (clk), .D (new_AGEMA_signal_17600), .Q (new_AGEMA_signal_17601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9780 ( .C (clk), .D (new_AGEMA_signal_17604), .Q (new_AGEMA_signal_17605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9784 ( .C (clk), .D (new_AGEMA_signal_17608), .Q (new_AGEMA_signal_17609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9788 ( .C (clk), .D (new_AGEMA_signal_17612), .Q (new_AGEMA_signal_17613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9792 ( .C (clk), .D (new_AGEMA_signal_17616), .Q (new_AGEMA_signal_17617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9796 ( .C (clk), .D (new_AGEMA_signal_17620), .Q (new_AGEMA_signal_17621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9800 ( .C (clk), .D (new_AGEMA_signal_17624), .Q (new_AGEMA_signal_17625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9804 ( .C (clk), .D (new_AGEMA_signal_17628), .Q (new_AGEMA_signal_17629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9808 ( .C (clk), .D (new_AGEMA_signal_17632), .Q (new_AGEMA_signal_17633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9812 ( .C (clk), .D (new_AGEMA_signal_17636), .Q (new_AGEMA_signal_17637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9816 ( .C (clk), .D (new_AGEMA_signal_17640), .Q (new_AGEMA_signal_17641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9820 ( .C (clk), .D (new_AGEMA_signal_17644), .Q (new_AGEMA_signal_17645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9824 ( .C (clk), .D (new_AGEMA_signal_17648), .Q (new_AGEMA_signal_17649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9828 ( .C (clk), .D (new_AGEMA_signal_17652), .Q (new_AGEMA_signal_17653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9832 ( .C (clk), .D (new_AGEMA_signal_17656), .Q (new_AGEMA_signal_17657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9836 ( .C (clk), .D (new_AGEMA_signal_17660), .Q (new_AGEMA_signal_17661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9840 ( .C (clk), .D (new_AGEMA_signal_17664), .Q (new_AGEMA_signal_17665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9844 ( .C (clk), .D (new_AGEMA_signal_17668), .Q (new_AGEMA_signal_17669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9848 ( .C (clk), .D (new_AGEMA_signal_17672), .Q (new_AGEMA_signal_17673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9852 ( .C (clk), .D (new_AGEMA_signal_17676), .Q (new_AGEMA_signal_17677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9856 ( .C (clk), .D (new_AGEMA_signal_17680), .Q (new_AGEMA_signal_17681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9860 ( .C (clk), .D (new_AGEMA_signal_17684), .Q (new_AGEMA_signal_17685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9864 ( .C (clk), .D (new_AGEMA_signal_17688), .Q (new_AGEMA_signal_17689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9868 ( .C (clk), .D (new_AGEMA_signal_17692), .Q (new_AGEMA_signal_17693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9872 ( .C (clk), .D (new_AGEMA_signal_17696), .Q (new_AGEMA_signal_17697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_9876 ( .C (clk), .D (new_AGEMA_signal_17700), .Q (new_AGEMA_signal_17701) ) ;
    buf_clk new_AGEMA_reg_buffer_9880 ( .C (clk), .D (new_AGEMA_signal_17704), .Q (new_AGEMA_signal_17705) ) ;
    buf_clk new_AGEMA_reg_buffer_9884 ( .C (clk), .D (new_AGEMA_signal_17708), .Q (new_AGEMA_signal_17709) ) ;
    buf_clk new_AGEMA_reg_buffer_9888 ( .C (clk), .D (new_AGEMA_signal_17712), .Q (new_AGEMA_signal_17713) ) ;
    buf_clk new_AGEMA_reg_buffer_9892 ( .C (clk), .D (new_AGEMA_signal_17716), .Q (new_AGEMA_signal_17717) ) ;
    buf_clk new_AGEMA_reg_buffer_9896 ( .C (clk), .D (new_AGEMA_signal_17720), .Q (new_AGEMA_signal_17721) ) ;
    buf_clk new_AGEMA_reg_buffer_9900 ( .C (clk), .D (new_AGEMA_signal_17724), .Q (new_AGEMA_signal_17725) ) ;
    buf_clk new_AGEMA_reg_buffer_9904 ( .C (clk), .D (new_AGEMA_signal_17728), .Q (new_AGEMA_signal_17729) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7794, new_AGEMA_signal_7793, new_AGEMA_signal_7792, RoundReg_Inst_ff_SDE_0_next_state}), .clk (clk), .Q ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8145, new_AGEMA_signal_8144, new_AGEMA_signal_8143, RoundReg_Inst_ff_SDE_1_next_state}), .clk (clk), .Q ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7800, new_AGEMA_signal_7799, new_AGEMA_signal_7798, RoundReg_Inst_ff_SDE_2_next_state}), .clk (clk), .Q ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8151, new_AGEMA_signal_8150, new_AGEMA_signal_8149, RoundReg_Inst_ff_SDE_3_next_state}), .clk (clk), .Q ({ciphertext_s3[35], ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8157, new_AGEMA_signal_8156, new_AGEMA_signal_8155, RoundReg_Inst_ff_SDE_4_next_state}), .clk (clk), .Q ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7806, new_AGEMA_signal_7805, new_AGEMA_signal_7804, RoundReg_Inst_ff_SDE_5_next_state}), .clk (clk), .Q ({ciphertext_s3[37], ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7812, new_AGEMA_signal_7811, new_AGEMA_signal_7810, RoundReg_Inst_ff_SDE_6_next_state}), .clk (clk), .Q ({ciphertext_s3[38], ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7818, new_AGEMA_signal_7817, new_AGEMA_signal_7816, RoundReg_Inst_ff_SDE_7_next_state}), .clk (clk), .Q ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7824, new_AGEMA_signal_7823, new_AGEMA_signal_7822, RoundReg_Inst_ff_SDE_8_next_state}), .clk (clk), .Q ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8163, new_AGEMA_signal_8162, new_AGEMA_signal_8161, RoundReg_Inst_ff_SDE_9_next_state}), .clk (clk), .Q ({ciphertext_s3[73], ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7830, new_AGEMA_signal_7829, new_AGEMA_signal_7828, RoundReg_Inst_ff_SDE_10_next_state}), .clk (clk), .Q ({ciphertext_s3[74], ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8169, new_AGEMA_signal_8168, new_AGEMA_signal_8167, RoundReg_Inst_ff_SDE_11_next_state}), .clk (clk), .Q ({ciphertext_s3[75], ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8175, new_AGEMA_signal_8174, new_AGEMA_signal_8173, RoundReg_Inst_ff_SDE_12_next_state}), .clk (clk), .Q ({ciphertext_s3[76], ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7836, new_AGEMA_signal_7835, new_AGEMA_signal_7834, RoundReg_Inst_ff_SDE_13_next_state}), .clk (clk), .Q ({ciphertext_s3[77], ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7842, new_AGEMA_signal_7841, new_AGEMA_signal_7840, RoundReg_Inst_ff_SDE_14_next_state}), .clk (clk), .Q ({ciphertext_s3[78], ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7848, new_AGEMA_signal_7847, new_AGEMA_signal_7846, RoundReg_Inst_ff_SDE_15_next_state}), .clk (clk), .Q ({ciphertext_s3[79], ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, new_AGEMA_signal_7852, RoundReg_Inst_ff_SDE_16_next_state}), .clk (clk), .Q ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8181, new_AGEMA_signal_8180, new_AGEMA_signal_8179, RoundReg_Inst_ff_SDE_17_next_state}), .clk (clk), .Q ({ciphertext_s3[113], ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7860, new_AGEMA_signal_7859, new_AGEMA_signal_7858, RoundReg_Inst_ff_SDE_18_next_state}), .clk (clk), .Q ({ciphertext_s3[114], ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8187, new_AGEMA_signal_8186, new_AGEMA_signal_8185, RoundReg_Inst_ff_SDE_19_next_state}), .clk (clk), .Q ({ciphertext_s3[115], ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8193, new_AGEMA_signal_8192, new_AGEMA_signal_8191, RoundReg_Inst_ff_SDE_20_next_state}), .clk (clk), .Q ({ciphertext_s3[116], ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7866, new_AGEMA_signal_7865, new_AGEMA_signal_7864, RoundReg_Inst_ff_SDE_21_next_state}), .clk (clk), .Q ({ciphertext_s3[117], ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7872, new_AGEMA_signal_7871, new_AGEMA_signal_7870, RoundReg_Inst_ff_SDE_22_next_state}), .clk (clk), .Q ({ciphertext_s3[118], ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7878, new_AGEMA_signal_7877, new_AGEMA_signal_7876, RoundReg_Inst_ff_SDE_23_next_state}), .clk (clk), .Q ({ciphertext_s3[119], ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7884, new_AGEMA_signal_7883, new_AGEMA_signal_7882, RoundReg_Inst_ff_SDE_24_next_state}), .clk (clk), .Q ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8199, new_AGEMA_signal_8198, new_AGEMA_signal_8197, RoundReg_Inst_ff_SDE_25_next_state}), .clk (clk), .Q ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7890, new_AGEMA_signal_7889, new_AGEMA_signal_7888, RoundReg_Inst_ff_SDE_26_next_state}), .clk (clk), .Q ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8205, new_AGEMA_signal_8204, new_AGEMA_signal_8203, RoundReg_Inst_ff_SDE_27_next_state}), .clk (clk), .Q ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8211, new_AGEMA_signal_8210, new_AGEMA_signal_8209, RoundReg_Inst_ff_SDE_28_next_state}), .clk (clk), .Q ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7896, new_AGEMA_signal_7895, new_AGEMA_signal_7894, RoundReg_Inst_ff_SDE_29_next_state}), .clk (clk), .Q ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7902, new_AGEMA_signal_7901, new_AGEMA_signal_7900, RoundReg_Inst_ff_SDE_30_next_state}), .clk (clk), .Q ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, new_AGEMA_signal_7906, RoundReg_Inst_ff_SDE_31_next_state}), .clk (clk), .Q ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16181, new_AGEMA_signal_16177, new_AGEMA_signal_16173, new_AGEMA_signal_16169}), .clk (clk), .Q ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16197, new_AGEMA_signal_16193, new_AGEMA_signal_16189, new_AGEMA_signal_16185}), .clk (clk), .Q ({ciphertext_s3[65], ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16213, new_AGEMA_signal_16209, new_AGEMA_signal_16205, new_AGEMA_signal_16201}), .clk (clk), .Q ({ciphertext_s3[66], ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16229, new_AGEMA_signal_16225, new_AGEMA_signal_16221, new_AGEMA_signal_16217}), .clk (clk), .Q ({ciphertext_s3[67], ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16245, new_AGEMA_signal_16241, new_AGEMA_signal_16237, new_AGEMA_signal_16233}), .clk (clk), .Q ({ciphertext_s3[68], ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16261, new_AGEMA_signal_16257, new_AGEMA_signal_16253, new_AGEMA_signal_16249}), .clk (clk), .Q ({ciphertext_s3[69], ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16277, new_AGEMA_signal_16273, new_AGEMA_signal_16269, new_AGEMA_signal_16265}), .clk (clk), .Q ({ciphertext_s3[70], ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16293, new_AGEMA_signal_16289, new_AGEMA_signal_16285, new_AGEMA_signal_16281}), .clk (clk), .Q ({ciphertext_s3[71], ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16309, new_AGEMA_signal_16305, new_AGEMA_signal_16301, new_AGEMA_signal_16297}), .clk (clk), .Q ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16325, new_AGEMA_signal_16321, new_AGEMA_signal_16317, new_AGEMA_signal_16313}), .clk (clk), .Q ({ciphertext_s3[105], ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16341, new_AGEMA_signal_16337, new_AGEMA_signal_16333, new_AGEMA_signal_16329}), .clk (clk), .Q ({ciphertext_s3[106], ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16357, new_AGEMA_signal_16353, new_AGEMA_signal_16349, new_AGEMA_signal_16345}), .clk (clk), .Q ({ciphertext_s3[107], ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16373, new_AGEMA_signal_16369, new_AGEMA_signal_16365, new_AGEMA_signal_16361}), .clk (clk), .Q ({ciphertext_s3[108], ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16389, new_AGEMA_signal_16385, new_AGEMA_signal_16381, new_AGEMA_signal_16377}), .clk (clk), .Q ({ciphertext_s3[109], ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16405, new_AGEMA_signal_16401, new_AGEMA_signal_16397, new_AGEMA_signal_16393}), .clk (clk), .Q ({ciphertext_s3[110], ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16421, new_AGEMA_signal_16417, new_AGEMA_signal_16413, new_AGEMA_signal_16409}), .clk (clk), .Q ({ciphertext_s3[111], ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16437, new_AGEMA_signal_16433, new_AGEMA_signal_16429, new_AGEMA_signal_16425}), .clk (clk), .Q ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16453, new_AGEMA_signal_16449, new_AGEMA_signal_16445, new_AGEMA_signal_16441}), .clk (clk), .Q ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16469, new_AGEMA_signal_16465, new_AGEMA_signal_16461, new_AGEMA_signal_16457}), .clk (clk), .Q ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16485, new_AGEMA_signal_16481, new_AGEMA_signal_16477, new_AGEMA_signal_16473}), .clk (clk), .Q ({ciphertext_s3[19], ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16501, new_AGEMA_signal_16497, new_AGEMA_signal_16493, new_AGEMA_signal_16489}), .clk (clk), .Q ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16517, new_AGEMA_signal_16513, new_AGEMA_signal_16509, new_AGEMA_signal_16505}), .clk (clk), .Q ({ciphertext_s3[21], ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16533, new_AGEMA_signal_16529, new_AGEMA_signal_16525, new_AGEMA_signal_16521}), .clk (clk), .Q ({ciphertext_s3[22], ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16549, new_AGEMA_signal_16545, new_AGEMA_signal_16541, new_AGEMA_signal_16537}), .clk (clk), .Q ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16565, new_AGEMA_signal_16561, new_AGEMA_signal_16557, new_AGEMA_signal_16553}), .clk (clk), .Q ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16581, new_AGEMA_signal_16577, new_AGEMA_signal_16573, new_AGEMA_signal_16569}), .clk (clk), .Q ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16597, new_AGEMA_signal_16593, new_AGEMA_signal_16589, new_AGEMA_signal_16585}), .clk (clk), .Q ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16613, new_AGEMA_signal_16609, new_AGEMA_signal_16605, new_AGEMA_signal_16601}), .clk (clk), .Q ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16629, new_AGEMA_signal_16625, new_AGEMA_signal_16621, new_AGEMA_signal_16617}), .clk (clk), .Q ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16645, new_AGEMA_signal_16641, new_AGEMA_signal_16637, new_AGEMA_signal_16633}), .clk (clk), .Q ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16661, new_AGEMA_signal_16657, new_AGEMA_signal_16653, new_AGEMA_signal_16649}), .clk (clk), .Q ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16677, new_AGEMA_signal_16673, new_AGEMA_signal_16669, new_AGEMA_signal_16665}), .clk (clk), .Q ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16693, new_AGEMA_signal_16689, new_AGEMA_signal_16685, new_AGEMA_signal_16681}), .clk (clk), .Q ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16709, new_AGEMA_signal_16705, new_AGEMA_signal_16701, new_AGEMA_signal_16697}), .clk (clk), .Q ({ciphertext_s3[97], ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16725, new_AGEMA_signal_16721, new_AGEMA_signal_16717, new_AGEMA_signal_16713}), .clk (clk), .Q ({ciphertext_s3[98], ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16741, new_AGEMA_signal_16737, new_AGEMA_signal_16733, new_AGEMA_signal_16729}), .clk (clk), .Q ({ciphertext_s3[99], ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16757, new_AGEMA_signal_16753, new_AGEMA_signal_16749, new_AGEMA_signal_16745}), .clk (clk), .Q ({ciphertext_s3[100], ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16773, new_AGEMA_signal_16769, new_AGEMA_signal_16765, new_AGEMA_signal_16761}), .clk (clk), .Q ({ciphertext_s3[101], ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16789, new_AGEMA_signal_16785, new_AGEMA_signal_16781, new_AGEMA_signal_16777}), .clk (clk), .Q ({ciphertext_s3[102], ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16805, new_AGEMA_signal_16801, new_AGEMA_signal_16797, new_AGEMA_signal_16793}), .clk (clk), .Q ({ciphertext_s3[103], ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16821, new_AGEMA_signal_16817, new_AGEMA_signal_16813, new_AGEMA_signal_16809}), .clk (clk), .Q ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16837, new_AGEMA_signal_16833, new_AGEMA_signal_16829, new_AGEMA_signal_16825}), .clk (clk), .Q ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16853, new_AGEMA_signal_16849, new_AGEMA_signal_16845, new_AGEMA_signal_16841}), .clk (clk), .Q ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16869, new_AGEMA_signal_16865, new_AGEMA_signal_16861, new_AGEMA_signal_16857}), .clk (clk), .Q ({ciphertext_s3[11], ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16885, new_AGEMA_signal_16881, new_AGEMA_signal_16877, new_AGEMA_signal_16873}), .clk (clk), .Q ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16901, new_AGEMA_signal_16897, new_AGEMA_signal_16893, new_AGEMA_signal_16889}), .clk (clk), .Q ({ciphertext_s3[13], ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16917, new_AGEMA_signal_16913, new_AGEMA_signal_16909, new_AGEMA_signal_16905}), .clk (clk), .Q ({ciphertext_s3[14], ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16933, new_AGEMA_signal_16929, new_AGEMA_signal_16925, new_AGEMA_signal_16921}), .clk (clk), .Q ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16949, new_AGEMA_signal_16945, new_AGEMA_signal_16941, new_AGEMA_signal_16937}), .clk (clk), .Q ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16965, new_AGEMA_signal_16961, new_AGEMA_signal_16957, new_AGEMA_signal_16953}), .clk (clk), .Q ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16981, new_AGEMA_signal_16977, new_AGEMA_signal_16973, new_AGEMA_signal_16969}), .clk (clk), .Q ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_16997, new_AGEMA_signal_16993, new_AGEMA_signal_16989, new_AGEMA_signal_16985}), .clk (clk), .Q ({ciphertext_s3[51], ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17013, new_AGEMA_signal_17009, new_AGEMA_signal_17005, new_AGEMA_signal_17001}), .clk (clk), .Q ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17029, new_AGEMA_signal_17025, new_AGEMA_signal_17021, new_AGEMA_signal_17017}), .clk (clk), .Q ({ciphertext_s3[53], ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17045, new_AGEMA_signal_17041, new_AGEMA_signal_17037, new_AGEMA_signal_17033}), .clk (clk), .Q ({ciphertext_s3[54], ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17061, new_AGEMA_signal_17057, new_AGEMA_signal_17053, new_AGEMA_signal_17049}), .clk (clk), .Q ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17077, new_AGEMA_signal_17073, new_AGEMA_signal_17069, new_AGEMA_signal_17065}), .clk (clk), .Q ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17093, new_AGEMA_signal_17089, new_AGEMA_signal_17085, new_AGEMA_signal_17081}), .clk (clk), .Q ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17109, new_AGEMA_signal_17105, new_AGEMA_signal_17101, new_AGEMA_signal_17097}), .clk (clk), .Q ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17125, new_AGEMA_signal_17121, new_AGEMA_signal_17117, new_AGEMA_signal_17113}), .clk (clk), .Q ({ciphertext_s3[91], ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17141, new_AGEMA_signal_17137, new_AGEMA_signal_17133, new_AGEMA_signal_17129}), .clk (clk), .Q ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17157, new_AGEMA_signal_17153, new_AGEMA_signal_17149, new_AGEMA_signal_17145}), .clk (clk), .Q ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17173, new_AGEMA_signal_17169, new_AGEMA_signal_17165, new_AGEMA_signal_17161}), .clk (clk), .Q ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17189, new_AGEMA_signal_17185, new_AGEMA_signal_17181, new_AGEMA_signal_17177}), .clk (clk), .Q ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17205, new_AGEMA_signal_17201, new_AGEMA_signal_17197, new_AGEMA_signal_17193}), .clk (clk), .Q ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17221, new_AGEMA_signal_17217, new_AGEMA_signal_17213, new_AGEMA_signal_17209}), .clk (clk), .Q ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17237, new_AGEMA_signal_17233, new_AGEMA_signal_17229, new_AGEMA_signal_17225}), .clk (clk), .Q ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17253, new_AGEMA_signal_17249, new_AGEMA_signal_17245, new_AGEMA_signal_17241}), .clk (clk), .Q ({ciphertext_s3[3], ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17269, new_AGEMA_signal_17265, new_AGEMA_signal_17261, new_AGEMA_signal_17257}), .clk (clk), .Q ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17285, new_AGEMA_signal_17281, new_AGEMA_signal_17277, new_AGEMA_signal_17273}), .clk (clk), .Q ({ciphertext_s3[5], ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17301, new_AGEMA_signal_17297, new_AGEMA_signal_17293, new_AGEMA_signal_17289}), .clk (clk), .Q ({ciphertext_s3[6], ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17317, new_AGEMA_signal_17313, new_AGEMA_signal_17309, new_AGEMA_signal_17305}), .clk (clk), .Q ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17333, new_AGEMA_signal_17329, new_AGEMA_signal_17325, new_AGEMA_signal_17321}), .clk (clk), .Q ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17349, new_AGEMA_signal_17345, new_AGEMA_signal_17341, new_AGEMA_signal_17337}), .clk (clk), .Q ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17365, new_AGEMA_signal_17361, new_AGEMA_signal_17357, new_AGEMA_signal_17353}), .clk (clk), .Q ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17381, new_AGEMA_signal_17377, new_AGEMA_signal_17373, new_AGEMA_signal_17369}), .clk (clk), .Q ({ciphertext_s3[43], ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17397, new_AGEMA_signal_17393, new_AGEMA_signal_17389, new_AGEMA_signal_17385}), .clk (clk), .Q ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17413, new_AGEMA_signal_17409, new_AGEMA_signal_17405, new_AGEMA_signal_17401}), .clk (clk), .Q ({ciphertext_s3[45], ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17429, new_AGEMA_signal_17425, new_AGEMA_signal_17421, new_AGEMA_signal_17417}), .clk (clk), .Q ({ciphertext_s3[46], ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17445, new_AGEMA_signal_17441, new_AGEMA_signal_17437, new_AGEMA_signal_17433}), .clk (clk), .Q ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17461, new_AGEMA_signal_17457, new_AGEMA_signal_17453, new_AGEMA_signal_17449}), .clk (clk), .Q ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17477, new_AGEMA_signal_17473, new_AGEMA_signal_17469, new_AGEMA_signal_17465}), .clk (clk), .Q ({ciphertext_s3[81], ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17493, new_AGEMA_signal_17489, new_AGEMA_signal_17485, new_AGEMA_signal_17481}), .clk (clk), .Q ({ciphertext_s3[82], ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17509, new_AGEMA_signal_17505, new_AGEMA_signal_17501, new_AGEMA_signal_17497}), .clk (clk), .Q ({ciphertext_s3[83], ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17525, new_AGEMA_signal_17521, new_AGEMA_signal_17517, new_AGEMA_signal_17513}), .clk (clk), .Q ({ciphertext_s3[84], ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17541, new_AGEMA_signal_17537, new_AGEMA_signal_17533, new_AGEMA_signal_17529}), .clk (clk), .Q ({ciphertext_s3[85], ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17557, new_AGEMA_signal_17553, new_AGEMA_signal_17549, new_AGEMA_signal_17545}), .clk (clk), .Q ({ciphertext_s3[86], ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17573, new_AGEMA_signal_17569, new_AGEMA_signal_17565, new_AGEMA_signal_17561}), .clk (clk), .Q ({ciphertext_s3[87], ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17589, new_AGEMA_signal_17585, new_AGEMA_signal_17581, new_AGEMA_signal_17577}), .clk (clk), .Q ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17605, new_AGEMA_signal_17601, new_AGEMA_signal_17597, new_AGEMA_signal_17593}), .clk (clk), .Q ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17621, new_AGEMA_signal_17617, new_AGEMA_signal_17613, new_AGEMA_signal_17609}), .clk (clk), .Q ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17637, new_AGEMA_signal_17633, new_AGEMA_signal_17629, new_AGEMA_signal_17625}), .clk (clk), .Q ({ciphertext_s3[123], ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17653, new_AGEMA_signal_17649, new_AGEMA_signal_17645, new_AGEMA_signal_17641}), .clk (clk), .Q ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17669, new_AGEMA_signal_17665, new_AGEMA_signal_17661, new_AGEMA_signal_17657}), .clk (clk), .Q ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17685, new_AGEMA_signal_17681, new_AGEMA_signal_17677, new_AGEMA_signal_17673}), .clk (clk), .Q ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) RoundReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_17701, new_AGEMA_signal_17697, new_AGEMA_signal_17693, new_AGEMA_signal_17689}), .clk (clk), .Q ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7494, new_AGEMA_signal_7493, new_AGEMA_signal_7492, KeyReg_Inst_ff_SDE_0_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, new_AGEMA_signal_2341, KSSubBytesInput[16]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7950, new_AGEMA_signal_7949, new_AGEMA_signal_7948, KeyReg_Inst_ff_SDE_1_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2694, new_AGEMA_signal_2693, new_AGEMA_signal_2692, KSSubBytesInput[17]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7956, new_AGEMA_signal_7955, new_AGEMA_signal_7954, KeyReg_Inst_ff_SDE_2_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, new_AGEMA_signal_2791, KSSubBytesInput[18]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, new_AGEMA_signal_7960, KeyReg_Inst_ff_SDE_3_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2892, new_AGEMA_signal_2891, new_AGEMA_signal_2890, KSSubBytesInput[19]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7968, new_AGEMA_signal_7967, new_AGEMA_signal_7966, KeyReg_Inst_ff_SDE_4_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, new_AGEMA_signal_2989, KSSubBytesInput[20]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7974, new_AGEMA_signal_7973, new_AGEMA_signal_7972, KeyReg_Inst_ff_SDE_5_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3090, new_AGEMA_signal_3089, new_AGEMA_signal_3088, KSSubBytesInput[21]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7980, new_AGEMA_signal_7979, new_AGEMA_signal_7978, KeyReg_Inst_ff_SDE_6_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, new_AGEMA_signal_3187, KSSubBytesInput[22]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7986, new_AGEMA_signal_7985, new_AGEMA_signal_7984, KeyReg_Inst_ff_SDE_7_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3288, new_AGEMA_signal_3287, new_AGEMA_signal_3286, KSSubBytesInput[23]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7500, new_AGEMA_signal_7499, new_AGEMA_signal_7498, KeyReg_Inst_ff_SDE_8_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, new_AGEMA_signal_3385, KSSubBytesInput[8]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7992, new_AGEMA_signal_7991, new_AGEMA_signal_7990, KeyReg_Inst_ff_SDE_9_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3486, new_AGEMA_signal_3485, new_AGEMA_signal_3484, KSSubBytesInput[9]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7998, new_AGEMA_signal_7997, new_AGEMA_signal_7996, KeyReg_Inst_ff_SDE_10_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2442, new_AGEMA_signal_2441, new_AGEMA_signal_2440, KSSubBytesInput[10]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8004, new_AGEMA_signal_8003, new_AGEMA_signal_8002, KeyReg_Inst_ff_SDE_11_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, new_AGEMA_signal_2539, KSSubBytesInput[11]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8010, new_AGEMA_signal_8009, new_AGEMA_signal_8008, KeyReg_Inst_ff_SDE_12_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2622, new_AGEMA_signal_2621, new_AGEMA_signal_2620, KSSubBytesInput[12]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8016, new_AGEMA_signal_8015, new_AGEMA_signal_8014, KeyReg_Inst_ff_SDE_13_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, new_AGEMA_signal_2629, KSSubBytesInput[13]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8022, new_AGEMA_signal_8021, new_AGEMA_signal_8020, KeyReg_Inst_ff_SDE_14_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2640, new_AGEMA_signal_2639, new_AGEMA_signal_2638, KSSubBytesInput[14]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8028, new_AGEMA_signal_8027, new_AGEMA_signal_8026, KeyReg_Inst_ff_SDE_15_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, new_AGEMA_signal_2647, KSSubBytesInput[15]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7506, new_AGEMA_signal_7505, new_AGEMA_signal_7504, KeyReg_Inst_ff_SDE_16_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2658, new_AGEMA_signal_2657, new_AGEMA_signal_2656, KSSubBytesInput[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8034, new_AGEMA_signal_8033, new_AGEMA_signal_8032, KeyReg_Inst_ff_SDE_17_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, new_AGEMA_signal_2665, KSSubBytesInput[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8040, new_AGEMA_signal_8039, new_AGEMA_signal_8038, KeyReg_Inst_ff_SDE_18_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2676, new_AGEMA_signal_2675, new_AGEMA_signal_2674, KSSubBytesInput[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8046, new_AGEMA_signal_8045, new_AGEMA_signal_8044, KeyReg_Inst_ff_SDE_19_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, new_AGEMA_signal_2683, KSSubBytesInput[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8052, new_AGEMA_signal_8051, new_AGEMA_signal_8050, KeyReg_Inst_ff_SDE_20_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, new_AGEMA_signal_2701, KSSubBytesInput[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8058, new_AGEMA_signal_8057, new_AGEMA_signal_8056, KeyReg_Inst_ff_SDE_21_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2712, new_AGEMA_signal_2711, new_AGEMA_signal_2710, KSSubBytesInput[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8064, new_AGEMA_signal_8063, new_AGEMA_signal_8062, KeyReg_Inst_ff_SDE_22_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, new_AGEMA_signal_2719, KSSubBytesInput[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8070, new_AGEMA_signal_8069, new_AGEMA_signal_8068, KeyReg_Inst_ff_SDE_23_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2730, new_AGEMA_signal_2729, new_AGEMA_signal_2728, KSSubBytesInput[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8076, new_AGEMA_signal_8075, new_AGEMA_signal_8074, KeyReg_Inst_ff_SDE_24_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, new_AGEMA_signal_2737, KSSubBytesInput[24]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8217, new_AGEMA_signal_8216, new_AGEMA_signal_8215, KeyReg_Inst_ff_SDE_25_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2748, new_AGEMA_signal_2747, new_AGEMA_signal_2746, KSSubBytesInput[25]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8223, new_AGEMA_signal_8222, new_AGEMA_signal_8221, KeyReg_Inst_ff_SDE_26_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, new_AGEMA_signal_2755, KSSubBytesInput[26]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8229, new_AGEMA_signal_8228, new_AGEMA_signal_8227, KeyReg_Inst_ff_SDE_27_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2766, new_AGEMA_signal_2765, new_AGEMA_signal_2764, KSSubBytesInput[27]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8235, new_AGEMA_signal_8234, new_AGEMA_signal_8233, KeyReg_Inst_ff_SDE_28_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, new_AGEMA_signal_2773, KSSubBytesInput[28]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8241, new_AGEMA_signal_8240, new_AGEMA_signal_8239, KeyReg_Inst_ff_SDE_29_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2784, new_AGEMA_signal_2783, new_AGEMA_signal_2782, KSSubBytesInput[29]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8247, new_AGEMA_signal_8246, new_AGEMA_signal_8245, KeyReg_Inst_ff_SDE_30_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2802, new_AGEMA_signal_2801, new_AGEMA_signal_2800, KSSubBytesInput[30]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8253, new_AGEMA_signal_8252, new_AGEMA_signal_8251, KeyReg_Inst_ff_SDE_31_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, new_AGEMA_signal_2809, KSSubBytesInput[31]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7023, new_AGEMA_signal_7022, new_AGEMA_signal_7021, KeyReg_Inst_ff_SDE_32_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2820, new_AGEMA_signal_2819, new_AGEMA_signal_2818, RoundKey[32]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7512, new_AGEMA_signal_7511, new_AGEMA_signal_7510, KeyReg_Inst_ff_SDE_33_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, new_AGEMA_signal_2827, RoundKey[33]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7518, new_AGEMA_signal_7517, new_AGEMA_signal_7516, KeyReg_Inst_ff_SDE_34_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2838, new_AGEMA_signal_2837, new_AGEMA_signal_2836, RoundKey[34]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7524, new_AGEMA_signal_7523, new_AGEMA_signal_7522, KeyReg_Inst_ff_SDE_35_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, new_AGEMA_signal_2845, RoundKey[35]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7530, new_AGEMA_signal_7529, new_AGEMA_signal_7528, KeyReg_Inst_ff_SDE_36_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2856, new_AGEMA_signal_2855, new_AGEMA_signal_2854, RoundKey[36]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7536, new_AGEMA_signal_7535, new_AGEMA_signal_7534, KeyReg_Inst_ff_SDE_37_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, new_AGEMA_signal_2863, RoundKey[37]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7542, new_AGEMA_signal_7541, new_AGEMA_signal_7540, KeyReg_Inst_ff_SDE_38_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2874, new_AGEMA_signal_2873, new_AGEMA_signal_2872, RoundKey[38]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7548, new_AGEMA_signal_7547, new_AGEMA_signal_7546, KeyReg_Inst_ff_SDE_39_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, new_AGEMA_signal_2881, RoundKey[39]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7029, new_AGEMA_signal_7028, new_AGEMA_signal_7027, KeyReg_Inst_ff_SDE_40_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, new_AGEMA_signal_2899, RoundKey[40]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7554, new_AGEMA_signal_7553, new_AGEMA_signal_7552, KeyReg_Inst_ff_SDE_41_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2910, new_AGEMA_signal_2909, new_AGEMA_signal_2908, RoundKey[41]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7560, new_AGEMA_signal_7559, new_AGEMA_signal_7558, KeyReg_Inst_ff_SDE_42_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, new_AGEMA_signal_2917, RoundKey[42]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7566, new_AGEMA_signal_7565, new_AGEMA_signal_7564, KeyReg_Inst_ff_SDE_43_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2928, new_AGEMA_signal_2927, new_AGEMA_signal_2926, RoundKey[43]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7572, new_AGEMA_signal_7571, new_AGEMA_signal_7570, KeyReg_Inst_ff_SDE_44_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, new_AGEMA_signal_2935, RoundKey[44]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7578, new_AGEMA_signal_7577, new_AGEMA_signal_7576, KeyReg_Inst_ff_SDE_45_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2946, new_AGEMA_signal_2945, new_AGEMA_signal_2944, RoundKey[45]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7584, new_AGEMA_signal_7583, new_AGEMA_signal_7582, KeyReg_Inst_ff_SDE_46_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, new_AGEMA_signal_2953, RoundKey[46]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7590, new_AGEMA_signal_7589, new_AGEMA_signal_7588, KeyReg_Inst_ff_SDE_47_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2964, new_AGEMA_signal_2963, new_AGEMA_signal_2962, RoundKey[47]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7035, new_AGEMA_signal_7034, new_AGEMA_signal_7033, KeyReg_Inst_ff_SDE_48_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, new_AGEMA_signal_2971, RoundKey[48]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7596, new_AGEMA_signal_7595, new_AGEMA_signal_7594, KeyReg_Inst_ff_SDE_49_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2982, new_AGEMA_signal_2981, new_AGEMA_signal_2980, RoundKey[49]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7602, new_AGEMA_signal_7601, new_AGEMA_signal_7600, KeyReg_Inst_ff_SDE_50_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3000, new_AGEMA_signal_2999, new_AGEMA_signal_2998, RoundKey[50]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7608, new_AGEMA_signal_7607, new_AGEMA_signal_7606, KeyReg_Inst_ff_SDE_51_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, new_AGEMA_signal_3007, RoundKey[51]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7614, new_AGEMA_signal_7613, new_AGEMA_signal_7612, KeyReg_Inst_ff_SDE_52_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3018, new_AGEMA_signal_3017, new_AGEMA_signal_3016, RoundKey[52]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7620, new_AGEMA_signal_7619, new_AGEMA_signal_7618, KeyReg_Inst_ff_SDE_53_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, new_AGEMA_signal_3025, RoundKey[53]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7626, new_AGEMA_signal_7625, new_AGEMA_signal_7624, KeyReg_Inst_ff_SDE_54_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3036, new_AGEMA_signal_3035, new_AGEMA_signal_3034, RoundKey[54]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7632, new_AGEMA_signal_7631, new_AGEMA_signal_7630, KeyReg_Inst_ff_SDE_55_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, new_AGEMA_signal_3043, RoundKey[55]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7638, new_AGEMA_signal_7637, new_AGEMA_signal_7636, KeyReg_Inst_ff_SDE_56_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3054, new_AGEMA_signal_3053, new_AGEMA_signal_3052, RoundKey[56]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8082, new_AGEMA_signal_8081, new_AGEMA_signal_8080, KeyReg_Inst_ff_SDE_57_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, new_AGEMA_signal_3061, RoundKey[57]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8088, new_AGEMA_signal_8087, new_AGEMA_signal_8086, KeyReg_Inst_ff_SDE_58_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3072, new_AGEMA_signal_3071, new_AGEMA_signal_3070, RoundKey[58]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8094, new_AGEMA_signal_8093, new_AGEMA_signal_8092, KeyReg_Inst_ff_SDE_59_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, new_AGEMA_signal_3079, RoundKey[59]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8100, new_AGEMA_signal_8099, new_AGEMA_signal_8098, KeyReg_Inst_ff_SDE_60_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, new_AGEMA_signal_3097, RoundKey[60]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8106, new_AGEMA_signal_8105, new_AGEMA_signal_8104, KeyReg_Inst_ff_SDE_61_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3108, new_AGEMA_signal_3107, new_AGEMA_signal_3106, RoundKey[61]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8112, new_AGEMA_signal_8111, new_AGEMA_signal_8110, KeyReg_Inst_ff_SDE_62_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, new_AGEMA_signal_3115, RoundKey[62]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8118, new_AGEMA_signal_8117, new_AGEMA_signal_8116, KeyReg_Inst_ff_SDE_63_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3126, new_AGEMA_signal_3125, new_AGEMA_signal_3124, RoundKey[63]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6585, new_AGEMA_signal_6584, new_AGEMA_signal_6583, KeyReg_Inst_ff_SDE_64_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, new_AGEMA_signal_3133, RoundKey[64]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7041, new_AGEMA_signal_7040, new_AGEMA_signal_7039, KeyReg_Inst_ff_SDE_65_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3144, new_AGEMA_signal_3143, new_AGEMA_signal_3142, RoundKey[65]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7047, new_AGEMA_signal_7046, new_AGEMA_signal_7045, KeyReg_Inst_ff_SDE_66_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, new_AGEMA_signal_3151, RoundKey[66]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7053, new_AGEMA_signal_7052, new_AGEMA_signal_7051, KeyReg_Inst_ff_SDE_67_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3162, new_AGEMA_signal_3161, new_AGEMA_signal_3160, RoundKey[67]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7059, new_AGEMA_signal_7058, new_AGEMA_signal_7057, KeyReg_Inst_ff_SDE_68_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, new_AGEMA_signal_3169, RoundKey[68]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7065, new_AGEMA_signal_7064, new_AGEMA_signal_7063, KeyReg_Inst_ff_SDE_69_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3180, new_AGEMA_signal_3179, new_AGEMA_signal_3178, RoundKey[69]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7071, new_AGEMA_signal_7070, new_AGEMA_signal_7069, KeyReg_Inst_ff_SDE_70_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3198, new_AGEMA_signal_3197, new_AGEMA_signal_3196, RoundKey[70]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7077, new_AGEMA_signal_7076, new_AGEMA_signal_7075, KeyReg_Inst_ff_SDE_71_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, new_AGEMA_signal_3205, RoundKey[71]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6591, new_AGEMA_signal_6590, new_AGEMA_signal_6589, KeyReg_Inst_ff_SDE_72_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3216, new_AGEMA_signal_3215, new_AGEMA_signal_3214, RoundKey[72]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7083, new_AGEMA_signal_7082, new_AGEMA_signal_7081, KeyReg_Inst_ff_SDE_73_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, new_AGEMA_signal_3223, RoundKey[73]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7089, new_AGEMA_signal_7088, new_AGEMA_signal_7087, KeyReg_Inst_ff_SDE_74_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3234, new_AGEMA_signal_3233, new_AGEMA_signal_3232, RoundKey[74]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7095, new_AGEMA_signal_7094, new_AGEMA_signal_7093, KeyReg_Inst_ff_SDE_75_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, new_AGEMA_signal_3241, RoundKey[75]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7101, new_AGEMA_signal_7100, new_AGEMA_signal_7099, KeyReg_Inst_ff_SDE_76_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3252, new_AGEMA_signal_3251, new_AGEMA_signal_3250, RoundKey[76]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7107, new_AGEMA_signal_7106, new_AGEMA_signal_7105, KeyReg_Inst_ff_SDE_77_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, new_AGEMA_signal_3259, RoundKey[77]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7113, new_AGEMA_signal_7112, new_AGEMA_signal_7111, KeyReg_Inst_ff_SDE_78_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3270, new_AGEMA_signal_3269, new_AGEMA_signal_3268, RoundKey[78]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7119, new_AGEMA_signal_7118, new_AGEMA_signal_7117, KeyReg_Inst_ff_SDE_79_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, new_AGEMA_signal_3277, RoundKey[79]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6597, new_AGEMA_signal_6596, new_AGEMA_signal_6595, KeyReg_Inst_ff_SDE_80_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, new_AGEMA_signal_3295, RoundKey[80]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7125, new_AGEMA_signal_7124, new_AGEMA_signal_7123, KeyReg_Inst_ff_SDE_81_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3306, new_AGEMA_signal_3305, new_AGEMA_signal_3304, RoundKey[81]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7131, new_AGEMA_signal_7130, new_AGEMA_signal_7129, KeyReg_Inst_ff_SDE_82_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, new_AGEMA_signal_3313, RoundKey[82]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7137, new_AGEMA_signal_7136, new_AGEMA_signal_7135, KeyReg_Inst_ff_SDE_83_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3324, new_AGEMA_signal_3323, new_AGEMA_signal_3322, RoundKey[83]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7143, new_AGEMA_signal_7142, new_AGEMA_signal_7141, KeyReg_Inst_ff_SDE_84_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, new_AGEMA_signal_3331, RoundKey[84]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7149, new_AGEMA_signal_7148, new_AGEMA_signal_7147, KeyReg_Inst_ff_SDE_85_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3342, new_AGEMA_signal_3341, new_AGEMA_signal_3340, RoundKey[85]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7155, new_AGEMA_signal_7154, new_AGEMA_signal_7153, KeyReg_Inst_ff_SDE_86_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, new_AGEMA_signal_3349, RoundKey[86]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7161, new_AGEMA_signal_7160, new_AGEMA_signal_7159, KeyReg_Inst_ff_SDE_87_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3360, new_AGEMA_signal_3359, new_AGEMA_signal_3358, RoundKey[87]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7167, new_AGEMA_signal_7166, new_AGEMA_signal_7165, KeyReg_Inst_ff_SDE_88_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, new_AGEMA_signal_3367, RoundKey[88]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7644, new_AGEMA_signal_7643, new_AGEMA_signal_7642, KeyReg_Inst_ff_SDE_89_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3378, new_AGEMA_signal_3377, new_AGEMA_signal_3376, RoundKey[89]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7650, new_AGEMA_signal_7649, new_AGEMA_signal_7648, KeyReg_Inst_ff_SDE_90_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3396, new_AGEMA_signal_3395, new_AGEMA_signal_3394, RoundKey[90]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7656, new_AGEMA_signal_7655, new_AGEMA_signal_7654, KeyReg_Inst_ff_SDE_91_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, new_AGEMA_signal_3403, RoundKey[91]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7662, new_AGEMA_signal_7661, new_AGEMA_signal_7660, KeyReg_Inst_ff_SDE_92_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3414, new_AGEMA_signal_3413, new_AGEMA_signal_3412, RoundKey[92]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7668, new_AGEMA_signal_7667, new_AGEMA_signal_7666, KeyReg_Inst_ff_SDE_93_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, new_AGEMA_signal_3421, RoundKey[93]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7674, new_AGEMA_signal_7673, new_AGEMA_signal_7672, KeyReg_Inst_ff_SDE_94_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3432, new_AGEMA_signal_3431, new_AGEMA_signal_3430, RoundKey[94]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7680, new_AGEMA_signal_7679, new_AGEMA_signal_7678, KeyReg_Inst_ff_SDE_95_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, new_AGEMA_signal_3439, RoundKey[95]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6300, new_AGEMA_signal_6299, new_AGEMA_signal_6298, KeyReg_Inst_ff_SDE_96_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3450, new_AGEMA_signal_3449, new_AGEMA_signal_3448, RoundKey[96]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6603, new_AGEMA_signal_6602, new_AGEMA_signal_6601, KeyReg_Inst_ff_SDE_97_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, new_AGEMA_signal_3457, RoundKey[97]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6609, new_AGEMA_signal_6608, new_AGEMA_signal_6607, KeyReg_Inst_ff_SDE_98_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3468, new_AGEMA_signal_3467, new_AGEMA_signal_3466, RoundKey[98]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6615, new_AGEMA_signal_6614, new_AGEMA_signal_6613, KeyReg_Inst_ff_SDE_99_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, new_AGEMA_signal_3475, RoundKey[99]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6621, new_AGEMA_signal_6620, new_AGEMA_signal_6619, KeyReg_Inst_ff_SDE_100_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2352, new_AGEMA_signal_2351, new_AGEMA_signal_2350, RoundKey[100]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6627, new_AGEMA_signal_6626, new_AGEMA_signal_6625, KeyReg_Inst_ff_SDE_101_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, new_AGEMA_signal_2359, RoundKey[101]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6633, new_AGEMA_signal_6632, new_AGEMA_signal_6631, KeyReg_Inst_ff_SDE_102_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2370, new_AGEMA_signal_2369, new_AGEMA_signal_2368, RoundKey[102]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6639, new_AGEMA_signal_6638, new_AGEMA_signal_6637, KeyReg_Inst_ff_SDE_103_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, new_AGEMA_signal_2377, RoundKey[103]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6306, new_AGEMA_signal_6305, new_AGEMA_signal_6304, KeyReg_Inst_ff_SDE_104_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2388, new_AGEMA_signal_2387, new_AGEMA_signal_2386, RoundKey[104]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6645, new_AGEMA_signal_6644, new_AGEMA_signal_6643, KeyReg_Inst_ff_SDE_105_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, new_AGEMA_signal_2395, RoundKey[105]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6651, new_AGEMA_signal_6650, new_AGEMA_signal_6649, KeyReg_Inst_ff_SDE_106_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2406, new_AGEMA_signal_2405, new_AGEMA_signal_2404, RoundKey[106]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6657, new_AGEMA_signal_6656, new_AGEMA_signal_6655, KeyReg_Inst_ff_SDE_107_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, new_AGEMA_signal_2413, RoundKey[107]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6663, new_AGEMA_signal_6662, new_AGEMA_signal_6661, KeyReg_Inst_ff_SDE_108_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2424, new_AGEMA_signal_2423, new_AGEMA_signal_2422, RoundKey[108]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6669, new_AGEMA_signal_6668, new_AGEMA_signal_6667, KeyReg_Inst_ff_SDE_109_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, new_AGEMA_signal_2431, RoundKey[109]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6675, new_AGEMA_signal_6674, new_AGEMA_signal_6673, KeyReg_Inst_ff_SDE_110_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, new_AGEMA_signal_2449, RoundKey[110]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6681, new_AGEMA_signal_6680, new_AGEMA_signal_6679, KeyReg_Inst_ff_SDE_111_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2460, new_AGEMA_signal_2459, new_AGEMA_signal_2458, RoundKey[111]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6312, new_AGEMA_signal_6311, new_AGEMA_signal_6310, KeyReg_Inst_ff_SDE_112_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, new_AGEMA_signal_2467, RoundKey[112]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6687, new_AGEMA_signal_6686, new_AGEMA_signal_6685, KeyReg_Inst_ff_SDE_113_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2478, new_AGEMA_signal_2477, new_AGEMA_signal_2476, RoundKey[113]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6693, new_AGEMA_signal_6692, new_AGEMA_signal_6691, KeyReg_Inst_ff_SDE_114_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, new_AGEMA_signal_2485, RoundKey[114]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6699, new_AGEMA_signal_6698, new_AGEMA_signal_6697, KeyReg_Inst_ff_SDE_115_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2496, new_AGEMA_signal_2495, new_AGEMA_signal_2494, RoundKey[115]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6705, new_AGEMA_signal_6704, new_AGEMA_signal_6703, KeyReg_Inst_ff_SDE_116_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, new_AGEMA_signal_2503, RoundKey[116]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6711, new_AGEMA_signal_6710, new_AGEMA_signal_6709, KeyReg_Inst_ff_SDE_117_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2514, new_AGEMA_signal_2513, new_AGEMA_signal_2512, RoundKey[117]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6717, new_AGEMA_signal_6716, new_AGEMA_signal_6715, KeyReg_Inst_ff_SDE_118_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, new_AGEMA_signal_2521, RoundKey[118]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6723, new_AGEMA_signal_6722, new_AGEMA_signal_6721, KeyReg_Inst_ff_SDE_119_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2532, new_AGEMA_signal_2531, new_AGEMA_signal_2530, RoundKey[119]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6729, new_AGEMA_signal_6728, new_AGEMA_signal_6727, KeyReg_Inst_ff_SDE_120_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2550, new_AGEMA_signal_2549, new_AGEMA_signal_2548, RoundKey[120]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7173, new_AGEMA_signal_7172, new_AGEMA_signal_7171, KeyReg_Inst_ff_SDE_121_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, new_AGEMA_signal_2557, RoundKey[121]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7179, new_AGEMA_signal_7178, new_AGEMA_signal_7177, KeyReg_Inst_ff_SDE_122_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2568, new_AGEMA_signal_2567, new_AGEMA_signal_2566, RoundKey[122]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7185, new_AGEMA_signal_7184, new_AGEMA_signal_7183, KeyReg_Inst_ff_SDE_123_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, new_AGEMA_signal_2575, RoundKey[123]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7191, new_AGEMA_signal_7190, new_AGEMA_signal_7189, KeyReg_Inst_ff_SDE_124_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2586, new_AGEMA_signal_2585, new_AGEMA_signal_2584, RoundKey[124]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7197, new_AGEMA_signal_7196, new_AGEMA_signal_7195, KeyReg_Inst_ff_SDE_125_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, new_AGEMA_signal_2593, RoundKey[125]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7203, new_AGEMA_signal_7202, new_AGEMA_signal_7201, KeyReg_Inst_ff_SDE_126_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2604, new_AGEMA_signal_2603, new_AGEMA_signal_2602, RoundKey[126]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) KeyReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7209, new_AGEMA_signal_7208, new_AGEMA_signal_7207, KeyReg_Inst_ff_SDE_127_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, new_AGEMA_signal_2611, RoundKey[127]}) ) ;
    DFF_X1 RoundCounterIns_count_reg_0__FF_FF ( .D (new_AGEMA_signal_17705), .CK (clk), .Q (RoundCounter[0]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_1__FF_FF ( .D (new_AGEMA_signal_17709), .CK (clk), .Q (RoundCounter[1]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_2__FF_FF ( .D (new_AGEMA_signal_17713), .CK (clk), .Q (RoundCounter[2]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_3__FF_FF ( .D (new_AGEMA_signal_17717), .CK (clk), .Q (RoundCounter[3]), .QN () ) ;
    DFF_X1 InRoundCounterIns_count_reg_0__FF_FF ( .D (new_AGEMA_signal_17721), .CK (clk), .Q (InRoundCounter[0]), .QN () ) ;
    DFF_X1 InRoundCounterIns_count_reg_1__FF_FF ( .D (new_AGEMA_signal_17725), .CK (clk), .Q (InRoundCounter[1]), .QN () ) ;
    DFF_X1 InRoundCounterIns_count_reg_2__FF_FF ( .D (new_AGEMA_signal_17729), .CK (clk), .Q (InRoundCounter[2]), .QN () ) ;
endmodule
