module Reg1(x, y);
 input [135:0] x;
 output [134:0] y;

  assign y[0] = x[135];
  register_stage #(.WIDTH(134)) inst_0(.clk(x[134]), .D({x[0],x[1],x[2],x[3],x[4],x[5],x[6],x[17],x[28],x[39],x[50],x[61],x[66],x[67],x[68],x[69],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[18],x[19],x[20],x[21],x[22],x[23],x[24],x[25],x[26],x[27],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[40],x[41],x[42],x[43],x[44],x[45],x[46],x[47],x[48],x[49],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[62],x[63],x[64],x[65],x[70],x[81],x[92],x[103],x[114],x[125],x[130],x[131],x[132],x[133],x[71],x[72],x[73],x[74],x[75],x[76],x[77],x[78],x[79],x[80],x[82],x[83],x[84],x[85],x[86],x[87],x[88],x[89],x[90],x[91],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[104],x[105],x[106],x[107],x[108],x[109],x[110],x[111],x[112],x[113],x[115],x[116],x[117],x[118],x[119],x[120],x[121],x[122],x[123],x[124],x[126],x[127],x[128],x[129]}), .Q({y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134]}));
endmodule

module Reg2(x, y);
 input [540:0] x;
 output [539:0] y;

  assign y[0] = x[537];
  assign y[1] = x[538];
  assign y[2] = x[539];
  assign y[3] = x[540];
  register_stage #(.WIDTH(536)) inst_0(.clk(x[536]), .D({x[0],x[1],x[2],x[3],x[4],x[5],x[6],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[22],x[23],x[24],x[25],x[26],x[27],x[68],x[69],x[70],x[71],x[112],x[113],x[114],x[115],x[156],x[157],x[158],x[159],x[200],x[201],x[202],x[203],x[244],x[245],x[246],x[247],x[264],x[265],x[266],x[267],x[268],x[269],x[270],x[271],x[272],x[273],x[274],x[275],x[276],x[277],x[278],x[279],x[28],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[44],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[61],x[62],x[63],x[64],x[65],x[66],x[67],x[72],x[73],x[74],x[75],x[76],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[84],x[85],x[86],x[87],x[88],x[89],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[103],x[104],x[105],x[106],x[107],x[108],x[109],x[110],x[111],x[116],x[117],x[118],x[119],x[120],x[121],x[122],x[123],x[124],x[125],x[126],x[127],x[128],x[129],x[130],x[131],x[132],x[133],x[134],x[135],x[136],x[137],x[138],x[139],x[140],x[141],x[142],x[143],x[144],x[145],x[146],x[147],x[148],x[149],x[150],x[151],x[152],x[153],x[154],x[155],x[160],x[161],x[162],x[163],x[164],x[165],x[166],x[167],x[168],x[169],x[170],x[171],x[172],x[173],x[174],x[175],x[176],x[177],x[178],x[179],x[180],x[181],x[182],x[183],x[184],x[185],x[186],x[187],x[188],x[189],x[190],x[191],x[192],x[193],x[194],x[195],x[196],x[197],x[198],x[199],x[204],x[205],x[206],x[207],x[208],x[209],x[210],x[211],x[212],x[213],x[214],x[215],x[216],x[217],x[218],x[219],x[220],x[221],x[222],x[223],x[224],x[225],x[226],x[227],x[228],x[229],x[230],x[231],x[232],x[233],x[234],x[235],x[236],x[237],x[238],x[239],x[240],x[241],x[242],x[243],x[248],x[249],x[250],x[251],x[252],x[253],x[254],x[255],x[256],x[257],x[258],x[259],x[260],x[261],x[262],x[263],x[280],x[281],x[282],x[283],x[324],x[325],x[326],x[327],x[368],x[369],x[370],x[371],x[412],x[413],x[414],x[415],x[456],x[457],x[458],x[459],x[500],x[501],x[502],x[503],x[520],x[521],x[522],x[523],x[524],x[525],x[526],x[527],x[528],x[529],x[530],x[531],x[532],x[533],x[534],x[535],x[284],x[285],x[286],x[287],x[288],x[289],x[290],x[291],x[292],x[293],x[294],x[295],x[296],x[297],x[298],x[299],x[300],x[301],x[302],x[303],x[304],x[305],x[306],x[307],x[308],x[309],x[310],x[311],x[312],x[313],x[314],x[315],x[316],x[317],x[318],x[319],x[320],x[321],x[322],x[323],x[328],x[329],x[330],x[331],x[332],x[333],x[334],x[335],x[336],x[337],x[338],x[339],x[340],x[341],x[342],x[343],x[344],x[345],x[346],x[347],x[348],x[349],x[350],x[351],x[352],x[353],x[354],x[355],x[356],x[357],x[358],x[359],x[360],x[361],x[362],x[363],x[364],x[365],x[366],x[367],x[372],x[373],x[374],x[375],x[376],x[377],x[378],x[379],x[380],x[381],x[382],x[383],x[384],x[385],x[386],x[387],x[388],x[389],x[390],x[391],x[392],x[393],x[394],x[395],x[396],x[397],x[398],x[399],x[400],x[401],x[402],x[403],x[404],x[405],x[406],x[407],x[408],x[409],x[410],x[411],x[416],x[417],x[418],x[419],x[420],x[421],x[422],x[423],x[424],x[425],x[426],x[427],x[428],x[429],x[430],x[431],x[432],x[433],x[434],x[435],x[436],x[437],x[438],x[439],x[440],x[441],x[442],x[443],x[444],x[445],x[446],x[447],x[448],x[449],x[450],x[451],x[452],x[453],x[454],x[455],x[460],x[461],x[462],x[463],x[464],x[465],x[466],x[467],x[468],x[469],x[470],x[471],x[472],x[473],x[474],x[475],x[476],x[477],x[478],x[479],x[480],x[481],x[482],x[483],x[484],x[485],x[486],x[487],x[488],x[489],x[490],x[491],x[492],x[493],x[494],x[495],x[496],x[497],x[498],x[499],x[504],x[505],x[506],x[507],x[508],x[509],x[510],x[511],x[512],x[513],x[514],x[515],x[516],x[517],x[518],x[519]}), .Q({y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149],y[150],y[151],y[152],y[153],y[154],y[155],y[156],y[157],y[158],y[159],y[160],y[161],y[162],y[163],y[164],y[165],y[166],y[167],y[168],y[169],y[170],y[171],y[172],y[173],y[174],y[175],y[176],y[177],y[178],y[179],y[180],y[181],y[182],y[183],y[184],y[185],y[186],y[187],y[188],y[189],y[190],y[191],y[192],y[193],y[194],y[195],y[196],y[197],y[198],y[199],y[200],y[201],y[202],y[203],y[204],y[205],y[206],y[207],y[208],y[209],y[210],y[211],y[212],y[213],y[214],y[215],y[216],y[217],y[218],y[219],y[220],y[221],y[222],y[223],y[224],y[225],y[226],y[227],y[228],y[229],y[230],y[231],y[232],y[233],y[234],y[235],y[236],y[237],y[238],y[239],y[240],y[241],y[242],y[243],y[244],y[245],y[246],y[247],y[248],y[249],y[250],y[251],y[252],y[253],y[254],y[255],y[256],y[257],y[258],y[259],y[260],y[261],y[262],y[263],y[264],y[265],y[266],y[267],y[268],y[269],y[270],y[271],y[272],y[273],y[274],y[275],y[276],y[277],y[278],y[279],y[280],y[281],y[282],y[283],y[284],y[285],y[286],y[287],y[288],y[289],y[290],y[291],y[292],y[293],y[294],y[295],y[296],y[297],y[298],y[299],y[300],y[301],y[302],y[303],y[304],y[305],y[306],y[307],y[308],y[309],y[310],y[311],y[312],y[313],y[314],y[315],y[316],y[317],y[318],y[319],y[320],y[321],y[322],y[323],y[324],y[325],y[326],y[327],y[328],y[329],y[330],y[331],y[332],y[333],y[334],y[335],y[336],y[337],y[338],y[339],y[340],y[341],y[342],y[343],y[344],y[345],y[346],y[347],y[348],y[349],y[350],y[351],y[352],y[353],y[354],y[355],y[356],y[357],y[358],y[359],y[360],y[361],y[362],y[363],y[364],y[365],y[366],y[367],y[368],y[369],y[370],y[371],y[372],y[373],y[374],y[375],y[376],y[377],y[378],y[379],y[380],y[381],y[382],y[383],y[384],y[385],y[386],y[387],y[388],y[389],y[390],y[391],y[392],y[393],y[394],y[395],y[396],y[397],y[398],y[399],y[400],y[401],y[402],y[403],y[404],y[405],y[406],y[407],y[408],y[409],y[410],y[411],y[412],y[413],y[414],y[415],y[416],y[417],y[418],y[419],y[420],y[421],y[422],y[423],y[424],y[425],y[426],y[427],y[428],y[429],y[430],y[431],y[432],y[433],y[434],y[435],y[436],y[437],y[438],y[439],y[440],y[441],y[442],y[443],y[444],y[445],y[446],y[447],y[448],y[449],y[450],y[451],y[452],y[453],y[454],y[455],y[456],y[457],y[458],y[459],y[460],y[461],y[462],y[463],y[464],y[465],y[466],y[467],y[468],y[469],y[470],y[471],y[472],y[473],y[474],y[475],y[476],y[477],y[478],y[479],y[480],y[481],y[482],y[483],y[484],y[485],y[486],y[487],y[488],y[489],y[490],y[491],y[492],y[493],y[494],y[495],y[496],y[497],y[498],y[499],y[500],y[501],y[502],y[503],y[504],y[505],y[506],y[507],y[508],y[509],y[510],y[511],y[512],y[513],y[514],y[515],y[516],y[517],y[518],y[519],y[520],y[521],y[522],y[523],y[524],y[525],y[526],y[527],y[528],y[529],y[530],y[531],y[532],y[533],y[534],y[535],y[536],y[537],y[538],y[539]}));
endmodule

module Fx0(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx1(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx2(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx3(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx4(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx5(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx6(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx7(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx8(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx9(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx10(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx11(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx12(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx13(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx14(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx15(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx16(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx17(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx18(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx19(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx20(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx21(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx22(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx23(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx24(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx25(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx26(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx27(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx28(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx29(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx30(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx31(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx32(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx33(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx34(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx35(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx36(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx37(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx38(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx39(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx40(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx41(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx42(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx43(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx44(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx45(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx46(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx47(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx48(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx49(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx50(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx51(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx52(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx53(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx54(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx55(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx56(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx57(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx58(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx59(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx60(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx61(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx62(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx63(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx64(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx65(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx66(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx67(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx68(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx69(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx70(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx71(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx72(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx73(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx74(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx75(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx76(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx77(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx78(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx79(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx80(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx81(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx82(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx83(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx84(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx85(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx86(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx87(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx88(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx89(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx90(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx91(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx92(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx93(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx94(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx95(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx96(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx97(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx98(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx99(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx100(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx101(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx102(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx103(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx104(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx105(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx106(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx107(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx108(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx109(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx110(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx111(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx112(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx113(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx114(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx115(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx116(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx117(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx118(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx119(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx120(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx121(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx122(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx123(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx124(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx125(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx126(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx127(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx128(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx129(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx130(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx131(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx132(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx133(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx134(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx135(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx136(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx137(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx138(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx139(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx140(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx141(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx142(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx143(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx144(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx145(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx146(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx147(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx148(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx149(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx150(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx151(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx152(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx153(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx154(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx155(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx156(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx157(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx158(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx159(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx160(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx161(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx162(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx163(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx164(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx165(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx166(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx167(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx168(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx169(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx170(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx171(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx172(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx173(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx174(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx175(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx176(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx177(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx178(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx179(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx180(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx181(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx182(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx183(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx184(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx185(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx186(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx187(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx188(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx189(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx190(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx191(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx192(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx193(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx194(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx195(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx196(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx197(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx198(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx199(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx200(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx201(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx202(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx203(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx204(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx205(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx206(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx207(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx208(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx209(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx210(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx211(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx212(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx213(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx214(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx215(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx216(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx217(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx218(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx219(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx220(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx221(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx222(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx223(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx224(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx225(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx226(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx227(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx228(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx229(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx230(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx231(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx232(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx233(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx234(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx235(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx236(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx237(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx238(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx239(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx240(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx241(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx242(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx243(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx244(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx245(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx246(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx247(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx248(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx249(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx250(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx251(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx252(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx253(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx254(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx255(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx256(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx257(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx258(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx259(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx260(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx261(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx262(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx263(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx264(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx265(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx266(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx267(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx268(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx269(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx270(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx271(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx272(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx273(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx274(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx275(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx276(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx277(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx278(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx279(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx280(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx281(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx282(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx283(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx284(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx285(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx286(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx287(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx288(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx289(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx290(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx291(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx292(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx293(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx294(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx295(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx296(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx297(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx298(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx299(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx300(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx301(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx302(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx303(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx304(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx305(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx306(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx307(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx308(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx309(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx310(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx311(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx312(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx313(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx314(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx315(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx316(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx317(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx318(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx319(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx320(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx321(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx322(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx323(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx324(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx325(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx326(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx327(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx328(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx329(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx330(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx331(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx332(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx333(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx334(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx335(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx336(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx337(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx338(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx339(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx340(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx341(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx342(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx343(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx344(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx345(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx346(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx347(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx348(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx349(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx350(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx351(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx352(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx353(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx354(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx355(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx356(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx357(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx358(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx359(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx360(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx361(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx362(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx363(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx364(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx365(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx366(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx367(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx368(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx369(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx370(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx371(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx372(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx373(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx374(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx375(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx376(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx377(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx378(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx379(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx380(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx381(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx382(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx383(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx384(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx385(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx386(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx387(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx388(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx389(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx390(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx391(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx392(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx393(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx394(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx395(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx396(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx397(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx398(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx399(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx400(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx401(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx402(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx403(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx404(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx405(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx406(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx407(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx408(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx409(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx410(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx411(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx412(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx413(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx414(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx415(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx416(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx417(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx418(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx419(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx420(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx421(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx422(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx423(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx424(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx425(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx426(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx427(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx428(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx429(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx430(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx431(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx432(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx433(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx434(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx435(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx436(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx437(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx438(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx439(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx440(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx441(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx442(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx443(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx444(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx445(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx446(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx447(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx448(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx449(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx450(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx451(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx452(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx453(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx454(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx455(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx456(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx457(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx458(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx459(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx460(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx461(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx462(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx463(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx464(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx465(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx466(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx467(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx468(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx469(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx470(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx471(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx472(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx473(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx474(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx475(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx476(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx477(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx478(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx479(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx480(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx481(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx482(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx483(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx484(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx485(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx486(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx487(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx488(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx489(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx490(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx491(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx492(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx493(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx494(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx495(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx496(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx497(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx498(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx499(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx500(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx501(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx502(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx503(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx504(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx505(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx506(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx507(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx508(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx509(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx510(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx511(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx512(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx513(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx514(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx515(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx516(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx517(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx518(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx519(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx520(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx521(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx522(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx523(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx524(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx525(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx526(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx527(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx528(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx529(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx530(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx531(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx532(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx533(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx534(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx535(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx536(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx537(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx538(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx539(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module FX(x, y);
 input [674:0] x;
 output [539:0] y;

  Fx0 Fx0_inst(.x({x[1], x[0]}), .y(y[0]));
  Fx1 Fx1_inst(.x({x[2], x[0]}), .y(y[1]));
  Fx2 Fx2_inst(.x({x[3], x[0]}), .y(y[2]));
  Fx3 Fx3_inst(.x({x[4], x[0]}), .y(y[3]));
  Fx4 Fx4_inst(.x({x[6], x[5]}), .y(y[4]));
  Fx5 Fx5_inst(.x({x[7], x[5]}), .y(y[5]));
  Fx6 Fx6_inst(.x({x[8], x[5]}), .y(y[6]));
  Fx7 Fx7_inst(.x({x[9], x[5]}), .y(y[7]));
  Fx8 Fx8_inst(.x({x[11], x[10]}), .y(y[8]));
  Fx9 Fx9_inst(.x({x[12], x[10]}), .y(y[9]));
  Fx10 Fx10_inst(.x({x[13], x[10]}), .y(y[10]));
  Fx11 Fx11_inst(.x({x[14], x[10]}), .y(y[11]));
  Fx12 Fx12_inst(.x({x[16], x[15]}), .y(y[12]));
  Fx13 Fx13_inst(.x({x[17], x[15]}), .y(y[13]));
  Fx14 Fx14_inst(.x({x[18], x[15]}), .y(y[14]));
  Fx15 Fx15_inst(.x({x[19], x[15]}), .y(y[15]));
  Fx16 Fx16_inst(.x({x[21], x[20]}), .y(y[16]));
  Fx17 Fx17_inst(.x({x[22], x[20]}), .y(y[17]));
  Fx18 Fx18_inst(.x({x[23], x[20]}), .y(y[18]));
  Fx19 Fx19_inst(.x({x[24], x[20]}), .y(y[19]));
  Fx20 Fx20_inst(.x({x[26], x[25]}), .y(y[20]));
  Fx21 Fx21_inst(.x({x[27], x[25]}), .y(y[21]));
  Fx22 Fx22_inst(.x({x[28], x[25]}), .y(y[22]));
  Fx23 Fx23_inst(.x({x[29], x[25]}), .y(y[23]));
  Fx24 Fx24_inst(.x({x[31], x[30]}), .y(y[24]));
  Fx25 Fx25_inst(.x({x[32], x[30]}), .y(y[25]));
  Fx26 Fx26_inst(.x({x[33], x[30]}), .y(y[26]));
  Fx27 Fx27_inst(.x({x[34], x[30]}), .y(y[27]));
  Fx28 Fx28_inst(.x({x[36], x[35]}), .y(y[28]));
  Fx29 Fx29_inst(.x({x[37], x[35]}), .y(y[29]));
  Fx30 Fx30_inst(.x({x[38], x[35]}), .y(y[30]));
  Fx31 Fx31_inst(.x({x[39], x[35]}), .y(y[31]));
  Fx32 Fx32_inst(.x({x[41], x[40]}), .y(y[32]));
  Fx33 Fx33_inst(.x({x[42], x[40]}), .y(y[33]));
  Fx34 Fx34_inst(.x({x[43], x[40]}), .y(y[34]));
  Fx35 Fx35_inst(.x({x[44], x[40]}), .y(y[35]));
  Fx36 Fx36_inst(.x({x[46], x[45]}), .y(y[36]));
  Fx37 Fx37_inst(.x({x[47], x[45]}), .y(y[37]));
  Fx38 Fx38_inst(.x({x[48], x[45]}), .y(y[38]));
  Fx39 Fx39_inst(.x({x[49], x[45]}), .y(y[39]));
  Fx40 Fx40_inst(.x({x[51], x[50]}), .y(y[40]));
  Fx41 Fx41_inst(.x({x[52], x[50]}), .y(y[41]));
  Fx42 Fx42_inst(.x({x[53], x[50]}), .y(y[42]));
  Fx43 Fx43_inst(.x({x[54], x[50]}), .y(y[43]));
  Fx44 Fx44_inst(.x({x[56], x[55]}), .y(y[44]));
  Fx45 Fx45_inst(.x({x[57], x[55]}), .y(y[45]));
  Fx46 Fx46_inst(.x({x[58], x[55]}), .y(y[46]));
  Fx47 Fx47_inst(.x({x[59], x[55]}), .y(y[47]));
  Fx48 Fx48_inst(.x({x[61], x[60]}), .y(y[48]));
  Fx49 Fx49_inst(.x({x[62], x[60]}), .y(y[49]));
  Fx50 Fx50_inst(.x({x[63], x[60]}), .y(y[50]));
  Fx51 Fx51_inst(.x({x[64], x[60]}), .y(y[51]));
  Fx52 Fx52_inst(.x({x[66], x[65]}), .y(y[52]));
  Fx53 Fx53_inst(.x({x[67], x[65]}), .y(y[53]));
  Fx54 Fx54_inst(.x({x[68], x[65]}), .y(y[54]));
  Fx55 Fx55_inst(.x({x[69], x[65]}), .y(y[55]));
  Fx56 Fx56_inst(.x({x[71], x[70]}), .y(y[56]));
  Fx57 Fx57_inst(.x({x[72], x[70]}), .y(y[57]));
  Fx58 Fx58_inst(.x({x[73], x[70]}), .y(y[58]));
  Fx59 Fx59_inst(.x({x[74], x[70]}), .y(y[59]));
  Fx60 Fx60_inst(.x({x[76], x[75]}), .y(y[60]));
  Fx61 Fx61_inst(.x({x[77], x[75]}), .y(y[61]));
  Fx62 Fx62_inst(.x({x[78], x[75]}), .y(y[62]));
  Fx63 Fx63_inst(.x({x[79], x[75]}), .y(y[63]));
  Fx64 Fx64_inst(.x({x[81], x[80]}), .y(y[64]));
  Fx65 Fx65_inst(.x({x[82], x[80]}), .y(y[65]));
  Fx66 Fx66_inst(.x({x[83], x[80]}), .y(y[66]));
  Fx67 Fx67_inst(.x({x[84], x[80]}), .y(y[67]));
  Fx68 Fx68_inst(.x({x[86], x[85]}), .y(y[68]));
  Fx69 Fx69_inst(.x({x[87], x[85]}), .y(y[69]));
  Fx70 Fx70_inst(.x({x[88], x[85]}), .y(y[70]));
  Fx71 Fx71_inst(.x({x[89], x[85]}), .y(y[71]));
  Fx72 Fx72_inst(.x({x[91], x[90]}), .y(y[72]));
  Fx73 Fx73_inst(.x({x[92], x[90]}), .y(y[73]));
  Fx74 Fx74_inst(.x({x[93], x[90]}), .y(y[74]));
  Fx75 Fx75_inst(.x({x[94], x[90]}), .y(y[75]));
  Fx76 Fx76_inst(.x({x[96], x[95]}), .y(y[76]));
  Fx77 Fx77_inst(.x({x[97], x[95]}), .y(y[77]));
  Fx78 Fx78_inst(.x({x[98], x[95]}), .y(y[78]));
  Fx79 Fx79_inst(.x({x[99], x[95]}), .y(y[79]));
  Fx80 Fx80_inst(.x({x[101], x[100]}), .y(y[80]));
  Fx81 Fx81_inst(.x({x[102], x[100]}), .y(y[81]));
  Fx82 Fx82_inst(.x({x[103], x[100]}), .y(y[82]));
  Fx83 Fx83_inst(.x({x[104], x[100]}), .y(y[83]));
  Fx84 Fx84_inst(.x({x[106], x[105]}), .y(y[84]));
  Fx85 Fx85_inst(.x({x[107], x[105]}), .y(y[85]));
  Fx86 Fx86_inst(.x({x[108], x[105]}), .y(y[86]));
  Fx87 Fx87_inst(.x({x[109], x[105]}), .y(y[87]));
  Fx88 Fx88_inst(.x({x[111], x[110]}), .y(y[88]));
  Fx89 Fx89_inst(.x({x[112], x[110]}), .y(y[89]));
  Fx90 Fx90_inst(.x({x[113], x[110]}), .y(y[90]));
  Fx91 Fx91_inst(.x({x[114], x[110]}), .y(y[91]));
  Fx92 Fx92_inst(.x({x[116], x[115]}), .y(y[92]));
  Fx93 Fx93_inst(.x({x[117], x[115]}), .y(y[93]));
  Fx94 Fx94_inst(.x({x[118], x[115]}), .y(y[94]));
  Fx95 Fx95_inst(.x({x[119], x[115]}), .y(y[95]));
  Fx96 Fx96_inst(.x({x[121], x[120]}), .y(y[96]));
  Fx97 Fx97_inst(.x({x[122], x[120]}), .y(y[97]));
  Fx98 Fx98_inst(.x({x[123], x[120]}), .y(y[98]));
  Fx99 Fx99_inst(.x({x[124], x[120]}), .y(y[99]));
  Fx100 Fx100_inst(.x({x[126], x[125]}), .y(y[100]));
  Fx101 Fx101_inst(.x({x[127], x[125]}), .y(y[101]));
  Fx102 Fx102_inst(.x({x[128], x[125]}), .y(y[102]));
  Fx103 Fx103_inst(.x({x[129], x[125]}), .y(y[103]));
  Fx104 Fx104_inst(.x({x[131], x[130]}), .y(y[104]));
  Fx105 Fx105_inst(.x({x[132], x[130]}), .y(y[105]));
  Fx106 Fx106_inst(.x({x[133], x[130]}), .y(y[106]));
  Fx107 Fx107_inst(.x({x[134], x[130]}), .y(y[107]));
  Fx108 Fx108_inst(.x({x[136], x[135]}), .y(y[108]));
  Fx109 Fx109_inst(.x({x[137], x[135]}), .y(y[109]));
  Fx110 Fx110_inst(.x({x[138], x[135]}), .y(y[110]));
  Fx111 Fx111_inst(.x({x[139], x[135]}), .y(y[111]));
  Fx112 Fx112_inst(.x({x[141], x[140]}), .y(y[112]));
  Fx113 Fx113_inst(.x({x[142], x[140]}), .y(y[113]));
  Fx114 Fx114_inst(.x({x[143], x[140]}), .y(y[114]));
  Fx115 Fx115_inst(.x({x[144], x[140]}), .y(y[115]));
  Fx116 Fx116_inst(.x({x[146], x[145]}), .y(y[116]));
  Fx117 Fx117_inst(.x({x[147], x[145]}), .y(y[117]));
  Fx118 Fx118_inst(.x({x[148], x[145]}), .y(y[118]));
  Fx119 Fx119_inst(.x({x[149], x[145]}), .y(y[119]));
  Fx120 Fx120_inst(.x({x[151], x[150]}), .y(y[120]));
  Fx121 Fx121_inst(.x({x[152], x[150]}), .y(y[121]));
  Fx122 Fx122_inst(.x({x[153], x[150]}), .y(y[122]));
  Fx123 Fx123_inst(.x({x[154], x[150]}), .y(y[123]));
  Fx124 Fx124_inst(.x({x[156], x[155]}), .y(y[124]));
  Fx125 Fx125_inst(.x({x[157], x[155]}), .y(y[125]));
  Fx126 Fx126_inst(.x({x[158], x[155]}), .y(y[126]));
  Fx127 Fx127_inst(.x({x[159], x[155]}), .y(y[127]));
  Fx128 Fx128_inst(.x({x[161], x[160]}), .y(y[128]));
  Fx129 Fx129_inst(.x({x[162], x[160]}), .y(y[129]));
  Fx130 Fx130_inst(.x({x[163], x[160]}), .y(y[130]));
  Fx131 Fx131_inst(.x({x[164], x[160]}), .y(y[131]));
  Fx132 Fx132_inst(.x({x[166], x[165]}), .y(y[132]));
  Fx133 Fx133_inst(.x({x[167], x[165]}), .y(y[133]));
  Fx134 Fx134_inst(.x({x[168], x[165]}), .y(y[134]));
  Fx135 Fx135_inst(.x({x[169], x[165]}), .y(y[135]));
  Fx136 Fx136_inst(.x({x[171], x[170]}), .y(y[136]));
  Fx137 Fx137_inst(.x({x[172], x[170]}), .y(y[137]));
  Fx138 Fx138_inst(.x({x[173], x[170]}), .y(y[138]));
  Fx139 Fx139_inst(.x({x[174], x[170]}), .y(y[139]));
  Fx140 Fx140_inst(.x({x[176], x[175]}), .y(y[140]));
  Fx141 Fx141_inst(.x({x[177], x[175]}), .y(y[141]));
  Fx142 Fx142_inst(.x({x[178], x[175]}), .y(y[142]));
  Fx143 Fx143_inst(.x({x[179], x[175]}), .y(y[143]));
  Fx144 Fx144_inst(.x({x[181], x[180]}), .y(y[144]));
  Fx145 Fx145_inst(.x({x[182], x[180]}), .y(y[145]));
  Fx146 Fx146_inst(.x({x[183], x[180]}), .y(y[146]));
  Fx147 Fx147_inst(.x({x[184], x[180]}), .y(y[147]));
  Fx148 Fx148_inst(.x({x[186], x[185]}), .y(y[148]));
  Fx149 Fx149_inst(.x({x[187], x[185]}), .y(y[149]));
  Fx150 Fx150_inst(.x({x[188], x[185]}), .y(y[150]));
  Fx151 Fx151_inst(.x({x[189], x[185]}), .y(y[151]));
  Fx152 Fx152_inst(.x({x[191], x[190]}), .y(y[152]));
  Fx153 Fx153_inst(.x({x[192], x[190]}), .y(y[153]));
  Fx154 Fx154_inst(.x({x[193], x[190]}), .y(y[154]));
  Fx155 Fx155_inst(.x({x[194], x[190]}), .y(y[155]));
  Fx156 Fx156_inst(.x({x[196], x[195]}), .y(y[156]));
  Fx157 Fx157_inst(.x({x[197], x[195]}), .y(y[157]));
  Fx158 Fx158_inst(.x({x[198], x[195]}), .y(y[158]));
  Fx159 Fx159_inst(.x({x[199], x[195]}), .y(y[159]));
  Fx160 Fx160_inst(.x({x[201], x[200]}), .y(y[160]));
  Fx161 Fx161_inst(.x({x[202], x[200]}), .y(y[161]));
  Fx162 Fx162_inst(.x({x[203], x[200]}), .y(y[162]));
  Fx163 Fx163_inst(.x({x[204], x[200]}), .y(y[163]));
  Fx164 Fx164_inst(.x({x[206], x[205]}), .y(y[164]));
  Fx165 Fx165_inst(.x({x[207], x[205]}), .y(y[165]));
  Fx166 Fx166_inst(.x({x[208], x[205]}), .y(y[166]));
  Fx167 Fx167_inst(.x({x[209], x[205]}), .y(y[167]));
  Fx168 Fx168_inst(.x({x[211], x[210]}), .y(y[168]));
  Fx169 Fx169_inst(.x({x[212], x[210]}), .y(y[169]));
  Fx170 Fx170_inst(.x({x[213], x[210]}), .y(y[170]));
  Fx171 Fx171_inst(.x({x[214], x[210]}), .y(y[171]));
  Fx172 Fx172_inst(.x({x[216], x[215]}), .y(y[172]));
  Fx173 Fx173_inst(.x({x[217], x[215]}), .y(y[173]));
  Fx174 Fx174_inst(.x({x[218], x[215]}), .y(y[174]));
  Fx175 Fx175_inst(.x({x[219], x[215]}), .y(y[175]));
  Fx176 Fx176_inst(.x({x[221], x[220]}), .y(y[176]));
  Fx177 Fx177_inst(.x({x[222], x[220]}), .y(y[177]));
  Fx178 Fx178_inst(.x({x[223], x[220]}), .y(y[178]));
  Fx179 Fx179_inst(.x({x[224], x[220]}), .y(y[179]));
  Fx180 Fx180_inst(.x({x[226], x[225]}), .y(y[180]));
  Fx181 Fx181_inst(.x({x[227], x[225]}), .y(y[181]));
  Fx182 Fx182_inst(.x({x[228], x[225]}), .y(y[182]));
  Fx183 Fx183_inst(.x({x[229], x[225]}), .y(y[183]));
  Fx184 Fx184_inst(.x({x[231], x[230]}), .y(y[184]));
  Fx185 Fx185_inst(.x({x[232], x[230]}), .y(y[185]));
  Fx186 Fx186_inst(.x({x[233], x[230]}), .y(y[186]));
  Fx187 Fx187_inst(.x({x[234], x[230]}), .y(y[187]));
  Fx188 Fx188_inst(.x({x[236], x[235]}), .y(y[188]));
  Fx189 Fx189_inst(.x({x[237], x[235]}), .y(y[189]));
  Fx190 Fx190_inst(.x({x[238], x[235]}), .y(y[190]));
  Fx191 Fx191_inst(.x({x[239], x[235]}), .y(y[191]));
  Fx192 Fx192_inst(.x({x[241], x[240]}), .y(y[192]));
  Fx193 Fx193_inst(.x({x[242], x[240]}), .y(y[193]));
  Fx194 Fx194_inst(.x({x[243], x[240]}), .y(y[194]));
  Fx195 Fx195_inst(.x({x[244], x[240]}), .y(y[195]));
  Fx196 Fx196_inst(.x({x[246], x[245]}), .y(y[196]));
  Fx197 Fx197_inst(.x({x[247], x[245]}), .y(y[197]));
  Fx198 Fx198_inst(.x({x[248], x[245]}), .y(y[198]));
  Fx199 Fx199_inst(.x({x[249], x[245]}), .y(y[199]));
  Fx200 Fx200_inst(.x({x[251], x[250]}), .y(y[200]));
  Fx201 Fx201_inst(.x({x[252], x[250]}), .y(y[201]));
  Fx202 Fx202_inst(.x({x[253], x[250]}), .y(y[202]));
  Fx203 Fx203_inst(.x({x[254], x[250]}), .y(y[203]));
  Fx204 Fx204_inst(.x({x[256], x[255]}), .y(y[204]));
  Fx205 Fx205_inst(.x({x[257], x[255]}), .y(y[205]));
  Fx206 Fx206_inst(.x({x[258], x[255]}), .y(y[206]));
  Fx207 Fx207_inst(.x({x[259], x[255]}), .y(y[207]));
  Fx208 Fx208_inst(.x({x[261], x[260]}), .y(y[208]));
  Fx209 Fx209_inst(.x({x[262], x[260]}), .y(y[209]));
  Fx210 Fx210_inst(.x({x[263], x[260]}), .y(y[210]));
  Fx211 Fx211_inst(.x({x[264], x[260]}), .y(y[211]));
  Fx212 Fx212_inst(.x({x[266], x[265]}), .y(y[212]));
  Fx213 Fx213_inst(.x({x[267], x[265]}), .y(y[213]));
  Fx214 Fx214_inst(.x({x[268], x[265]}), .y(y[214]));
  Fx215 Fx215_inst(.x({x[269], x[265]}), .y(y[215]));
  Fx216 Fx216_inst(.x({x[271], x[270]}), .y(y[216]));
  Fx217 Fx217_inst(.x({x[272], x[270]}), .y(y[217]));
  Fx218 Fx218_inst(.x({x[273], x[270]}), .y(y[218]));
  Fx219 Fx219_inst(.x({x[274], x[270]}), .y(y[219]));
  Fx220 Fx220_inst(.x({x[276], x[275]}), .y(y[220]));
  Fx221 Fx221_inst(.x({x[277], x[275]}), .y(y[221]));
  Fx222 Fx222_inst(.x({x[278], x[275]}), .y(y[222]));
  Fx223 Fx223_inst(.x({x[279], x[275]}), .y(y[223]));
  Fx224 Fx224_inst(.x({x[281], x[280]}), .y(y[224]));
  Fx225 Fx225_inst(.x({x[282], x[280]}), .y(y[225]));
  Fx226 Fx226_inst(.x({x[283], x[280]}), .y(y[226]));
  Fx227 Fx227_inst(.x({x[284], x[280]}), .y(y[227]));
  Fx228 Fx228_inst(.x({x[286], x[285]}), .y(y[228]));
  Fx229 Fx229_inst(.x({x[287], x[285]}), .y(y[229]));
  Fx230 Fx230_inst(.x({x[288], x[285]}), .y(y[230]));
  Fx231 Fx231_inst(.x({x[289], x[285]}), .y(y[231]));
  Fx232 Fx232_inst(.x({x[291], x[290]}), .y(y[232]));
  Fx233 Fx233_inst(.x({x[292], x[290]}), .y(y[233]));
  Fx234 Fx234_inst(.x({x[293], x[290]}), .y(y[234]));
  Fx235 Fx235_inst(.x({x[294], x[290]}), .y(y[235]));
  Fx236 Fx236_inst(.x({x[296], x[295]}), .y(y[236]));
  Fx237 Fx237_inst(.x({x[297], x[295]}), .y(y[237]));
  Fx238 Fx238_inst(.x({x[298], x[295]}), .y(y[238]));
  Fx239 Fx239_inst(.x({x[299], x[295]}), .y(y[239]));
  Fx240 Fx240_inst(.x({x[301], x[300]}), .y(y[240]));
  Fx241 Fx241_inst(.x({x[302], x[300]}), .y(y[241]));
  Fx242 Fx242_inst(.x({x[303], x[300]}), .y(y[242]));
  Fx243 Fx243_inst(.x({x[304], x[300]}), .y(y[243]));
  Fx244 Fx244_inst(.x({x[306], x[305]}), .y(y[244]));
  Fx245 Fx245_inst(.x({x[307], x[305]}), .y(y[245]));
  Fx246 Fx246_inst(.x({x[308], x[305]}), .y(y[246]));
  Fx247 Fx247_inst(.x({x[309], x[305]}), .y(y[247]));
  Fx248 Fx248_inst(.x({x[311], x[310]}), .y(y[248]));
  Fx249 Fx249_inst(.x({x[312], x[310]}), .y(y[249]));
  Fx250 Fx250_inst(.x({x[313], x[310]}), .y(y[250]));
  Fx251 Fx251_inst(.x({x[314], x[310]}), .y(y[251]));
  Fx252 Fx252_inst(.x({x[316], x[315]}), .y(y[252]));
  Fx253 Fx253_inst(.x({x[317], x[315]}), .y(y[253]));
  Fx254 Fx254_inst(.x({x[318], x[315]}), .y(y[254]));
  Fx255 Fx255_inst(.x({x[319], x[315]}), .y(y[255]));
  Fx256 Fx256_inst(.x({x[321], x[320]}), .y(y[256]));
  Fx257 Fx257_inst(.x({x[322], x[320]}), .y(y[257]));
  Fx258 Fx258_inst(.x({x[323], x[320]}), .y(y[258]));
  Fx259 Fx259_inst(.x({x[324], x[320]}), .y(y[259]));
  Fx260 Fx260_inst(.x({x[326], x[325]}), .y(y[260]));
  Fx261 Fx261_inst(.x({x[327], x[325]}), .y(y[261]));
  Fx262 Fx262_inst(.x({x[328], x[325]}), .y(y[262]));
  Fx263 Fx263_inst(.x({x[329], x[325]}), .y(y[263]));
  Fx264 Fx264_inst(.x({x[331], x[330]}), .y(y[264]));
  Fx265 Fx265_inst(.x({x[332], x[330]}), .y(y[265]));
  Fx266 Fx266_inst(.x({x[333], x[330]}), .y(y[266]));
  Fx267 Fx267_inst(.x({x[334], x[330]}), .y(y[267]));
  Fx268 Fx268_inst(.x({x[336], x[335]}), .y(y[268]));
  Fx269 Fx269_inst(.x({x[337], x[335]}), .y(y[269]));
  Fx270 Fx270_inst(.x({x[338], x[335]}), .y(y[270]));
  Fx271 Fx271_inst(.x({x[339], x[335]}), .y(y[271]));
  Fx272 Fx272_inst(.x({x[341], x[340]}), .y(y[272]));
  Fx273 Fx273_inst(.x({x[342], x[340]}), .y(y[273]));
  Fx274 Fx274_inst(.x({x[343], x[340]}), .y(y[274]));
  Fx275 Fx275_inst(.x({x[344], x[340]}), .y(y[275]));
  Fx276 Fx276_inst(.x({x[346], x[345]}), .y(y[276]));
  Fx277 Fx277_inst(.x({x[347], x[345]}), .y(y[277]));
  Fx278 Fx278_inst(.x({x[348], x[345]}), .y(y[278]));
  Fx279 Fx279_inst(.x({x[349], x[345]}), .y(y[279]));
  Fx280 Fx280_inst(.x({x[351], x[350]}), .y(y[280]));
  Fx281 Fx281_inst(.x({x[352], x[350]}), .y(y[281]));
  Fx282 Fx282_inst(.x({x[353], x[350]}), .y(y[282]));
  Fx283 Fx283_inst(.x({x[354], x[350]}), .y(y[283]));
  Fx284 Fx284_inst(.x({x[356], x[355]}), .y(y[284]));
  Fx285 Fx285_inst(.x({x[357], x[355]}), .y(y[285]));
  Fx286 Fx286_inst(.x({x[358], x[355]}), .y(y[286]));
  Fx287 Fx287_inst(.x({x[359], x[355]}), .y(y[287]));
  Fx288 Fx288_inst(.x({x[361], x[360]}), .y(y[288]));
  Fx289 Fx289_inst(.x({x[362], x[360]}), .y(y[289]));
  Fx290 Fx290_inst(.x({x[363], x[360]}), .y(y[290]));
  Fx291 Fx291_inst(.x({x[364], x[360]}), .y(y[291]));
  Fx292 Fx292_inst(.x({x[366], x[365]}), .y(y[292]));
  Fx293 Fx293_inst(.x({x[367], x[365]}), .y(y[293]));
  Fx294 Fx294_inst(.x({x[368], x[365]}), .y(y[294]));
  Fx295 Fx295_inst(.x({x[369], x[365]}), .y(y[295]));
  Fx296 Fx296_inst(.x({x[371], x[370]}), .y(y[296]));
  Fx297 Fx297_inst(.x({x[372], x[370]}), .y(y[297]));
  Fx298 Fx298_inst(.x({x[373], x[370]}), .y(y[298]));
  Fx299 Fx299_inst(.x({x[374], x[370]}), .y(y[299]));
  Fx300 Fx300_inst(.x({x[376], x[375]}), .y(y[300]));
  Fx301 Fx301_inst(.x({x[377], x[375]}), .y(y[301]));
  Fx302 Fx302_inst(.x({x[378], x[375]}), .y(y[302]));
  Fx303 Fx303_inst(.x({x[379], x[375]}), .y(y[303]));
  Fx304 Fx304_inst(.x({x[381], x[380]}), .y(y[304]));
  Fx305 Fx305_inst(.x({x[382], x[380]}), .y(y[305]));
  Fx306 Fx306_inst(.x({x[383], x[380]}), .y(y[306]));
  Fx307 Fx307_inst(.x({x[384], x[380]}), .y(y[307]));
  Fx308 Fx308_inst(.x({x[386], x[385]}), .y(y[308]));
  Fx309 Fx309_inst(.x({x[387], x[385]}), .y(y[309]));
  Fx310 Fx310_inst(.x({x[388], x[385]}), .y(y[310]));
  Fx311 Fx311_inst(.x({x[389], x[385]}), .y(y[311]));
  Fx312 Fx312_inst(.x({x[391], x[390]}), .y(y[312]));
  Fx313 Fx313_inst(.x({x[392], x[390]}), .y(y[313]));
  Fx314 Fx314_inst(.x({x[393], x[390]}), .y(y[314]));
  Fx315 Fx315_inst(.x({x[394], x[390]}), .y(y[315]));
  Fx316 Fx316_inst(.x({x[396], x[395]}), .y(y[316]));
  Fx317 Fx317_inst(.x({x[397], x[395]}), .y(y[317]));
  Fx318 Fx318_inst(.x({x[398], x[395]}), .y(y[318]));
  Fx319 Fx319_inst(.x({x[399], x[395]}), .y(y[319]));
  Fx320 Fx320_inst(.x({x[401], x[400]}), .y(y[320]));
  Fx321 Fx321_inst(.x({x[402], x[400]}), .y(y[321]));
  Fx322 Fx322_inst(.x({x[403], x[400]}), .y(y[322]));
  Fx323 Fx323_inst(.x({x[404], x[400]}), .y(y[323]));
  Fx324 Fx324_inst(.x({x[406], x[405]}), .y(y[324]));
  Fx325 Fx325_inst(.x({x[407], x[405]}), .y(y[325]));
  Fx326 Fx326_inst(.x({x[408], x[405]}), .y(y[326]));
  Fx327 Fx327_inst(.x({x[409], x[405]}), .y(y[327]));
  Fx328 Fx328_inst(.x({x[411], x[410]}), .y(y[328]));
  Fx329 Fx329_inst(.x({x[412], x[410]}), .y(y[329]));
  Fx330 Fx330_inst(.x({x[413], x[410]}), .y(y[330]));
  Fx331 Fx331_inst(.x({x[414], x[410]}), .y(y[331]));
  Fx332 Fx332_inst(.x({x[416], x[415]}), .y(y[332]));
  Fx333 Fx333_inst(.x({x[417], x[415]}), .y(y[333]));
  Fx334 Fx334_inst(.x({x[418], x[415]}), .y(y[334]));
  Fx335 Fx335_inst(.x({x[419], x[415]}), .y(y[335]));
  Fx336 Fx336_inst(.x({x[421], x[420]}), .y(y[336]));
  Fx337 Fx337_inst(.x({x[422], x[420]}), .y(y[337]));
  Fx338 Fx338_inst(.x({x[423], x[420]}), .y(y[338]));
  Fx339 Fx339_inst(.x({x[424], x[420]}), .y(y[339]));
  Fx340 Fx340_inst(.x({x[426], x[425]}), .y(y[340]));
  Fx341 Fx341_inst(.x({x[427], x[425]}), .y(y[341]));
  Fx342 Fx342_inst(.x({x[428], x[425]}), .y(y[342]));
  Fx343 Fx343_inst(.x({x[429], x[425]}), .y(y[343]));
  Fx344 Fx344_inst(.x({x[431], x[430]}), .y(y[344]));
  Fx345 Fx345_inst(.x({x[432], x[430]}), .y(y[345]));
  Fx346 Fx346_inst(.x({x[433], x[430]}), .y(y[346]));
  Fx347 Fx347_inst(.x({x[434], x[430]}), .y(y[347]));
  Fx348 Fx348_inst(.x({x[436], x[435]}), .y(y[348]));
  Fx349 Fx349_inst(.x({x[437], x[435]}), .y(y[349]));
  Fx350 Fx350_inst(.x({x[438], x[435]}), .y(y[350]));
  Fx351 Fx351_inst(.x({x[439], x[435]}), .y(y[351]));
  Fx352 Fx352_inst(.x({x[441], x[440]}), .y(y[352]));
  Fx353 Fx353_inst(.x({x[442], x[440]}), .y(y[353]));
  Fx354 Fx354_inst(.x({x[443], x[440]}), .y(y[354]));
  Fx355 Fx355_inst(.x({x[444], x[440]}), .y(y[355]));
  Fx356 Fx356_inst(.x({x[446], x[445]}), .y(y[356]));
  Fx357 Fx357_inst(.x({x[447], x[445]}), .y(y[357]));
  Fx358 Fx358_inst(.x({x[448], x[445]}), .y(y[358]));
  Fx359 Fx359_inst(.x({x[449], x[445]}), .y(y[359]));
  Fx360 Fx360_inst(.x({x[451], x[450]}), .y(y[360]));
  Fx361 Fx361_inst(.x({x[452], x[450]}), .y(y[361]));
  Fx362 Fx362_inst(.x({x[453], x[450]}), .y(y[362]));
  Fx363 Fx363_inst(.x({x[454], x[450]}), .y(y[363]));
  Fx364 Fx364_inst(.x({x[456], x[455]}), .y(y[364]));
  Fx365 Fx365_inst(.x({x[457], x[455]}), .y(y[365]));
  Fx366 Fx366_inst(.x({x[458], x[455]}), .y(y[366]));
  Fx367 Fx367_inst(.x({x[459], x[455]}), .y(y[367]));
  Fx368 Fx368_inst(.x({x[461], x[460]}), .y(y[368]));
  Fx369 Fx369_inst(.x({x[462], x[460]}), .y(y[369]));
  Fx370 Fx370_inst(.x({x[463], x[460]}), .y(y[370]));
  Fx371 Fx371_inst(.x({x[464], x[460]}), .y(y[371]));
  Fx372 Fx372_inst(.x({x[466], x[465]}), .y(y[372]));
  Fx373 Fx373_inst(.x({x[467], x[465]}), .y(y[373]));
  Fx374 Fx374_inst(.x({x[468], x[465]}), .y(y[374]));
  Fx375 Fx375_inst(.x({x[469], x[465]}), .y(y[375]));
  Fx376 Fx376_inst(.x({x[471], x[470]}), .y(y[376]));
  Fx377 Fx377_inst(.x({x[472], x[470]}), .y(y[377]));
  Fx378 Fx378_inst(.x({x[473], x[470]}), .y(y[378]));
  Fx379 Fx379_inst(.x({x[474], x[470]}), .y(y[379]));
  Fx380 Fx380_inst(.x({x[476], x[475]}), .y(y[380]));
  Fx381 Fx381_inst(.x({x[477], x[475]}), .y(y[381]));
  Fx382 Fx382_inst(.x({x[478], x[475]}), .y(y[382]));
  Fx383 Fx383_inst(.x({x[479], x[475]}), .y(y[383]));
  Fx384 Fx384_inst(.x({x[481], x[480]}), .y(y[384]));
  Fx385 Fx385_inst(.x({x[482], x[480]}), .y(y[385]));
  Fx386 Fx386_inst(.x({x[483], x[480]}), .y(y[386]));
  Fx387 Fx387_inst(.x({x[484], x[480]}), .y(y[387]));
  Fx388 Fx388_inst(.x({x[486], x[485]}), .y(y[388]));
  Fx389 Fx389_inst(.x({x[487], x[485]}), .y(y[389]));
  Fx390 Fx390_inst(.x({x[488], x[485]}), .y(y[390]));
  Fx391 Fx391_inst(.x({x[489], x[485]}), .y(y[391]));
  Fx392 Fx392_inst(.x({x[491], x[490]}), .y(y[392]));
  Fx393 Fx393_inst(.x({x[492], x[490]}), .y(y[393]));
  Fx394 Fx394_inst(.x({x[493], x[490]}), .y(y[394]));
  Fx395 Fx395_inst(.x({x[494], x[490]}), .y(y[395]));
  Fx396 Fx396_inst(.x({x[496], x[495]}), .y(y[396]));
  Fx397 Fx397_inst(.x({x[497], x[495]}), .y(y[397]));
  Fx398 Fx398_inst(.x({x[498], x[495]}), .y(y[398]));
  Fx399 Fx399_inst(.x({x[499], x[495]}), .y(y[399]));
  Fx400 Fx400_inst(.x({x[501], x[500]}), .y(y[400]));
  Fx401 Fx401_inst(.x({x[502], x[500]}), .y(y[401]));
  Fx402 Fx402_inst(.x({x[503], x[500]}), .y(y[402]));
  Fx403 Fx403_inst(.x({x[504], x[500]}), .y(y[403]));
  Fx404 Fx404_inst(.x({x[506], x[505]}), .y(y[404]));
  Fx405 Fx405_inst(.x({x[507], x[505]}), .y(y[405]));
  Fx406 Fx406_inst(.x({x[508], x[505]}), .y(y[406]));
  Fx407 Fx407_inst(.x({x[509], x[505]}), .y(y[407]));
  Fx408 Fx408_inst(.x({x[511], x[510]}), .y(y[408]));
  Fx409 Fx409_inst(.x({x[512], x[510]}), .y(y[409]));
  Fx410 Fx410_inst(.x({x[513], x[510]}), .y(y[410]));
  Fx411 Fx411_inst(.x({x[514], x[510]}), .y(y[411]));
  Fx412 Fx412_inst(.x({x[516], x[515]}), .y(y[412]));
  Fx413 Fx413_inst(.x({x[517], x[515]}), .y(y[413]));
  Fx414 Fx414_inst(.x({x[518], x[515]}), .y(y[414]));
  Fx415 Fx415_inst(.x({x[519], x[515]}), .y(y[415]));
  Fx416 Fx416_inst(.x({x[521], x[520]}), .y(y[416]));
  Fx417 Fx417_inst(.x({x[522], x[520]}), .y(y[417]));
  Fx418 Fx418_inst(.x({x[523], x[520]}), .y(y[418]));
  Fx419 Fx419_inst(.x({x[524], x[520]}), .y(y[419]));
  Fx420 Fx420_inst(.x({x[526], x[525]}), .y(y[420]));
  Fx421 Fx421_inst(.x({x[527], x[525]}), .y(y[421]));
  Fx422 Fx422_inst(.x({x[528], x[525]}), .y(y[422]));
  Fx423 Fx423_inst(.x({x[529], x[525]}), .y(y[423]));
  Fx424 Fx424_inst(.x({x[531], x[530]}), .y(y[424]));
  Fx425 Fx425_inst(.x({x[532], x[530]}), .y(y[425]));
  Fx426 Fx426_inst(.x({x[533], x[530]}), .y(y[426]));
  Fx427 Fx427_inst(.x({x[534], x[530]}), .y(y[427]));
  Fx428 Fx428_inst(.x({x[536], x[535]}), .y(y[428]));
  Fx429 Fx429_inst(.x({x[537], x[535]}), .y(y[429]));
  Fx430 Fx430_inst(.x({x[538], x[535]}), .y(y[430]));
  Fx431 Fx431_inst(.x({x[539], x[535]}), .y(y[431]));
  Fx432 Fx432_inst(.x({x[541], x[540]}), .y(y[432]));
  Fx433 Fx433_inst(.x({x[542], x[540]}), .y(y[433]));
  Fx434 Fx434_inst(.x({x[543], x[540]}), .y(y[434]));
  Fx435 Fx435_inst(.x({x[544], x[540]}), .y(y[435]));
  Fx436 Fx436_inst(.x({x[546], x[545]}), .y(y[436]));
  Fx437 Fx437_inst(.x({x[547], x[545]}), .y(y[437]));
  Fx438 Fx438_inst(.x({x[548], x[545]}), .y(y[438]));
  Fx439 Fx439_inst(.x({x[549], x[545]}), .y(y[439]));
  Fx440 Fx440_inst(.x({x[551], x[550]}), .y(y[440]));
  Fx441 Fx441_inst(.x({x[552], x[550]}), .y(y[441]));
  Fx442 Fx442_inst(.x({x[553], x[550]}), .y(y[442]));
  Fx443 Fx443_inst(.x({x[554], x[550]}), .y(y[443]));
  Fx444 Fx444_inst(.x({x[556], x[555]}), .y(y[444]));
  Fx445 Fx445_inst(.x({x[557], x[555]}), .y(y[445]));
  Fx446 Fx446_inst(.x({x[558], x[555]}), .y(y[446]));
  Fx447 Fx447_inst(.x({x[559], x[555]}), .y(y[447]));
  Fx448 Fx448_inst(.x({x[561], x[560]}), .y(y[448]));
  Fx449 Fx449_inst(.x({x[562], x[560]}), .y(y[449]));
  Fx450 Fx450_inst(.x({x[563], x[560]}), .y(y[450]));
  Fx451 Fx451_inst(.x({x[564], x[560]}), .y(y[451]));
  Fx452 Fx452_inst(.x({x[566], x[565]}), .y(y[452]));
  Fx453 Fx453_inst(.x({x[567], x[565]}), .y(y[453]));
  Fx454 Fx454_inst(.x({x[568], x[565]}), .y(y[454]));
  Fx455 Fx455_inst(.x({x[569], x[565]}), .y(y[455]));
  Fx456 Fx456_inst(.x({x[571], x[570]}), .y(y[456]));
  Fx457 Fx457_inst(.x({x[572], x[570]}), .y(y[457]));
  Fx458 Fx458_inst(.x({x[573], x[570]}), .y(y[458]));
  Fx459 Fx459_inst(.x({x[574], x[570]}), .y(y[459]));
  Fx460 Fx460_inst(.x({x[576], x[575]}), .y(y[460]));
  Fx461 Fx461_inst(.x({x[577], x[575]}), .y(y[461]));
  Fx462 Fx462_inst(.x({x[578], x[575]}), .y(y[462]));
  Fx463 Fx463_inst(.x({x[579], x[575]}), .y(y[463]));
  Fx464 Fx464_inst(.x({x[581], x[580]}), .y(y[464]));
  Fx465 Fx465_inst(.x({x[582], x[580]}), .y(y[465]));
  Fx466 Fx466_inst(.x({x[583], x[580]}), .y(y[466]));
  Fx467 Fx467_inst(.x({x[584], x[580]}), .y(y[467]));
  Fx468 Fx468_inst(.x({x[586], x[585]}), .y(y[468]));
  Fx469 Fx469_inst(.x({x[587], x[585]}), .y(y[469]));
  Fx470 Fx470_inst(.x({x[588], x[585]}), .y(y[470]));
  Fx471 Fx471_inst(.x({x[589], x[585]}), .y(y[471]));
  Fx472 Fx472_inst(.x({x[591], x[590]}), .y(y[472]));
  Fx473 Fx473_inst(.x({x[592], x[590]}), .y(y[473]));
  Fx474 Fx474_inst(.x({x[593], x[590]}), .y(y[474]));
  Fx475 Fx475_inst(.x({x[594], x[590]}), .y(y[475]));
  Fx476 Fx476_inst(.x({x[596], x[595]}), .y(y[476]));
  Fx477 Fx477_inst(.x({x[597], x[595]}), .y(y[477]));
  Fx478 Fx478_inst(.x({x[598], x[595]}), .y(y[478]));
  Fx479 Fx479_inst(.x({x[599], x[595]}), .y(y[479]));
  Fx480 Fx480_inst(.x({x[601], x[600]}), .y(y[480]));
  Fx481 Fx481_inst(.x({x[602], x[600]}), .y(y[481]));
  Fx482 Fx482_inst(.x({x[603], x[600]}), .y(y[482]));
  Fx483 Fx483_inst(.x({x[604], x[600]}), .y(y[483]));
  Fx484 Fx484_inst(.x({x[606], x[605]}), .y(y[484]));
  Fx485 Fx485_inst(.x({x[607], x[605]}), .y(y[485]));
  Fx486 Fx486_inst(.x({x[608], x[605]}), .y(y[486]));
  Fx487 Fx487_inst(.x({x[609], x[605]}), .y(y[487]));
  Fx488 Fx488_inst(.x({x[611], x[610]}), .y(y[488]));
  Fx489 Fx489_inst(.x({x[612], x[610]}), .y(y[489]));
  Fx490 Fx490_inst(.x({x[613], x[610]}), .y(y[490]));
  Fx491 Fx491_inst(.x({x[614], x[610]}), .y(y[491]));
  Fx492 Fx492_inst(.x({x[616], x[615]}), .y(y[492]));
  Fx493 Fx493_inst(.x({x[617], x[615]}), .y(y[493]));
  Fx494 Fx494_inst(.x({x[618], x[615]}), .y(y[494]));
  Fx495 Fx495_inst(.x({x[619], x[615]}), .y(y[495]));
  Fx496 Fx496_inst(.x({x[621], x[620]}), .y(y[496]));
  Fx497 Fx497_inst(.x({x[622], x[620]}), .y(y[497]));
  Fx498 Fx498_inst(.x({x[623], x[620]}), .y(y[498]));
  Fx499 Fx499_inst(.x({x[624], x[620]}), .y(y[499]));
  Fx500 Fx500_inst(.x({x[626], x[625]}), .y(y[500]));
  Fx501 Fx501_inst(.x({x[627], x[625]}), .y(y[501]));
  Fx502 Fx502_inst(.x({x[628], x[625]}), .y(y[502]));
  Fx503 Fx503_inst(.x({x[629], x[625]}), .y(y[503]));
  Fx504 Fx504_inst(.x({x[631], x[630]}), .y(y[504]));
  Fx505 Fx505_inst(.x({x[632], x[630]}), .y(y[505]));
  Fx506 Fx506_inst(.x({x[633], x[630]}), .y(y[506]));
  Fx507 Fx507_inst(.x({x[634], x[630]}), .y(y[507]));
  Fx508 Fx508_inst(.x({x[636], x[635]}), .y(y[508]));
  Fx509 Fx509_inst(.x({x[637], x[635]}), .y(y[509]));
  Fx510 Fx510_inst(.x({x[638], x[635]}), .y(y[510]));
  Fx511 Fx511_inst(.x({x[639], x[635]}), .y(y[511]));
  Fx512 Fx512_inst(.x({x[641], x[640]}), .y(y[512]));
  Fx513 Fx513_inst(.x({x[642], x[640]}), .y(y[513]));
  Fx514 Fx514_inst(.x({x[643], x[640]}), .y(y[514]));
  Fx515 Fx515_inst(.x({x[644], x[640]}), .y(y[515]));
  Fx516 Fx516_inst(.x({x[646], x[645]}), .y(y[516]));
  Fx517 Fx517_inst(.x({x[647], x[645]}), .y(y[517]));
  Fx518 Fx518_inst(.x({x[648], x[645]}), .y(y[518]));
  Fx519 Fx519_inst(.x({x[649], x[645]}), .y(y[519]));
  Fx520 Fx520_inst(.x({x[651], x[650]}), .y(y[520]));
  Fx521 Fx521_inst(.x({x[652], x[650]}), .y(y[521]));
  Fx522 Fx522_inst(.x({x[653], x[650]}), .y(y[522]));
  Fx523 Fx523_inst(.x({x[654], x[650]}), .y(y[523]));
  Fx524 Fx524_inst(.x({x[656], x[655]}), .y(y[524]));
  Fx525 Fx525_inst(.x({x[657], x[655]}), .y(y[525]));
  Fx526 Fx526_inst(.x({x[658], x[655]}), .y(y[526]));
  Fx527 Fx527_inst(.x({x[659], x[655]}), .y(y[527]));
  Fx528 Fx528_inst(.x({x[661], x[660]}), .y(y[528]));
  Fx529 Fx529_inst(.x({x[662], x[660]}), .y(y[529]));
  Fx530 Fx530_inst(.x({x[663], x[660]}), .y(y[530]));
  Fx531 Fx531_inst(.x({x[664], x[660]}), .y(y[531]));
  Fx532 Fx532_inst(.x({x[666], x[665]}), .y(y[532]));
  Fx533 Fx533_inst(.x({x[667], x[665]}), .y(y[533]));
  Fx534 Fx534_inst(.x({x[668], x[665]}), .y(y[534]));
  Fx535 Fx535_inst(.x({x[669], x[665]}), .y(y[535]));
  Fx536 Fx536_inst(.x({x[671], x[670]}), .y(y[536]));
  Fx537 Fx537_inst(.x({x[672], x[670]}), .y(y[537]));
  Fx538 Fx538_inst(.x({x[673], x[670]}), .y(y[538]));
  Fx539 Fx539_inst(.x({x[674], x[670]}), .y(y[539]));
endmodule

module R1ind0(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind1(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind2(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind3(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind4(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind5(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind6(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind7(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind8(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind9(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind10(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind11(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind12(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind13(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind14(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind15(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind16(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind17(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind18(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind19(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind20(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind21(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind22(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind23(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind24(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind25(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind26(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind27(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind28(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind29(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind30(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind31(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind32(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind33(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind34(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind35(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind36(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind37(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind38(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind39(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind40(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind41(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind42(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind43(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind44(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind45(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind46(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind47(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind48(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind49(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind50(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind51(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind52(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind53(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind54(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind55(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind56(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind57(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind58(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind59(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind60(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind61(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind62(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind63(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind64(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign y = t[0];
endmodule

module R1ind65(x, y);
 input [29:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[16] ^ x[29];
  assign t[11] = (x[0] & x[1] & x[2]) | (x[0] & x[1] & x[3]) | (x[0] & x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[12] = (x[5] & x[6] & x[7]) | (x[5] & x[6] & x[8]) | (x[5] & x[7] & x[8]) | (x[6] & x[7] & x[8]);
  assign t[13] = (x[10] & x[11] & x[12]) | (x[10] & x[11] & x[13]) | (x[10] & x[12] & x[13]) | (x[11] & x[12] & x[13]);
  assign t[14] = (x[15] & x[16] & x[17]) | (x[15] & x[16] & x[18]) | (x[15] & x[17] & x[18]) | (x[16] & x[17] & x[18]);
  assign t[15] = (x[20] & x[21] & x[22]) | (x[20] & x[21] & x[23]) | (x[20] & x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[16] = (x[25] & x[26] & x[27]) | (x[25] & x[26] & x[28]) | (x[25] & x[27] & x[28]) | (x[26] & x[27] & x[28]);
  assign t[1] = ~(t[5] & t[6]);
  assign t[2] = ~(t[7] | t[8]);
  assign t[3] = ~(t[9] | t[4]);
  assign t[4] = ~(t[10]);
  assign t[5] = t[11] ^ x[4];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[14];
  assign t[8] = t[14] ^ x[19];
  assign t[9] = t[15] ^ x[24];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind66(x, y);
 input [30:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[5] ? t[6] : t[1];
  assign t[10] = t[16] ^ x[30];
  assign t[11] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[12] = (x[6] & x[7] & x[8]) | (x[6] & x[7] & x[9]) | (x[6] & x[8] & x[9]) | (x[7] & x[8] & x[9]);
  assign t[13] = (x[11] & x[12] & x[13]) | (x[11] & x[12] & x[14]) | (x[11] & x[13] & x[14]) | (x[12] & x[13] & x[14]);
  assign t[14] = (x[16] & x[17] & x[18]) | (x[16] & x[17] & x[19]) | (x[16] & x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[15] = (x[21] & x[22] & x[23]) | (x[21] & x[22] & x[24]) | (x[21] & x[23] & x[24]) | (x[22] & x[23] & x[24]);
  assign t[16] = (x[26] & x[27] & x[28]) | (x[26] & x[27] & x[29]) | (x[26] & x[28] & x[29]) | (x[27] & x[28] & x[29]);
  assign t[1] = ~(t[6] & t[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = t[7] & t[8];
  assign t[4] = ~(t[9] | t[10]);
  assign t[5] = t[11] ^ x[5];
  assign t[6] = t[12] ^ x[10];
  assign t[7] = t[13] ^ x[15];
  assign t[8] = t[14] ^ x[20];
  assign t[9] = t[15] ^ x[25];
  assign y = ~(~x[0] & ~t[0]);
endmodule

module R1ind67(x, y);
 input [5:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind68(x, y);
 input [30:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] & t[5];
  assign t[10] = t[16] ^ x[30];
  assign t[11] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[12] = (x[6] & x[7] & x[8]) | (x[6] & x[7] & x[9]) | (x[6] & x[8] & x[9]) | (x[7] & x[8] & x[9]);
  assign t[13] = (x[11] & x[12] & x[13]) | (x[11] & x[12] & x[14]) | (x[11] & x[13] & x[14]) | (x[12] & x[13] & x[14]);
  assign t[14] = (x[16] & x[17] & x[18]) | (x[16] & x[17] & x[19]) | (x[16] & x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[15] = (x[21] & x[22] & x[23]) | (x[21] & x[22] & x[24]) | (x[21] & x[23] & x[24]) | (x[22] & x[23] & x[24]);
  assign t[16] = (x[26] & x[27] & x[28]) | (x[26] & x[27] & x[29]) | (x[26] & x[28] & x[29]) | (x[27] & x[28] & x[29]);
  assign t[1] = ~(t[2] & t[6]);
  assign t[2] = ~(t[7] | t[3]);
  assign t[3] = ~(t[8] & t[4]);
  assign t[4] = ~(t[9] | t[10]);
  assign t[5] = t[11] ^ x[5];
  assign t[6] = t[12] ^ x[10];
  assign t[7] = t[13] ^ x[15];
  assign t[8] = t[14] ^ x[20];
  assign t[9] = t[15] ^ x[25];
  assign y = ~x[0] & t[0];
endmodule

module R1ind69(x, y);
 input [5:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind70(x, y);
 input [5:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind71(x, y);
 input [30:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[5] | t[1];
  assign t[10] = t[16] ^ x[30];
  assign t[11] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[12] = (x[6] & x[7] & x[8]) | (x[6] & x[7] & x[9]) | (x[6] & x[8] & x[9]) | (x[7] & x[8] & x[9]);
  assign t[13] = (x[11] & x[12] & x[13]) | (x[11] & x[12] & x[14]) | (x[11] & x[13] & x[14]) | (x[12] & x[13] & x[14]);
  assign t[14] = (x[16] & x[17] & x[18]) | (x[16] & x[17] & x[19]) | (x[16] & x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[15] = (x[21] & x[22] & x[23]) | (x[21] & x[22] & x[24]) | (x[21] & x[23] & x[24]) | (x[22] & x[23] & x[24]);
  assign t[16] = (x[26] & x[27] & x[28]) | (x[26] & x[27] & x[29]) | (x[26] & x[28] & x[29]) | (x[27] & x[28] & x[29]);
  assign t[1] = ~(t[6] | t[2]);
  assign t[2] = ~(t[7] & t[3]);
  assign t[3] = ~(t[8] | t[4]);
  assign t[4] = ~(t[9] & t[10]);
  assign t[5] = t[11] ^ x[5];
  assign t[6] = t[12] ^ x[10];
  assign t[7] = t[13] ^ x[15];
  assign t[8] = t[14] ^ x[20];
  assign t[9] = t[15] ^ x[25];
  assign y = ~x[0] & t[0];
endmodule

module R1ind72(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind73(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind74(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind75(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind76(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind77(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind78(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind79(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind80(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind81(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind82(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind83(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind84(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind85(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind86(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind87(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind88(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind89(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind90(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind91(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind92(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind93(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind94(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind95(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind96(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind97(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind98(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind99(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind100(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind101(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind102(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind103(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind104(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind105(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind106(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind107(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind108(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind109(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind110(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind111(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind112(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind113(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind114(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind115(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind116(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind117(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind118(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind119(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind120(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind121(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind122(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind123(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind124(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind125(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind126(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind127(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind128(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind129(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind130(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind131(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind132(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind133(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind134(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind135(x, y);
 input [6:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[1] = (x[1] & x[2] & x[3]) | (x[1] & x[2] & x[4]) | (x[1] & x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign y = x[0] ? x[6] : t[0];
endmodule

module R1ind136(x, y);
 input [46:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[6];
  assign t[37] = t[46] ^ x[11];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[26];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = t[51] ^ x[36];
  assign t[43] = t[52] ^ x[41];
  assign t[44] = t[53] ^ x[46];
  assign t[45] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[46] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[47] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[48] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[49] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[51] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[52] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[53] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind137(x, y);
 input [46:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[37] ^ t[14];
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[12] = t[38] ^ t[39];
  assign t[13] = t[14] & t[19];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[37] ^ t[14]);
  assign t[16] = t[37] & t[20];
  assign t[17] = t[21] ^ t[22];
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[37] ^ t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[13];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[40] ^ t[29];
  assign t[25] = t[39] ^ t[41];
  assign t[26] = t[37] ^ t[12];
  assign t[27] = t[42] ^ t[43];
  assign t[28] = t[29] & t[32];
  assign t[29] = ~(t[43]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[40] ^ t[29]);
  assign t[31] = t[40] & t[33];
  assign t[32] = t[40] ^ t[34];
  assign t[33] = t[35] ^ t[28];
  assign t[34] = t[43] ^ t[44];
  assign t[35] = t[40] ^ t[27];
  assign t[36] = t[45] ^ x[6];
  assign t[37] = t[46] ^ x[11];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[26];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = t[51] ^ x[36];
  assign t[43] = t[52] ^ x[41];
  assign t[44] = t[53] ^ x[46];
  assign t[45] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[46] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[47] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[48] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[49] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[51] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[52] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[53] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind138(x, y);
 input [36:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[16];
  assign t[19] = t[26] ^ x[21];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[26];
  assign t[21] = t[28] ^ x[31];
  assign t[22] = t[29] ^ x[36];
  assign t[23] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[24] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[25] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[26] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[27] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[28] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[29] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind139(x, y);
 input [46:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[6];
  assign t[25] = t[34] ^ x[11];
  assign t[26] = t[35] ^ x[16];
  assign t[27] = t[36] ^ x[21];
  assign t[28] = t[37] ^ x[26];
  assign t[29] = t[38] ^ x[31];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[36];
  assign t[31] = t[40] ^ x[41];
  assign t[32] = t[41] ^ x[46];
  assign t[33] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[34] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[35] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[36] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[37] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[38] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[39] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[41] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind140(x, y);
 input [46:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[6];
  assign t[37] = t[46] ^ x[11];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[26];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = t[51] ^ x[36];
  assign t[43] = t[52] ^ x[41];
  assign t[44] = t[53] ^ x[46];
  assign t[45] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[46] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[47] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[48] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[49] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[51] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[52] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[53] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind141(x, y);
 input [46:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[17] & t[18];
  assign t[11] = t[19] ^ t[10];
  assign t[12] = t[38] ^ t[17];
  assign t[13] = t[20] ^ t[21];
  assign t[14] = t[22] ^ t[23];
  assign t[15] = t[39] ^ t[40];
  assign t[16] = t[17] & t[24];
  assign t[17] = ~(t[40]);
  assign t[18] = ~(t[38] ^ t[17]);
  assign t[19] = t[38] & t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[27];
  assign t[21] = t[28] & t[29];
  assign t[22] = t[30] ^ t[21];
  assign t[23] = t[41] ^ t[28];
  assign t[24] = t[38] ^ t[31];
  assign t[25] = t[32] ^ t[16];
  assign t[26] = t[42] ^ t[43];
  assign t[27] = t[28] & t[33];
  assign t[28] = ~(t[43]);
  assign t[29] = ~(t[41] ^ t[28]);
  assign t[2] = ~(t[4]);
  assign t[30] = t[41] & t[34];
  assign t[31] = t[40] ^ t[44];
  assign t[32] = t[38] ^ t[15];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[27];
  assign t[35] = t[43] ^ t[45];
  assign t[36] = t[41] ^ t[26];
  assign t[37] = t[46] ^ x[6];
  assign t[38] = t[47] ^ x[11];
  assign t[39] = t[48] ^ x[16];
  assign t[3] = ~(t[5] ^ t[37]);
  assign t[40] = t[49] ^ x[21];
  assign t[41] = t[50] ^ x[26];
  assign t[42] = t[51] ^ x[31];
  assign t[43] = t[52] ^ x[36];
  assign t[44] = t[53] ^ x[41];
  assign t[45] = t[54] ^ x[46];
  assign t[46] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[47] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[48] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[49] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[4] = ~(t[6] ^ t[7]);
  assign t[50] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[51] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[52] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[53] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[54] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] ^ t[12];
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[9] = t[15] ^ t[16];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind142(x, y);
 input [36:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[16];
  assign t[19] = t[26] ^ x[21];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[26];
  assign t[21] = t[28] ^ x[31];
  assign t[22] = t[29] ^ x[36];
  assign t[23] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[24] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[25] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[26] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[27] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[28] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[29] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind143(x, y);
 input [46:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[6];
  assign t[25] = t[34] ^ x[11];
  assign t[26] = t[35] ^ x[16];
  assign t[27] = t[36] ^ x[21];
  assign t[28] = t[37] ^ x[26];
  assign t[29] = t[38] ^ x[31];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[36];
  assign t[31] = t[40] ^ x[41];
  assign t[32] = t[41] ^ x[46];
  assign t[33] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[34] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[35] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[36] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[37] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[38] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[39] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[41] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind144(x, y);
 input [46:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[6];
  assign t[37] = t[46] ^ x[11];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[26];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = t[51] ^ x[36];
  assign t[43] = t[52] ^ x[41];
  assign t[44] = t[53] ^ x[46];
  assign t[45] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[46] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[47] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[48] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[49] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[51] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[52] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[53] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind145(x, y);
 input [46:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[37] ^ t[14];
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[12] = t[38] ^ t[39];
  assign t[13] = t[14] & t[19];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[37] ^ t[14]);
  assign t[16] = t[37] & t[20];
  assign t[17] = t[21] ^ t[22];
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[37] ^ t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[13];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[40] ^ t[29];
  assign t[25] = t[39] ^ t[41];
  assign t[26] = t[37] ^ t[12];
  assign t[27] = t[42] ^ t[43];
  assign t[28] = t[29] & t[32];
  assign t[29] = ~(t[43]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[40] ^ t[29]);
  assign t[31] = t[40] & t[33];
  assign t[32] = t[40] ^ t[34];
  assign t[33] = t[35] ^ t[28];
  assign t[34] = t[43] ^ t[44];
  assign t[35] = t[40] ^ t[27];
  assign t[36] = t[45] ^ x[6];
  assign t[37] = t[46] ^ x[11];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[26];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = t[51] ^ x[36];
  assign t[43] = t[52] ^ x[41];
  assign t[44] = t[53] ^ x[46];
  assign t[45] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[46] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[47] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[48] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[49] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[51] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[52] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[53] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind146(x, y);
 input [36:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[16];
  assign t[19] = t[26] ^ x[21];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[26];
  assign t[21] = t[28] ^ x[31];
  assign t[22] = t[29] ^ x[36];
  assign t[23] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[24] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[25] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[26] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[27] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[28] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[29] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind147(x, y);
 input [46:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[6];
  assign t[25] = t[34] ^ x[11];
  assign t[26] = t[35] ^ x[16];
  assign t[27] = t[36] ^ x[21];
  assign t[28] = t[37] ^ x[26];
  assign t[29] = t[38] ^ x[31];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[36];
  assign t[31] = t[40] ^ x[41];
  assign t[32] = t[41] ^ x[46];
  assign t[33] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[34] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[35] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[36] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[37] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[38] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[39] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[41] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind148(x, y);
 input [51:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = ~(t[17] ^ t[40]);
  assign t[12] = t[18] ^ t[19];
  assign t[13] = ~(t[41]);
  assign t[14] = ~(t[39] ^ t[13]);
  assign t[15] = t[42] ^ t[41];
  assign t[16] = ~(t[20] ^ t[9]);
  assign t[17] = ~t[21];
  assign t[18] = t[39] ^ t[15];
  assign t[19] = t[13] & t[20];
  assign t[1] = ~t[3];
  assign t[20] = t[39] ^ t[22];
  assign t[21] = t[23] ^ t[24];
  assign t[22] = t[41] ^ t[43];
  assign t[23] = t[25] ^ t[26];
  assign t[24] = t[27] & t[28];
  assign t[25] = t[44] & t[29];
  assign t[26] = t[30] & t[31];
  assign t[27] = t[32] ^ t[30];
  assign t[28] = t[33] ^ t[26];
  assign t[29] = t[34] ^ t[35];
  assign t[2] = t[4] ^ t[5];
  assign t[30] = ~(t[45]);
  assign t[31] = ~(t[44] ^ t[30]);
  assign t[32] = t[46] ^ t[45];
  assign t[33] = ~(t[36] ^ t[27]);
  assign t[34] = t[44] ^ t[32];
  assign t[35] = t[30] & t[36];
  assign t[36] = t[44] ^ t[37];
  assign t[37] = t[45] ^ t[47];
  assign t[38] = t[48] ^ x[6];
  assign t[39] = t[49] ^ x[11];
  assign t[3] = ~(t[6] ^ t[38]);
  assign t[40] = t[50] ^ x[16];
  assign t[41] = t[51] ^ x[21];
  assign t[42] = t[52] ^ x[26];
  assign t[43] = t[53] ^ x[31];
  assign t[44] = t[54] ^ x[36];
  assign t[45] = t[55] ^ x[41];
  assign t[46] = t[56] ^ x[46];
  assign t[47] = t[57] ^ x[51];
  assign t[48] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[49] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[51] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[52] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[53] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[54] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[55] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[56] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[57] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[39] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind149(x, y);
 input [51:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[39] ^ t[14];
  assign t[11] = ~(t[17] ^ t[40]);
  assign t[12] = t[41] ^ t[42];
  assign t[13] = t[14] & t[18];
  assign t[14] = ~(t[42]);
  assign t[15] = ~(t[39] ^ t[14]);
  assign t[16] = t[39] & t[19];
  assign t[17] = ~t[20];
  assign t[18] = t[39] ^ t[21];
  assign t[19] = t[22] ^ t[13];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23] ^ t[24]);
  assign t[21] = t[42] ^ t[43];
  assign t[22] = t[39] ^ t[12];
  assign t[23] = t[25] ^ t[26];
  assign t[24] = t[27] ^ t[28];
  assign t[25] = t[29] ^ t[30];
  assign t[26] = t[31] & t[32];
  assign t[27] = t[33] ^ t[26];
  assign t[28] = t[44] ^ t[31];
  assign t[29] = t[45] ^ t[46];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[31] & t[34];
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[44] ^ t[31]);
  assign t[33] = t[44] & t[35];
  assign t[34] = t[44] ^ t[36];
  assign t[35] = t[37] ^ t[30];
  assign t[36] = t[46] ^ t[47];
  assign t[37] = t[44] ^ t[29];
  assign t[38] = t[48] ^ x[6];
  assign t[39] = t[49] ^ x[11];
  assign t[3] = ~(t[6] ^ t[38]);
  assign t[40] = t[50] ^ x[16];
  assign t[41] = t[51] ^ x[21];
  assign t[42] = t[52] ^ x[26];
  assign t[43] = t[53] ^ x[31];
  assign t[44] = t[54] ^ x[36];
  assign t[45] = t[55] ^ x[41];
  assign t[46] = t[56] ^ x[46];
  assign t[47] = t[57] ^ x[51];
  assign t[48] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[49] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[51] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[52] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[53] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[54] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[55] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[56] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[57] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind150(x, y);
 input [41:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[22] ^ t[9]);
  assign t[11] = ~t[12];
  assign t[12] = ~(t[13]);
  assign t[13] = t[14] ^ t[15];
  assign t[14] = t[23] ^ t[24];
  assign t[15] = t[16] & t[17];
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[25] ^ t[16]);
  assign t[18] = t[26] ^ x[6];
  assign t[19] = t[27] ^ x[11];
  assign t[1] = ~t[3];
  assign t[20] = t[28] ^ x[16];
  assign t[21] = t[29] ^ x[21];
  assign t[22] = t[30] ^ x[26];
  assign t[23] = t[31] ^ x[31];
  assign t[24] = t[32] ^ x[36];
  assign t[25] = t[33] ^ x[41];
  assign t[26] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[27] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[28] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[29] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[2] = ~(t[4]);
  assign t[30] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[31] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[32] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[33] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[3] = ~(t[5] ^ t[18]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[19] ^ t[20];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11] ^ t[21]);
  assign t[9] = ~(t[19]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind151(x, y);
 input [51:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[29]);
  assign t[12] = ~(t[30] ^ t[11]);
  assign t[13] = ~t[15];
  assign t[14] = t[30] ^ t[16];
  assign t[15] = ~(t[17]);
  assign t[16] = t[29] ^ t[31];
  assign t[17] = t[18] ^ t[19];
  assign t[18] = t[20] ^ t[21];
  assign t[19] = t[22] & t[23];
  assign t[1] = ~t[3];
  assign t[20] = t[32] ^ t[33];
  assign t[21] = t[22] & t[24];
  assign t[22] = ~(t[33]);
  assign t[23] = ~(t[34] ^ t[22]);
  assign t[24] = t[34] ^ t[25];
  assign t[25] = t[33] ^ t[35];
  assign t[26] = t[36] ^ x[6];
  assign t[27] = t[37] ^ x[11];
  assign t[28] = t[38] ^ x[16];
  assign t[29] = t[39] ^ x[21];
  assign t[2] = ~(t[4]);
  assign t[30] = t[40] ^ x[26];
  assign t[31] = t[41] ^ x[31];
  assign t[32] = t[42] ^ x[36];
  assign t[33] = t[43] ^ x[41];
  assign t[34] = t[44] ^ x[46];
  assign t[35] = t[45] ^ x[51];
  assign t[36] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[37] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[38] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[39] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[3] = ~(t[5] ^ t[26]);
  assign t[40] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[41] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[42] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[43] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[44] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[45] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13] ^ t[27]);
  assign t[9] = t[28] ^ t[29];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind152(x, y);
 input [46:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[6];
  assign t[37] = t[46] ^ x[11];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[26];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = t[51] ^ x[36];
  assign t[43] = t[52] ^ x[41];
  assign t[44] = t[53] ^ x[46];
  assign t[45] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[46] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[47] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[48] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[49] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[51] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[52] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[53] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind153(x, y);
 input [46:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[37] ^ t[14];
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[12] = t[38] ^ t[39];
  assign t[13] = t[14] & t[19];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[37] ^ t[14]);
  assign t[16] = t[37] & t[20];
  assign t[17] = t[21] ^ t[22];
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[37] ^ t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[13];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[40] ^ t[29];
  assign t[25] = t[39] ^ t[41];
  assign t[26] = t[37] ^ t[12];
  assign t[27] = t[42] ^ t[43];
  assign t[28] = t[29] & t[32];
  assign t[29] = ~(t[43]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[40] ^ t[29]);
  assign t[31] = t[40] & t[33];
  assign t[32] = t[40] ^ t[34];
  assign t[33] = t[35] ^ t[28];
  assign t[34] = t[43] ^ t[44];
  assign t[35] = t[40] ^ t[27];
  assign t[36] = t[45] ^ x[6];
  assign t[37] = t[46] ^ x[11];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[26];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = t[51] ^ x[36];
  assign t[43] = t[52] ^ x[41];
  assign t[44] = t[53] ^ x[46];
  assign t[45] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[46] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[47] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[48] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[49] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[51] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[52] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[53] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind154(x, y);
 input [36:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[16];
  assign t[19] = t[26] ^ x[21];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[26];
  assign t[21] = t[28] ^ x[31];
  assign t[22] = t[29] ^ x[36];
  assign t[23] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[24] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[25] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[26] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[27] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[28] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[29] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind155(x, y);
 input [46:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[6];
  assign t[25] = t[34] ^ x[11];
  assign t[26] = t[35] ^ x[16];
  assign t[27] = t[36] ^ x[21];
  assign t[28] = t[37] ^ x[26];
  assign t[29] = t[38] ^ x[31];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[36];
  assign t[31] = t[40] ^ x[41];
  assign t[32] = t[41] ^ x[46];
  assign t[33] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[34] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[35] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[36] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[37] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[38] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[39] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[41] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind156(x, y);
 input [46:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[6];
  assign t[37] = t[46] ^ x[11];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[26];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = t[51] ^ x[36];
  assign t[43] = t[52] ^ x[41];
  assign t[44] = t[53] ^ x[46];
  assign t[45] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[46] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[47] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[48] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[49] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[51] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[52] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[53] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind157(x, y);
 input [46:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[17] & t[18];
  assign t[11] = t[19] ^ t[10];
  assign t[12] = t[38] ^ t[17];
  assign t[13] = t[20] ^ t[21];
  assign t[14] = t[22] ^ t[23];
  assign t[15] = t[39] ^ t[40];
  assign t[16] = t[17] & t[24];
  assign t[17] = ~(t[40]);
  assign t[18] = ~(t[38] ^ t[17]);
  assign t[19] = t[38] & t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[27];
  assign t[21] = t[28] & t[29];
  assign t[22] = t[30] ^ t[21];
  assign t[23] = t[41] ^ t[28];
  assign t[24] = t[38] ^ t[31];
  assign t[25] = t[32] ^ t[16];
  assign t[26] = t[42] ^ t[43];
  assign t[27] = t[28] & t[33];
  assign t[28] = ~(t[43]);
  assign t[29] = ~(t[41] ^ t[28]);
  assign t[2] = ~(t[4]);
  assign t[30] = t[41] & t[34];
  assign t[31] = t[40] ^ t[44];
  assign t[32] = t[38] ^ t[15];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[27];
  assign t[35] = t[43] ^ t[45];
  assign t[36] = t[41] ^ t[26];
  assign t[37] = t[46] ^ x[6];
  assign t[38] = t[47] ^ x[11];
  assign t[39] = t[48] ^ x[16];
  assign t[3] = ~(t[5] ^ t[37]);
  assign t[40] = t[49] ^ x[21];
  assign t[41] = t[50] ^ x[26];
  assign t[42] = t[51] ^ x[31];
  assign t[43] = t[52] ^ x[36];
  assign t[44] = t[53] ^ x[41];
  assign t[45] = t[54] ^ x[46];
  assign t[46] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[47] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[48] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[49] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[4] = ~(t[6] ^ t[7]);
  assign t[50] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[51] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[52] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[53] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[54] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] ^ t[12];
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[9] = t[15] ^ t[16];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind158(x, y);
 input [36:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[16];
  assign t[19] = t[26] ^ x[21];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[26];
  assign t[21] = t[28] ^ x[31];
  assign t[22] = t[29] ^ x[36];
  assign t[23] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[24] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[25] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[26] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[27] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[28] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[29] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind159(x, y);
 input [46:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[6];
  assign t[25] = t[34] ^ x[11];
  assign t[26] = t[35] ^ x[16];
  assign t[27] = t[36] ^ x[21];
  assign t[28] = t[37] ^ x[26];
  assign t[29] = t[38] ^ x[31];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[36];
  assign t[31] = t[40] ^ x[41];
  assign t[32] = t[41] ^ x[46];
  assign t[33] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[34] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[35] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[36] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[37] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[38] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[39] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[41] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind160(x, y);
 input [51:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = ~(t[17] ^ t[40]);
  assign t[12] = t[18] ^ t[19];
  assign t[13] = ~(t[41]);
  assign t[14] = ~(t[39] ^ t[13]);
  assign t[15] = t[42] ^ t[41];
  assign t[16] = ~(t[20] ^ t[9]);
  assign t[17] = ~t[21];
  assign t[18] = t[39] ^ t[15];
  assign t[19] = t[13] & t[20];
  assign t[1] = ~t[3];
  assign t[20] = t[39] ^ t[22];
  assign t[21] = t[23] ^ t[24];
  assign t[22] = t[41] ^ t[43];
  assign t[23] = t[25] ^ t[26];
  assign t[24] = t[27] & t[28];
  assign t[25] = t[44] & t[29];
  assign t[26] = t[30] & t[31];
  assign t[27] = t[32] ^ t[30];
  assign t[28] = t[33] ^ t[26];
  assign t[29] = t[34] ^ t[35];
  assign t[2] = t[4] ^ t[5];
  assign t[30] = ~(t[45]);
  assign t[31] = ~(t[44] ^ t[30]);
  assign t[32] = t[46] ^ t[45];
  assign t[33] = ~(t[36] ^ t[27]);
  assign t[34] = t[44] ^ t[32];
  assign t[35] = t[30] & t[36];
  assign t[36] = t[44] ^ t[37];
  assign t[37] = t[45] ^ t[47];
  assign t[38] = t[48] ^ x[6];
  assign t[39] = t[49] ^ x[11];
  assign t[3] = ~(t[6] ^ t[38]);
  assign t[40] = t[50] ^ x[16];
  assign t[41] = t[51] ^ x[21];
  assign t[42] = t[52] ^ x[26];
  assign t[43] = t[53] ^ x[31];
  assign t[44] = t[54] ^ x[36];
  assign t[45] = t[55] ^ x[41];
  assign t[46] = t[56] ^ x[46];
  assign t[47] = t[57] ^ x[51];
  assign t[48] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[49] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[51] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[52] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[53] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[54] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[55] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[56] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[57] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[39] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind161(x, y);
 input [51:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[39] ^ t[14];
  assign t[11] = ~(t[17] ^ t[40]);
  assign t[12] = t[41] ^ t[42];
  assign t[13] = t[14] & t[18];
  assign t[14] = ~(t[42]);
  assign t[15] = ~(t[39] ^ t[14]);
  assign t[16] = t[39] & t[19];
  assign t[17] = ~t[20];
  assign t[18] = t[39] ^ t[21];
  assign t[19] = t[22] ^ t[13];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23] ^ t[24]);
  assign t[21] = t[42] ^ t[43];
  assign t[22] = t[39] ^ t[12];
  assign t[23] = t[25] ^ t[26];
  assign t[24] = t[27] ^ t[28];
  assign t[25] = t[29] ^ t[30];
  assign t[26] = t[31] & t[32];
  assign t[27] = t[33] ^ t[26];
  assign t[28] = t[44] ^ t[31];
  assign t[29] = t[45] ^ t[46];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[31] & t[34];
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[44] ^ t[31]);
  assign t[33] = t[44] & t[35];
  assign t[34] = t[44] ^ t[36];
  assign t[35] = t[37] ^ t[30];
  assign t[36] = t[46] ^ t[47];
  assign t[37] = t[44] ^ t[29];
  assign t[38] = t[48] ^ x[6];
  assign t[39] = t[49] ^ x[11];
  assign t[3] = ~(t[6] ^ t[38]);
  assign t[40] = t[50] ^ x[16];
  assign t[41] = t[51] ^ x[21];
  assign t[42] = t[52] ^ x[26];
  assign t[43] = t[53] ^ x[31];
  assign t[44] = t[54] ^ x[36];
  assign t[45] = t[55] ^ x[41];
  assign t[46] = t[56] ^ x[46];
  assign t[47] = t[57] ^ x[51];
  assign t[48] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[49] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[51] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[52] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[53] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[54] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[55] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[56] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[57] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind162(x, y);
 input [36:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[21] ^ t[9]);
  assign t[11] = ~t[12];
  assign t[12] = ~(t[13]);
  assign t[13] = t[14] ^ t[15];
  assign t[14] = t[22] ^ t[23];
  assign t[15] = t[16] & t[17];
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[24] ^ t[16]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[16];
  assign t[21] = t[28] ^ x[21];
  assign t[22] = t[29] ^ x[26];
  assign t[23] = t[30] ^ x[31];
  assign t[24] = t[31] ^ x[36];
  assign t[25] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[26] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[27] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[28] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[29] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[2] = ~(t[4]);
  assign t[30] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[31] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[3] = ~(t[5] ^ t[18]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[19] ^ t[20];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~t[11];
  assign t[9] = ~(t[19]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind163(x, y);
 input [46:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[28]);
  assign t[12] = ~(t[29] ^ t[11]);
  assign t[13] = ~t[15];
  assign t[14] = t[29] ^ t[16];
  assign t[15] = ~(t[17]);
  assign t[16] = t[28] ^ t[30];
  assign t[17] = t[18] ^ t[19];
  assign t[18] = t[20] ^ t[21];
  assign t[19] = t[22] & t[23];
  assign t[1] = ~t[3];
  assign t[20] = t[31] ^ t[32];
  assign t[21] = t[22] & t[24];
  assign t[22] = ~(t[32]);
  assign t[23] = ~(t[33] ^ t[22]);
  assign t[24] = t[33] ^ t[25];
  assign t[25] = t[32] ^ t[34];
  assign t[26] = t[35] ^ x[6];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[16];
  assign t[29] = t[38] ^ x[21];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[26];
  assign t[31] = t[40] ^ x[31];
  assign t[32] = t[41] ^ x[36];
  assign t[33] = t[42] ^ x[41];
  assign t[34] = t[43] ^ x[46];
  assign t[35] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[36] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[37] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[38] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[39] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[3] = ~(t[5] ^ t[26]);
  assign t[40] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[41] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[42] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[43] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~t[13];
  assign t[9] = t[27] ^ t[28];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind164(x, y);
 input [46:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[6];
  assign t[37] = t[46] ^ x[11];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[26];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = t[51] ^ x[36];
  assign t[43] = t[52] ^ x[41];
  assign t[44] = t[53] ^ x[46];
  assign t[45] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[46] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[47] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[48] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[49] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[51] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[52] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[53] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind165(x, y);
 input [46:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[37] ^ t[14];
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[12] = t[38] ^ t[39];
  assign t[13] = t[14] & t[19];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[37] ^ t[14]);
  assign t[16] = t[37] & t[20];
  assign t[17] = t[21] ^ t[22];
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[37] ^ t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[13];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[40] ^ t[29];
  assign t[25] = t[39] ^ t[41];
  assign t[26] = t[37] ^ t[12];
  assign t[27] = t[42] ^ t[43];
  assign t[28] = t[29] & t[32];
  assign t[29] = ~(t[43]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[40] ^ t[29]);
  assign t[31] = t[40] & t[33];
  assign t[32] = t[40] ^ t[34];
  assign t[33] = t[35] ^ t[28];
  assign t[34] = t[43] ^ t[44];
  assign t[35] = t[40] ^ t[27];
  assign t[36] = t[45] ^ x[6];
  assign t[37] = t[46] ^ x[11];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[26];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = t[51] ^ x[36];
  assign t[43] = t[52] ^ x[41];
  assign t[44] = t[53] ^ x[46];
  assign t[45] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[46] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[47] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[48] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[49] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[51] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[52] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[53] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind166(x, y);
 input [36:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[16];
  assign t[19] = t[26] ^ x[21];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[26];
  assign t[21] = t[28] ^ x[31];
  assign t[22] = t[29] ^ x[36];
  assign t[23] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[24] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[25] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[26] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[27] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[28] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[29] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind167(x, y);
 input [46:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[6];
  assign t[25] = t[34] ^ x[11];
  assign t[26] = t[35] ^ x[16];
  assign t[27] = t[36] ^ x[21];
  assign t[28] = t[37] ^ x[26];
  assign t[29] = t[38] ^ x[31];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[36];
  assign t[31] = t[40] ^ x[41];
  assign t[32] = t[41] ^ x[46];
  assign t[33] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[34] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[35] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[36] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[37] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[38] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[39] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[41] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind168(x, y);
 input [26:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[24] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[25] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[26] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[27] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind169(x, y);
 input [26:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[24] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[25] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[26] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[27] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind170(x, y);
 input [21:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = t[14] ^ x[16];
  assign t[11] = t[15] ^ x[21];
  assign t[12] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[13] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[14] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[15] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[1] = ~t[2];
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind171(x, y);
 input [26:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = t[17] ^ x[6];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[16];
  assign t[15] = t[20] ^ x[21];
  assign t[16] = t[21] ^ x[26];
  assign t[17] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[18] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[19] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[1] = ~t[2];
  assign t[20] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[21] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind172(x, y);
 input [26:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[24] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[25] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[26] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[27] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind173(x, y);
 input [26:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[24] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[25] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[26] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[27] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind174(x, y);
 input [21:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = t[14] ^ x[16];
  assign t[11] = t[15] ^ x[21];
  assign t[12] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[13] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[14] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[15] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[1] = ~t[2];
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind175(x, y);
 input [26:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = t[17] ^ x[6];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[16];
  assign t[15] = t[20] ^ x[21];
  assign t[16] = t[21] ^ x[26];
  assign t[17] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[18] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[19] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[1] = ~t[2];
  assign t[20] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[21] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind176(x, y);
 input [26:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[24] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[25] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[26] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[27] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind177(x, y);
 input [26:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[24] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[25] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[26] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[27] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind178(x, y);
 input [21:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = t[14] ^ x[16];
  assign t[11] = t[15] ^ x[21];
  assign t[12] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[13] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[14] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[15] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[1] = ~t[2];
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind179(x, y);
 input [26:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = t[17] ^ x[6];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[16];
  assign t[15] = t[20] ^ x[21];
  assign t[16] = t[21] ^ x[26];
  assign t[17] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[18] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[19] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[1] = ~t[2];
  assign t[20] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[21] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind180(x, y);
 input [31:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[20]);
  assign t[10] = t[15] ^ t[8];
  assign t[11] = t[16] ^ t[17];
  assign t[12] = ~(t[23]);
  assign t[13] = ~(t[22] ^ t[12]);
  assign t[14] = t[24] ^ t[23];
  assign t[15] = ~(t[18] ^ t[9]);
  assign t[16] = t[22] ^ t[14];
  assign t[17] = t[12] & t[18];
  assign t[18] = t[22] ^ t[19];
  assign t[19] = t[23] ^ t[25];
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[11];
  assign t[22] = t[28] ^ x[16];
  assign t[23] = t[29] ^ x[21];
  assign t[24] = t[30] ^ x[26];
  assign t[25] = t[31] ^ x[31];
  assign t[26] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[27] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[28] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[29] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[2] = ~(t[3] ^ t[21]);
  assign t[30] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[31] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[3] = ~t[4];
  assign t[4] = t[5] ^ t[6];
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] & t[10];
  assign t[7] = t[22] & t[11];
  assign t[8] = t[12] & t[13];
  assign t[9] = t[14] ^ t[12];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind181(x, y);
 input [31:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[20]);
  assign t[10] = t[22] ^ t[13];
  assign t[11] = t[23] ^ t[24];
  assign t[12] = t[13] & t[16];
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[22] ^ t[13]);
  assign t[15] = t[22] & t[17];
  assign t[16] = t[22] ^ t[18];
  assign t[17] = t[19] ^ t[12];
  assign t[18] = t[24] ^ t[25];
  assign t[19] = t[22] ^ t[11];
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[6];
  assign t[21] = t[27] ^ x[11];
  assign t[22] = t[28] ^ x[16];
  assign t[23] = t[29] ^ x[21];
  assign t[24] = t[30] ^ x[26];
  assign t[25] = t[31] ^ x[31];
  assign t[26] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[27] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[28] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[29] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[2] = ~(t[3] ^ t[21]);
  assign t[30] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[31] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[3] = ~t[4];
  assign t[4] = ~(t[5] ^ t[6]);
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] ^ t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind182(x, y);
 input [26:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~(t[1] ^ t[10]);
  assign t[10] = t[15] ^ x[6];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[16];
  assign t[13] = t[18] ^ x[21];
  assign t[14] = t[19] ^ x[26];
  assign t[15] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[16] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[17] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[18] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[19] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[1] = ~t[2];
  assign t[2] = ~(t[3] ^ t[11]);
  assign t[3] = ~t[4];
  assign t[4] = ~(t[5]);
  assign t[5] = t[6] ^ t[7];
  assign t[6] = t[12] ^ t[13];
  assign t[7] = t[8] & t[9];
  assign t[8] = ~(t[12]);
  assign t[9] = ~(t[14] ^ t[8]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind183(x, y);
 input [31:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = ~(t[1] ^ t[14]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18] ^ t[10]);
  assign t[12] = t[18] ^ t[13];
  assign t[13] = t[17] ^ t[19];
  assign t[14] = t[20] ^ x[6];
  assign t[15] = t[21] ^ x[11];
  assign t[16] = t[22] ^ x[16];
  assign t[17] = t[23] ^ x[21];
  assign t[18] = t[24] ^ x[26];
  assign t[19] = t[25] ^ x[31];
  assign t[1] = ~t[2];
  assign t[20] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[21] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[22] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[23] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[24] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[25] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[2] = ~(t[3] ^ t[15]);
  assign t[3] = ~t[4];
  assign t[4] = ~(t[5]);
  assign t[5] = t[6] ^ t[7];
  assign t[6] = t[8] ^ t[9];
  assign t[7] = t[10] & t[11];
  assign t[8] = t[16] ^ t[17];
  assign t[9] = t[10] & t[12];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind184(x, y);
 input [66:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[19] & t[20];
  assign t[11] = t[21] ^ t[22];
  assign t[12] = t[23] & t[24];
  assign t[13] = t[53] & t[25];
  assign t[14] = t[26] & t[27];
  assign t[15] = t[28] ^ t[26];
  assign t[16] = t[29] ^ t[14];
  assign t[17] = t[54] & t[30];
  assign t[18] = t[31] & t[32];
  assign t[19] = t[33] ^ t[31];
  assign t[1] = ~(t[3] ^ t[52]);
  assign t[20] = t[34] ^ t[18];
  assign t[21] = t[55] & t[35];
  assign t[22] = t[36] & t[37];
  assign t[23] = t[38] ^ t[36];
  assign t[24] = t[39] ^ t[22];
  assign t[25] = t[40] ^ t[41];
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[53] ^ t[26]);
  assign t[28] = t[57] ^ t[56];
  assign t[29] = ~(t[42] ^ t[15]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[44];
  assign t[31] = ~(t[58]);
  assign t[32] = ~(t[54] ^ t[31]);
  assign t[33] = t[59] ^ t[58];
  assign t[34] = ~(t[45] ^ t[19]);
  assign t[35] = t[46] ^ t[47];
  assign t[36] = ~(t[60]);
  assign t[37] = ~(t[55] ^ t[36]);
  assign t[38] = t[61] ^ t[60];
  assign t[39] = ~(t[48] ^ t[23]);
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ t[28];
  assign t[41] = t[26] & t[42];
  assign t[42] = t[53] ^ t[49];
  assign t[43] = t[54] ^ t[33];
  assign t[44] = t[31] & t[45];
  assign t[45] = t[54] ^ t[50];
  assign t[46] = t[55] ^ t[38];
  assign t[47] = t[36] & t[48];
  assign t[48] = t[55] ^ t[51];
  assign t[49] = t[56] ^ t[62];
  assign t[4] = t[7] ^ t[8];
  assign t[50] = t[58] ^ t[63];
  assign t[51] = t[60] ^ t[64];
  assign t[52] = t[65] ^ x[6];
  assign t[53] = t[66] ^ x[11];
  assign t[54] = t[67] ^ x[16];
  assign t[55] = t[68] ^ x[21];
  assign t[56] = t[69] ^ x[26];
  assign t[57] = t[70] ^ x[31];
  assign t[58] = t[71] ^ x[36];
  assign t[59] = t[72] ^ x[41];
  assign t[5] = t[9] ^ t[10];
  assign t[60] = t[73] ^ x[46];
  assign t[61] = t[74] ^ x[51];
  assign t[62] = t[75] ^ x[56];
  assign t[63] = t[76] ^ x[61];
  assign t[64] = t[77] ^ x[66];
  assign t[65] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[66] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[67] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[68] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[69] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[71] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[72] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[73] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[74] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[75] = (x[52] & x[53] & x[54]) | (x[52] & x[53] & x[55]) | (x[52] & x[54] & x[55]) | (x[53] & x[54] & x[55]);
  assign t[76] = (x[57] & x[58] & x[59]) | (x[57] & x[58] & x[60]) | (x[57] & x[59] & x[60]) | (x[58] & x[59] & x[60]);
  assign t[77] = (x[62] & x[63] & x[64]) | (x[62] & x[63] & x[65]) | (x[62] & x[64] & x[65]) | (x[63] & x[64] & x[65]);
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[15] & t[16];
  assign t[9] = t[17] ^ t[18];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind185(x, y);
 input [66:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[19] ^ t[20];
  assign t[11] = t[21] ^ t[22];
  assign t[12] = t[23] ^ t[24];
  assign t[13] = t[25] ^ t[26];
  assign t[14] = t[27] & t[28];
  assign t[15] = t[29] ^ t[14];
  assign t[16] = t[53] ^ t[27];
  assign t[17] = t[30] ^ t[31];
  assign t[18] = t[32] & t[33];
  assign t[19] = t[34] ^ t[18];
  assign t[1] = ~(t[3] ^ t[52]);
  assign t[20] = t[54] ^ t[32];
  assign t[21] = t[35] ^ t[36];
  assign t[22] = t[37] & t[38];
  assign t[23] = t[39] ^ t[22];
  assign t[24] = t[55] ^ t[37];
  assign t[25] = t[56] ^ t[57];
  assign t[26] = t[27] & t[40];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[53] ^ t[27]);
  assign t[29] = t[53] & t[41];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[58] ^ t[59];
  assign t[31] = t[32] & t[42];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[54] ^ t[32]);
  assign t[34] = t[54] & t[43];
  assign t[35] = t[60] ^ t[61];
  assign t[36] = t[37] & t[44];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[55] ^ t[37]);
  assign t[39] = t[55] & t[45];
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ t[46];
  assign t[41] = t[47] ^ t[26];
  assign t[42] = t[54] ^ t[48];
  assign t[43] = t[49] ^ t[31];
  assign t[44] = t[55] ^ t[50];
  assign t[45] = t[51] ^ t[36];
  assign t[46] = t[57] ^ t[62];
  assign t[47] = t[53] ^ t[25];
  assign t[48] = t[59] ^ t[63];
  assign t[49] = t[54] ^ t[30];
  assign t[4] = ~(t[7] ^ t[8]);
  assign t[50] = t[61] ^ t[64];
  assign t[51] = t[55] ^ t[35];
  assign t[52] = t[65] ^ x[6];
  assign t[53] = t[66] ^ x[11];
  assign t[54] = t[67] ^ x[16];
  assign t[55] = t[68] ^ x[21];
  assign t[56] = t[69] ^ x[26];
  assign t[57] = t[70] ^ x[31];
  assign t[58] = t[71] ^ x[36];
  assign t[59] = t[72] ^ x[41];
  assign t[5] = ~(t[9] ^ t[10]);
  assign t[60] = t[73] ^ x[46];
  assign t[61] = t[74] ^ x[51];
  assign t[62] = t[75] ^ x[56];
  assign t[63] = t[76] ^ x[61];
  assign t[64] = t[77] ^ x[66];
  assign t[65] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[66] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[67] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[68] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[69] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[71] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[72] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[73] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[74] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[75] = (x[52] & x[53] & x[54]) | (x[52] & x[53] & x[55]) | (x[52] & x[54] & x[55]) | (x[53] & x[54] & x[55]);
  assign t[76] = (x[57] & x[58] & x[59]) | (x[57] & x[58] & x[60]) | (x[57] & x[59] & x[60]) | (x[58] & x[59] & x[60]);
  assign t[77] = (x[62] & x[63] & x[64]) | (x[62] & x[63] & x[65]) | (x[62] & x[64] & x[65]) | (x[63] & x[64] & x[65]);
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[15] ^ t[16];
  assign t[9] = t[17] ^ t[18];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind186(x, y);
 input [51:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[23] ^ t[24];
  assign t[11] = t[16] & t[17];
  assign t[12] = t[25] ^ t[26];
  assign t[13] = t[18] & t[19];
  assign t[14] = t[27] ^ t[28];
  assign t[15] = t[20] & t[21];
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[29] ^ t[16]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[30] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[22]);
  assign t[20] = ~(t[27]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[32] ^ x[6];
  assign t[23] = t[33] ^ x[11];
  assign t[24] = t[34] ^ x[16];
  assign t[25] = t[35] ^ x[21];
  assign t[26] = t[36] ^ x[26];
  assign t[27] = t[37] ^ x[31];
  assign t[28] = t[38] ^ x[36];
  assign t[29] = t[39] ^ x[41];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[46];
  assign t[31] = t[41] ^ x[51];
  assign t[32] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[33] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[34] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[35] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[36] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[37] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[38] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[39] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[3] = ~t[6];
  assign t[40] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[41] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[4] = ~(t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind187(x, y);
 input [66:0] x;
 output y;

 wire [59:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[17];
  assign t[11] = t[18] & t[19];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[22] & t[23];
  assign t[14] = t[24] ^ t[25];
  assign t[15] = t[26] & t[27];
  assign t[16] = t[35] ^ t[36];
  assign t[17] = t[18] & t[28];
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[37] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[34]);
  assign t[20] = t[38] ^ t[39];
  assign t[21] = t[22] & t[29];
  assign t[22] = ~(t[39]);
  assign t[23] = ~(t[40] ^ t[22]);
  assign t[24] = t[41] ^ t[42];
  assign t[25] = t[26] & t[30];
  assign t[26] = ~(t[42]);
  assign t[27] = ~(t[43] ^ t[26]);
  assign t[28] = t[37] ^ t[31];
  assign t[29] = t[40] ^ t[32];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[33];
  assign t[31] = t[36] ^ t[44];
  assign t[32] = t[39] ^ t[45];
  assign t[33] = t[42] ^ t[46];
  assign t[34] = t[47] ^ x[6];
  assign t[35] = t[48] ^ x[11];
  assign t[36] = t[49] ^ x[16];
  assign t[37] = t[50] ^ x[21];
  assign t[38] = t[51] ^ x[26];
  assign t[39] = t[52] ^ x[31];
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ x[36];
  assign t[41] = t[54] ^ x[41];
  assign t[42] = t[55] ^ x[46];
  assign t[43] = t[56] ^ x[51];
  assign t[44] = t[57] ^ x[56];
  assign t[45] = t[58] ^ x[61];
  assign t[46] = t[59] ^ x[66];
  assign t[47] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[48] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[49] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[4] = ~(t[7]);
  assign t[50] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[51] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[52] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[53] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[54] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[55] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[56] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[57] = (x[52] & x[53] & x[54]) | (x[52] & x[53] & x[55]) | (x[52] & x[54] & x[55]) | (x[53] & x[54] & x[55]);
  assign t[58] = (x[57] & x[58] & x[59]) | (x[57] & x[58] & x[60]) | (x[57] & x[59] & x[60]) | (x[58] & x[59] & x[60]);
  assign t[59] = (x[62] & x[63] & x[64]) | (x[62] & x[63] & x[65]) | (x[62] & x[64] & x[65]) | (x[63] & x[64] & x[65]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind188(x, y);
 input [66:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[19] & t[20];
  assign t[11] = t[21] ^ t[22];
  assign t[12] = t[23] & t[24];
  assign t[13] = t[53] & t[25];
  assign t[14] = t[26] & t[27];
  assign t[15] = t[28] ^ t[26];
  assign t[16] = t[29] ^ t[14];
  assign t[17] = t[54] & t[30];
  assign t[18] = t[31] & t[32];
  assign t[19] = t[33] ^ t[31];
  assign t[1] = ~(t[3] ^ t[52]);
  assign t[20] = t[34] ^ t[18];
  assign t[21] = t[55] & t[35];
  assign t[22] = t[36] & t[37];
  assign t[23] = t[38] ^ t[36];
  assign t[24] = t[39] ^ t[22];
  assign t[25] = t[40] ^ t[41];
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[53] ^ t[26]);
  assign t[28] = t[57] ^ t[56];
  assign t[29] = ~(t[42] ^ t[15]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[44];
  assign t[31] = ~(t[58]);
  assign t[32] = ~(t[54] ^ t[31]);
  assign t[33] = t[59] ^ t[58];
  assign t[34] = ~(t[45] ^ t[19]);
  assign t[35] = t[46] ^ t[47];
  assign t[36] = ~(t[60]);
  assign t[37] = ~(t[55] ^ t[36]);
  assign t[38] = t[61] ^ t[60];
  assign t[39] = ~(t[48] ^ t[23]);
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ t[28];
  assign t[41] = t[26] & t[42];
  assign t[42] = t[53] ^ t[49];
  assign t[43] = t[54] ^ t[33];
  assign t[44] = t[31] & t[45];
  assign t[45] = t[54] ^ t[50];
  assign t[46] = t[55] ^ t[38];
  assign t[47] = t[36] & t[48];
  assign t[48] = t[55] ^ t[51];
  assign t[49] = t[56] ^ t[62];
  assign t[4] = t[7] ^ t[8];
  assign t[50] = t[58] ^ t[63];
  assign t[51] = t[60] ^ t[64];
  assign t[52] = t[65] ^ x[6];
  assign t[53] = t[66] ^ x[11];
  assign t[54] = t[67] ^ x[16];
  assign t[55] = t[68] ^ x[21];
  assign t[56] = t[69] ^ x[26];
  assign t[57] = t[70] ^ x[31];
  assign t[58] = t[71] ^ x[36];
  assign t[59] = t[72] ^ x[41];
  assign t[5] = t[9] ^ t[10];
  assign t[60] = t[73] ^ x[46];
  assign t[61] = t[74] ^ x[51];
  assign t[62] = t[75] ^ x[56];
  assign t[63] = t[76] ^ x[61];
  assign t[64] = t[77] ^ x[66];
  assign t[65] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[66] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[67] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[68] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[69] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[71] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[72] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[73] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[74] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[75] = (x[52] & x[53] & x[54]) | (x[52] & x[53] & x[55]) | (x[52] & x[54] & x[55]) | (x[53] & x[54] & x[55]);
  assign t[76] = (x[57] & x[58] & x[59]) | (x[57] & x[58] & x[60]) | (x[57] & x[59] & x[60]) | (x[58] & x[59] & x[60]);
  assign t[77] = (x[62] & x[63] & x[64]) | (x[62] & x[63] & x[65]) | (x[62] & x[64] & x[65]) | (x[63] & x[64] & x[65]);
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[15] & t[16];
  assign t[9] = t[17] ^ t[18];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind189(x, y);
 input [66:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[20] ^ t[21];
  assign t[12] = t[22] ^ t[23];
  assign t[13] = t[24] ^ t[25];
  assign t[14] = t[26] ^ t[27];
  assign t[15] = t[28] & t[29];
  assign t[16] = t[30] ^ t[15];
  assign t[17] = t[54] ^ t[28];
  assign t[18] = t[31] ^ t[32];
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[3] ^ t[53]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[55] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[56] ^ t[38];
  assign t[26] = t[57] ^ t[58];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[58]);
  assign t[29] = ~(t[54] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[54] & t[42];
  assign t[31] = t[59] ^ t[60];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[60]);
  assign t[34] = ~(t[55] ^ t[33]);
  assign t[35] = t[55] & t[44];
  assign t[36] = t[61] ^ t[62];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[62]);
  assign t[39] = ~(t[56] ^ t[38]);
  assign t[3] = ~t[6];
  assign t[40] = t[56] & t[46];
  assign t[41] = t[54] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[55] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[56] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[58] ^ t[63];
  assign t[48] = t[54] ^ t[26];
  assign t[49] = t[60] ^ t[64];
  assign t[4] = ~(t[7]);
  assign t[50] = t[55] ^ t[31];
  assign t[51] = t[62] ^ t[65];
  assign t[52] = t[56] ^ t[36];
  assign t[53] = t[66] ^ x[6];
  assign t[54] = t[67] ^ x[11];
  assign t[55] = t[68] ^ x[16];
  assign t[56] = t[69] ^ x[21];
  assign t[57] = t[70] ^ x[26];
  assign t[58] = t[71] ^ x[31];
  assign t[59] = t[72] ^ x[36];
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = t[73] ^ x[41];
  assign t[61] = t[74] ^ x[46];
  assign t[62] = t[75] ^ x[51];
  assign t[63] = t[76] ^ x[56];
  assign t[64] = t[77] ^ x[61];
  assign t[65] = t[78] ^ x[66];
  assign t[66] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[67] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[68] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[69] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[71] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[72] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[73] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[74] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[75] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[76] = (x[52] & x[53] & x[54]) | (x[52] & x[53] & x[55]) | (x[52] & x[54] & x[55]) | (x[53] & x[54] & x[55]);
  assign t[77] = (x[57] & x[58] & x[59]) | (x[57] & x[58] & x[60]) | (x[57] & x[59] & x[60]) | (x[58] & x[59] & x[60]);
  assign t[78] = (x[62] & x[63] & x[64]) | (x[62] & x[63] & x[65]) | (x[62] & x[64] & x[65]) | (x[63] & x[64] & x[65]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[8] = t[14] ^ t[15];
  assign t[9] = t[16] ^ t[17];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind190(x, y);
 input [51:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[23] ^ t[24];
  assign t[11] = t[16] & t[17];
  assign t[12] = t[25] ^ t[26];
  assign t[13] = t[18] & t[19];
  assign t[14] = t[27] ^ t[28];
  assign t[15] = t[20] & t[21];
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[29] ^ t[16]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[30] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[22]);
  assign t[20] = ~(t[27]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[32] ^ x[6];
  assign t[23] = t[33] ^ x[11];
  assign t[24] = t[34] ^ x[16];
  assign t[25] = t[35] ^ x[21];
  assign t[26] = t[36] ^ x[26];
  assign t[27] = t[37] ^ x[31];
  assign t[28] = t[38] ^ x[36];
  assign t[29] = t[39] ^ x[41];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[46];
  assign t[31] = t[41] ^ x[51];
  assign t[32] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[33] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[34] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[35] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[36] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[37] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[38] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[39] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[3] = ~t[6];
  assign t[40] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[41] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[4] = ~(t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind191(x, y);
 input [66:0] x;
 output y;

 wire [59:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[17];
  assign t[11] = t[18] & t[19];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[22] & t[23];
  assign t[14] = t[24] ^ t[25];
  assign t[15] = t[26] & t[27];
  assign t[16] = t[35] ^ t[36];
  assign t[17] = t[18] & t[28];
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[37] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[34]);
  assign t[20] = t[38] ^ t[39];
  assign t[21] = t[22] & t[29];
  assign t[22] = ~(t[39]);
  assign t[23] = ~(t[40] ^ t[22]);
  assign t[24] = t[41] ^ t[42];
  assign t[25] = t[26] & t[30];
  assign t[26] = ~(t[42]);
  assign t[27] = ~(t[43] ^ t[26]);
  assign t[28] = t[37] ^ t[31];
  assign t[29] = t[40] ^ t[32];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[33];
  assign t[31] = t[36] ^ t[44];
  assign t[32] = t[39] ^ t[45];
  assign t[33] = t[42] ^ t[46];
  assign t[34] = t[47] ^ x[6];
  assign t[35] = t[48] ^ x[11];
  assign t[36] = t[49] ^ x[16];
  assign t[37] = t[50] ^ x[21];
  assign t[38] = t[51] ^ x[26];
  assign t[39] = t[52] ^ x[31];
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ x[36];
  assign t[41] = t[54] ^ x[41];
  assign t[42] = t[55] ^ x[46];
  assign t[43] = t[56] ^ x[51];
  assign t[44] = t[57] ^ x[56];
  assign t[45] = t[58] ^ x[61];
  assign t[46] = t[59] ^ x[66];
  assign t[47] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[48] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[49] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[4] = ~(t[7]);
  assign t[50] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[51] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[52] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[53] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[54] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[55] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[56] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[57] = (x[52] & x[53] & x[54]) | (x[52] & x[53] & x[55]) | (x[52] & x[54] & x[55]) | (x[53] & x[54] & x[55]);
  assign t[58] = (x[57] & x[58] & x[59]) | (x[57] & x[58] & x[60]) | (x[57] & x[59] & x[60]) | (x[58] & x[59] & x[60]);
  assign t[59] = (x[62] & x[63] & x[64]) | (x[62] & x[63] & x[65]) | (x[62] & x[64] & x[65]) | (x[63] & x[64] & x[65]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind192(x, y);
 input [66:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[19] & t[20];
  assign t[11] = t[21] ^ t[22];
  assign t[12] = t[23] & t[24];
  assign t[13] = t[53] & t[25];
  assign t[14] = t[26] & t[27];
  assign t[15] = t[28] ^ t[26];
  assign t[16] = t[29] ^ t[14];
  assign t[17] = t[54] & t[30];
  assign t[18] = t[31] & t[32];
  assign t[19] = t[33] ^ t[31];
  assign t[1] = ~(t[3] ^ t[52]);
  assign t[20] = t[34] ^ t[18];
  assign t[21] = t[55] & t[35];
  assign t[22] = t[36] & t[37];
  assign t[23] = t[38] ^ t[36];
  assign t[24] = t[39] ^ t[22];
  assign t[25] = t[40] ^ t[41];
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[53] ^ t[26]);
  assign t[28] = t[57] ^ t[56];
  assign t[29] = ~(t[42] ^ t[15]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[44];
  assign t[31] = ~(t[58]);
  assign t[32] = ~(t[54] ^ t[31]);
  assign t[33] = t[59] ^ t[58];
  assign t[34] = ~(t[45] ^ t[19]);
  assign t[35] = t[46] ^ t[47];
  assign t[36] = ~(t[60]);
  assign t[37] = ~(t[55] ^ t[36]);
  assign t[38] = t[61] ^ t[60];
  assign t[39] = ~(t[48] ^ t[23]);
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ t[28];
  assign t[41] = t[26] & t[42];
  assign t[42] = t[53] ^ t[49];
  assign t[43] = t[54] ^ t[33];
  assign t[44] = t[31] & t[45];
  assign t[45] = t[54] ^ t[50];
  assign t[46] = t[55] ^ t[38];
  assign t[47] = t[36] & t[48];
  assign t[48] = t[55] ^ t[51];
  assign t[49] = t[56] ^ t[62];
  assign t[4] = t[7] ^ t[8];
  assign t[50] = t[58] ^ t[63];
  assign t[51] = t[60] ^ t[64];
  assign t[52] = t[65] ^ x[6];
  assign t[53] = t[66] ^ x[11];
  assign t[54] = t[67] ^ x[16];
  assign t[55] = t[68] ^ x[21];
  assign t[56] = t[69] ^ x[26];
  assign t[57] = t[70] ^ x[31];
  assign t[58] = t[71] ^ x[36];
  assign t[59] = t[72] ^ x[41];
  assign t[5] = t[9] ^ t[10];
  assign t[60] = t[73] ^ x[46];
  assign t[61] = t[74] ^ x[51];
  assign t[62] = t[75] ^ x[56];
  assign t[63] = t[76] ^ x[61];
  assign t[64] = t[77] ^ x[66];
  assign t[65] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[66] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[67] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[68] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[69] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[71] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[72] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[73] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[74] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[75] = (x[52] & x[53] & x[54]) | (x[52] & x[53] & x[55]) | (x[52] & x[54] & x[55]) | (x[53] & x[54] & x[55]);
  assign t[76] = (x[57] & x[58] & x[59]) | (x[57] & x[58] & x[60]) | (x[57] & x[59] & x[60]) | (x[58] & x[59] & x[60]);
  assign t[77] = (x[62] & x[63] & x[64]) | (x[62] & x[63] & x[65]) | (x[62] & x[64] & x[65]) | (x[63] & x[64] & x[65]);
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[15] & t[16];
  assign t[9] = t[17] ^ t[18];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind193(x, y);
 input [66:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[19] ^ t[20];
  assign t[11] = t[21] ^ t[22];
  assign t[12] = t[23] ^ t[24];
  assign t[13] = t[25] ^ t[26];
  assign t[14] = t[27] & t[28];
  assign t[15] = t[29] ^ t[14];
  assign t[16] = t[53] ^ t[27];
  assign t[17] = t[30] ^ t[31];
  assign t[18] = t[32] & t[33];
  assign t[19] = t[34] ^ t[18];
  assign t[1] = ~(t[3] ^ t[52]);
  assign t[20] = t[54] ^ t[32];
  assign t[21] = t[35] ^ t[36];
  assign t[22] = t[37] & t[38];
  assign t[23] = t[39] ^ t[22];
  assign t[24] = t[55] ^ t[37];
  assign t[25] = t[56] ^ t[57];
  assign t[26] = t[27] & t[40];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[53] ^ t[27]);
  assign t[29] = t[53] & t[41];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[58] ^ t[59];
  assign t[31] = t[32] & t[42];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[54] ^ t[32]);
  assign t[34] = t[54] & t[43];
  assign t[35] = t[60] ^ t[61];
  assign t[36] = t[37] & t[44];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[55] ^ t[37]);
  assign t[39] = t[55] & t[45];
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ t[46];
  assign t[41] = t[47] ^ t[26];
  assign t[42] = t[54] ^ t[48];
  assign t[43] = t[49] ^ t[31];
  assign t[44] = t[55] ^ t[50];
  assign t[45] = t[51] ^ t[36];
  assign t[46] = t[57] ^ t[62];
  assign t[47] = t[53] ^ t[25];
  assign t[48] = t[59] ^ t[63];
  assign t[49] = t[54] ^ t[30];
  assign t[4] = ~(t[7] ^ t[8]);
  assign t[50] = t[61] ^ t[64];
  assign t[51] = t[55] ^ t[35];
  assign t[52] = t[65] ^ x[6];
  assign t[53] = t[66] ^ x[11];
  assign t[54] = t[67] ^ x[16];
  assign t[55] = t[68] ^ x[21];
  assign t[56] = t[69] ^ x[26];
  assign t[57] = t[70] ^ x[31];
  assign t[58] = t[71] ^ x[36];
  assign t[59] = t[72] ^ x[41];
  assign t[5] = ~(t[9] ^ t[10]);
  assign t[60] = t[73] ^ x[46];
  assign t[61] = t[74] ^ x[51];
  assign t[62] = t[75] ^ x[56];
  assign t[63] = t[76] ^ x[61];
  assign t[64] = t[77] ^ x[66];
  assign t[65] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[66] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[67] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[68] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[69] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[71] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[72] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[73] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[74] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[75] = (x[52] & x[53] & x[54]) | (x[52] & x[53] & x[55]) | (x[52] & x[54] & x[55]) | (x[53] & x[54] & x[55]);
  assign t[76] = (x[57] & x[58] & x[59]) | (x[57] & x[58] & x[60]) | (x[57] & x[59] & x[60]) | (x[58] & x[59] & x[60]);
  assign t[77] = (x[62] & x[63] & x[64]) | (x[62] & x[63] & x[65]) | (x[62] & x[64] & x[65]) | (x[63] & x[64] & x[65]);
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[15] ^ t[16];
  assign t[9] = t[17] ^ t[18];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind194(x, y);
 input [51:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[23] ^ t[24];
  assign t[11] = t[16] & t[17];
  assign t[12] = t[25] ^ t[26];
  assign t[13] = t[18] & t[19];
  assign t[14] = t[27] ^ t[28];
  assign t[15] = t[20] & t[21];
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[29] ^ t[16]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[30] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[22]);
  assign t[20] = ~(t[27]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[32] ^ x[6];
  assign t[23] = t[33] ^ x[11];
  assign t[24] = t[34] ^ x[16];
  assign t[25] = t[35] ^ x[21];
  assign t[26] = t[36] ^ x[26];
  assign t[27] = t[37] ^ x[31];
  assign t[28] = t[38] ^ x[36];
  assign t[29] = t[39] ^ x[41];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[46];
  assign t[31] = t[41] ^ x[51];
  assign t[32] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[33] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[34] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[35] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[36] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[37] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[38] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[39] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[3] = ~t[6];
  assign t[40] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[41] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[4] = ~(t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind195(x, y);
 input [66:0] x;
 output y;

 wire [59:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[17];
  assign t[11] = t[18] & t[19];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[22] & t[23];
  assign t[14] = t[24] ^ t[25];
  assign t[15] = t[26] & t[27];
  assign t[16] = t[35] ^ t[36];
  assign t[17] = t[18] & t[28];
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[37] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[34]);
  assign t[20] = t[38] ^ t[39];
  assign t[21] = t[22] & t[29];
  assign t[22] = ~(t[39]);
  assign t[23] = ~(t[40] ^ t[22]);
  assign t[24] = t[41] ^ t[42];
  assign t[25] = t[26] & t[30];
  assign t[26] = ~(t[42]);
  assign t[27] = ~(t[43] ^ t[26]);
  assign t[28] = t[37] ^ t[31];
  assign t[29] = t[40] ^ t[32];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[33];
  assign t[31] = t[36] ^ t[44];
  assign t[32] = t[39] ^ t[45];
  assign t[33] = t[42] ^ t[46];
  assign t[34] = t[47] ^ x[6];
  assign t[35] = t[48] ^ x[11];
  assign t[36] = t[49] ^ x[16];
  assign t[37] = t[50] ^ x[21];
  assign t[38] = t[51] ^ x[26];
  assign t[39] = t[52] ^ x[31];
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ x[36];
  assign t[41] = t[54] ^ x[41];
  assign t[42] = t[55] ^ x[46];
  assign t[43] = t[56] ^ x[51];
  assign t[44] = t[57] ^ x[56];
  assign t[45] = t[58] ^ x[61];
  assign t[46] = t[59] ^ x[66];
  assign t[47] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[48] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[49] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[4] = ~(t[7]);
  assign t[50] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[51] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[52] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[53] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[54] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[55] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[56] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[57] = (x[52] & x[53] & x[54]) | (x[52] & x[53] & x[55]) | (x[52] & x[54] & x[55]) | (x[53] & x[54] & x[55]);
  assign t[58] = (x[57] & x[58] & x[59]) | (x[57] & x[58] & x[60]) | (x[57] & x[59] & x[60]) | (x[58] & x[59] & x[60]);
  assign t[59] = (x[62] & x[63] & x[64]) | (x[62] & x[63] & x[65]) | (x[62] & x[64] & x[65]) | (x[63] & x[64] & x[65]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind196(x, y);
 input [71:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] & t[19];
  assign t[11] = ~t[20];
  assign t[12] = t[56] & t[21];
  assign t[13] = t[22] & t[23];
  assign t[14] = t[24] ^ t[22];
  assign t[15] = t[25] ^ t[13];
  assign t[16] = t[57] & t[26];
  assign t[17] = t[27] & t[28];
  assign t[18] = t[29] ^ t[27];
  assign t[19] = t[30] ^ t[17];
  assign t[1] = ~(t[3] ^ t[54]);
  assign t[20] = t[31] ^ t[32];
  assign t[21] = t[33] ^ t[34];
  assign t[22] = ~(t[58]);
  assign t[23] = ~(t[56] ^ t[22]);
  assign t[24] = t[59] ^ t[58];
  assign t[25] = ~(t[35] ^ t[14]);
  assign t[26] = t[36] ^ t[37];
  assign t[27] = ~(t[60]);
  assign t[28] = ~(t[57] ^ t[27]);
  assign t[29] = t[61] ^ t[60];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[38] ^ t[18]);
  assign t[31] = t[39] ^ t[40];
  assign t[32] = t[41] & t[42];
  assign t[33] = t[56] ^ t[24];
  assign t[34] = t[22] & t[35];
  assign t[35] = t[56] ^ t[43];
  assign t[36] = t[57] ^ t[29];
  assign t[37] = t[27] & t[38];
  assign t[38] = t[57] ^ t[44];
  assign t[39] = t[62] & t[45];
  assign t[3] = ~t[6];
  assign t[40] = t[46] & t[47];
  assign t[41] = t[48] ^ t[46];
  assign t[42] = t[49] ^ t[40];
  assign t[43] = t[58] ^ t[63];
  assign t[44] = t[60] ^ t[64];
  assign t[45] = t[50] ^ t[51];
  assign t[46] = ~(t[65]);
  assign t[47] = ~(t[62] ^ t[46]);
  assign t[48] = t[66] ^ t[65];
  assign t[49] = ~(t[52] ^ t[41]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = t[62] ^ t[48];
  assign t[51] = t[46] & t[52];
  assign t[52] = t[62] ^ t[53];
  assign t[53] = t[65] ^ t[67];
  assign t[54] = t[68] ^ x[6];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = t[71] ^ x[21];
  assign t[58] = t[72] ^ x[26];
  assign t[59] = t[73] ^ x[31];
  assign t[5] = t[9] ^ t[10];
  assign t[60] = t[74] ^ x[36];
  assign t[61] = t[75] ^ x[41];
  assign t[62] = t[76] ^ x[46];
  assign t[63] = t[77] ^ x[51];
  assign t[64] = t[78] ^ x[56];
  assign t[65] = t[79] ^ x[61];
  assign t[66] = t[80] ^ x[66];
  assign t[67] = t[81] ^ x[71];
  assign t[68] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[69] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[6] = ~(t[11] ^ t[55]);
  assign t[70] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[71] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[72] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[73] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[74] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[75] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[76] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[77] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[78] = (x[52] & x[53] & x[54]) | (x[52] & x[53] & x[55]) | (x[52] & x[54] & x[55]) | (x[53] & x[54] & x[55]);
  assign t[79] = (x[57] & x[58] & x[59]) | (x[57] & x[58] & x[60]) | (x[57] & x[59] & x[60]) | (x[58] & x[59] & x[60]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[62] & x[63] & x[64]) | (x[62] & x[63] & x[65]) | (x[62] & x[64] & x[65]) | (x[63] & x[64] & x[65]);
  assign t[81] = (x[67] & x[68] & x[69]) | (x[67] & x[68] & x[70]) | (x[67] & x[69] & x[70]) | (x[68] & x[69] & x[70]);
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[17];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind197(x, y);
 input [71:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = ~t[20];
  assign t[12] = t[21] ^ t[22];
  assign t[13] = t[23] & t[24];
  assign t[14] = t[25] ^ t[13];
  assign t[15] = t[56] ^ t[23];
  assign t[16] = t[26] ^ t[27];
  assign t[17] = t[28] & t[29];
  assign t[18] = t[30] ^ t[17];
  assign t[19] = t[57] ^ t[28];
  assign t[1] = ~(t[3] ^ t[54]);
  assign t[20] = ~(t[31] ^ t[32]);
  assign t[21] = t[58] ^ t[59];
  assign t[22] = t[23] & t[33];
  assign t[23] = ~(t[59]);
  assign t[24] = ~(t[56] ^ t[23]);
  assign t[25] = t[56] & t[34];
  assign t[26] = t[60] ^ t[61];
  assign t[27] = t[28] & t[35];
  assign t[28] = ~(t[61]);
  assign t[29] = ~(t[57] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[57] & t[36];
  assign t[31] = t[37] ^ t[38];
  assign t[32] = t[39] ^ t[40];
  assign t[33] = t[56] ^ t[41];
  assign t[34] = t[42] ^ t[22];
  assign t[35] = t[57] ^ t[43];
  assign t[36] = t[44] ^ t[27];
  assign t[37] = t[45] ^ t[46];
  assign t[38] = t[47] & t[48];
  assign t[39] = t[49] ^ t[38];
  assign t[3] = ~t[6];
  assign t[40] = t[62] ^ t[47];
  assign t[41] = t[59] ^ t[63];
  assign t[42] = t[56] ^ t[21];
  assign t[43] = t[61] ^ t[64];
  assign t[44] = t[57] ^ t[26];
  assign t[45] = t[65] ^ t[66];
  assign t[46] = t[47] & t[50];
  assign t[47] = ~(t[66]);
  assign t[48] = ~(t[62] ^ t[47]);
  assign t[49] = t[62] & t[51];
  assign t[4] = ~(t[7] ^ t[8]);
  assign t[50] = t[62] ^ t[52];
  assign t[51] = t[53] ^ t[46];
  assign t[52] = t[66] ^ t[67];
  assign t[53] = t[62] ^ t[45];
  assign t[54] = t[68] ^ x[6];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = t[71] ^ x[21];
  assign t[58] = t[72] ^ x[26];
  assign t[59] = t[73] ^ x[31];
  assign t[5] = ~(t[9] ^ t[10]);
  assign t[60] = t[74] ^ x[36];
  assign t[61] = t[75] ^ x[41];
  assign t[62] = t[76] ^ x[46];
  assign t[63] = t[77] ^ x[51];
  assign t[64] = t[78] ^ x[56];
  assign t[65] = t[79] ^ x[61];
  assign t[66] = t[80] ^ x[66];
  assign t[67] = t[81] ^ x[71];
  assign t[68] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[69] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[6] = ~(t[11] ^ t[55]);
  assign t[70] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[71] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[72] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[73] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[74] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[75] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[76] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[77] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[78] = (x[52] & x[53] & x[54]) | (x[52] & x[53] & x[55]) | (x[52] & x[54] & x[55]) | (x[53] & x[54] & x[55]);
  assign t[79] = (x[57] & x[58] & x[59]) | (x[57] & x[58] & x[60]) | (x[57] & x[59] & x[60]) | (x[58] & x[59] & x[60]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[62] & x[63] & x[64]) | (x[62] & x[63] & x[65]) | (x[62] & x[64] & x[65]) | (x[63] & x[64] & x[65]);
  assign t[81] = (x[67] & x[68] & x[69]) | (x[67] & x[68] & x[70]) | (x[67] & x[69] & x[70]) | (x[68] & x[69] & x[70]);
  assign t[8] = t[14] ^ t[15];
  assign t[9] = t[16] ^ t[17];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind198(x, y);
 input [56:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[26] ^ t[27];
  assign t[11] = t[15] & t[16];
  assign t[12] = t[28] ^ t[29];
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[19]);
  assign t[15] = ~(t[26]);
  assign t[16] = ~(t[30] ^ t[15]);
  assign t[17] = ~(t[28]);
  assign t[18] = ~(t[31] ^ t[17]);
  assign t[19] = t[20] ^ t[21];
  assign t[1] = ~(t[3] ^ t[24]);
  assign t[20] = t[32] ^ t[33];
  assign t[21] = t[22] & t[23];
  assign t[22] = ~(t[32]);
  assign t[23] = ~(t[34] ^ t[22]);
  assign t[24] = t[35] ^ x[6];
  assign t[25] = t[36] ^ x[11];
  assign t[26] = t[37] ^ x[16];
  assign t[27] = t[38] ^ x[21];
  assign t[28] = t[39] ^ x[26];
  assign t[29] = t[40] ^ x[31];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[41] ^ x[36];
  assign t[31] = t[42] ^ x[41];
  assign t[32] = t[43] ^ x[46];
  assign t[33] = t[44] ^ x[51];
  assign t[34] = t[45] ^ x[56];
  assign t[35] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[36] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[37] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[38] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[39] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[3] = ~t[6];
  assign t[40] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[41] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[42] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[43] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[44] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[45] = (x[52] & x[53] & x[54]) | (x[52] & x[53] & x[55]) | (x[52] & x[54] & x[55]) | (x[53] & x[54] & x[55]);
  assign t[4] = ~(t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] ^ t[25]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = ~t[14];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind199(x, y);
 input [71:0] x;
 output y;

 wire [63:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[15] ^ t[16];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = t[21] & t[22];
  assign t[14] = ~(t[23]);
  assign t[15] = t[38] ^ t[39];
  assign t[16] = t[17] & t[24];
  assign t[17] = ~(t[39]);
  assign t[18] = ~(t[40] ^ t[17]);
  assign t[19] = t[41] ^ t[42];
  assign t[1] = ~(t[3] ^ t[36]);
  assign t[20] = t[21] & t[25];
  assign t[21] = ~(t[42]);
  assign t[22] = ~(t[43] ^ t[21]);
  assign t[23] = t[26] ^ t[27];
  assign t[24] = t[40] ^ t[28];
  assign t[25] = t[43] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[39] ^ t[44];
  assign t[29] = t[42] ^ t[45];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[46] ^ t[47];
  assign t[31] = t[32] & t[34];
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[48] ^ t[32]);
  assign t[34] = t[48] ^ t[35];
  assign t[35] = t[47] ^ t[49];
  assign t[36] = t[50] ^ x[6];
  assign t[37] = t[51] ^ x[11];
  assign t[38] = t[52] ^ x[16];
  assign t[39] = t[53] ^ x[21];
  assign t[3] = ~t[6];
  assign t[40] = t[54] ^ x[26];
  assign t[41] = t[55] ^ x[31];
  assign t[42] = t[56] ^ x[36];
  assign t[43] = t[57] ^ x[41];
  assign t[44] = t[58] ^ x[46];
  assign t[45] = t[59] ^ x[51];
  assign t[46] = t[60] ^ x[56];
  assign t[47] = t[61] ^ x[61];
  assign t[48] = t[62] ^ x[66];
  assign t[49] = t[63] ^ x[71];
  assign t[4] = ~(t[7]);
  assign t[50] = (x[2] & x[3] & x[4]) | (x[2] & x[3] & x[5]) | (x[2] & x[4] & x[5]) | (x[3] & x[4] & x[5]);
  assign t[51] = (x[7] & x[8] & x[9]) | (x[7] & x[8] & x[10]) | (x[7] & x[9] & x[10]) | (x[8] & x[9] & x[10]);
  assign t[52] = (x[12] & x[13] & x[14]) | (x[12] & x[13] & x[15]) | (x[12] & x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[53] = (x[17] & x[18] & x[19]) | (x[17] & x[18] & x[20]) | (x[17] & x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[54] = (x[22] & x[23] & x[24]) | (x[22] & x[23] & x[25]) | (x[22] & x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[55] = (x[27] & x[28] & x[29]) | (x[27] & x[28] & x[30]) | (x[27] & x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[56] = (x[32] & x[33] & x[34]) | (x[32] & x[33] & x[35]) | (x[32] & x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[57] = (x[37] & x[38] & x[39]) | (x[37] & x[38] & x[40]) | (x[37] & x[39] & x[40]) | (x[38] & x[39] & x[40]);
  assign t[58] = (x[42] & x[43] & x[44]) | (x[42] & x[43] & x[45]) | (x[42] & x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[59] = (x[47] & x[48] & x[49]) | (x[47] & x[48] & x[50]) | (x[47] & x[49] & x[50]) | (x[48] & x[49] & x[50]);
  assign t[5] = ~(t[8]);
  assign t[60] = (x[52] & x[53] & x[54]) | (x[52] & x[53] & x[55]) | (x[52] & x[54] & x[55]) | (x[53] & x[54] & x[55]);
  assign t[61] = (x[57] & x[58] & x[59]) | (x[57] & x[58] & x[60]) | (x[57] & x[59] & x[60]) | (x[58] & x[59] & x[60]);
  assign t[62] = (x[62] & x[63] & x[64]) | (x[62] & x[63] & x[65]) | (x[62] & x[64] & x[65]) | (x[63] & x[64] & x[65]);
  assign t[63] = (x[67] & x[68] & x[69]) | (x[67] & x[68] & x[70]) | (x[67] & x[69] & x[70]) | (x[68] & x[69] & x[70]);
  assign t[6] = ~(t[9] ^ t[37]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = ~t[14];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1_ind(x, y);
 input [803:0] x;
 output [199:0] y;

  R1ind0 R1ind0_inst(.x({x[4], x[3], x[2], x[1], x[0]}), .y(y[0]));
  R1ind1 R1ind1_inst(.x({x[9], x[8], x[7], x[6], x[5]}), .y(y[1]));
  R1ind2 R1ind2_inst(.x({x[14], x[13], x[12], x[11], x[10]}), .y(y[2]));
  R1ind3 R1ind3_inst(.x({x[19], x[18], x[17], x[16], x[15]}), .y(y[3]));
  R1ind4 R1ind4_inst(.x({x[24], x[23], x[22], x[21], x[20]}), .y(y[4]));
  R1ind5 R1ind5_inst(.x({x[29], x[28], x[27], x[26], x[25]}), .y(y[5]));
  R1ind6 R1ind6_inst(.x({x[34], x[33], x[32], x[31], x[30]}), .y(y[6]));
  R1ind7 R1ind7_inst(.x({x[39], x[38], x[37], x[36], x[35]}), .y(y[7]));
  R1ind8 R1ind8_inst(.x({x[44], x[43], x[42], x[41], x[40]}), .y(y[8]));
  R1ind9 R1ind9_inst(.x({x[49], x[48], x[47], x[46], x[45]}), .y(y[9]));
  R1ind10 R1ind10_inst(.x({x[54], x[53], x[52], x[51], x[50]}), .y(y[10]));
  R1ind11 R1ind11_inst(.x({x[59], x[58], x[57], x[56], x[55]}), .y(y[11]));
  R1ind12 R1ind12_inst(.x({x[64], x[63], x[62], x[61], x[60]}), .y(y[12]));
  R1ind13 R1ind13_inst(.x({x[69], x[68], x[67], x[66], x[65]}), .y(y[13]));
  R1ind14 R1ind14_inst(.x({x[74], x[73], x[72], x[71], x[70]}), .y(y[14]));
  R1ind15 R1ind15_inst(.x({x[79], x[78], x[77], x[76], x[75]}), .y(y[15]));
  R1ind16 R1ind16_inst(.x({x[84], x[83], x[82], x[81], x[80]}), .y(y[16]));
  R1ind17 R1ind17_inst(.x({x[89], x[88], x[87], x[86], x[85]}), .y(y[17]));
  R1ind18 R1ind18_inst(.x({x[94], x[93], x[92], x[91], x[90]}), .y(y[18]));
  R1ind19 R1ind19_inst(.x({x[99], x[98], x[97], x[96], x[95]}), .y(y[19]));
  R1ind20 R1ind20_inst(.x({x[104], x[103], x[102], x[101], x[100]}), .y(y[20]));
  R1ind21 R1ind21_inst(.x({x[109], x[108], x[107], x[106], x[105]}), .y(y[21]));
  R1ind22 R1ind22_inst(.x({x[114], x[113], x[112], x[111], x[110]}), .y(y[22]));
  R1ind23 R1ind23_inst(.x({x[119], x[118], x[117], x[116], x[115]}), .y(y[23]));
  R1ind24 R1ind24_inst(.x({x[124], x[123], x[122], x[121], x[120]}), .y(y[24]));
  R1ind25 R1ind25_inst(.x({x[129], x[128], x[127], x[126], x[125]}), .y(y[25]));
  R1ind26 R1ind26_inst(.x({x[134], x[133], x[132], x[131], x[130]}), .y(y[26]));
  R1ind27 R1ind27_inst(.x({x[139], x[138], x[137], x[136], x[135]}), .y(y[27]));
  R1ind28 R1ind28_inst(.x({x[144], x[143], x[142], x[141], x[140]}), .y(y[28]));
  R1ind29 R1ind29_inst(.x({x[149], x[148], x[147], x[146], x[145]}), .y(y[29]));
  R1ind30 R1ind30_inst(.x({x[154], x[153], x[152], x[151], x[150]}), .y(y[30]));
  R1ind31 R1ind31_inst(.x({x[159], x[158], x[157], x[156], x[155]}), .y(y[31]));
  R1ind32 R1ind32_inst(.x({x[164], x[163], x[162], x[161], x[160]}), .y(y[32]));
  R1ind33 R1ind33_inst(.x({x[169], x[168], x[167], x[166], x[165]}), .y(y[33]));
  R1ind34 R1ind34_inst(.x({x[174], x[173], x[172], x[171], x[170]}), .y(y[34]));
  R1ind35 R1ind35_inst(.x({x[179], x[178], x[177], x[176], x[175]}), .y(y[35]));
  R1ind36 R1ind36_inst(.x({x[184], x[183], x[182], x[181], x[180]}), .y(y[36]));
  R1ind37 R1ind37_inst(.x({x[189], x[188], x[187], x[186], x[185]}), .y(y[37]));
  R1ind38 R1ind38_inst(.x({x[194], x[193], x[192], x[191], x[190]}), .y(y[38]));
  R1ind39 R1ind39_inst(.x({x[199], x[198], x[197], x[196], x[195]}), .y(y[39]));
  R1ind40 R1ind40_inst(.x({x[204], x[203], x[202], x[201], x[200]}), .y(y[40]));
  R1ind41 R1ind41_inst(.x({x[209], x[208], x[207], x[206], x[205]}), .y(y[41]));
  R1ind42 R1ind42_inst(.x({x[214], x[213], x[212], x[211], x[210]}), .y(y[42]));
  R1ind43 R1ind43_inst(.x({x[219], x[218], x[217], x[216], x[215]}), .y(y[43]));
  R1ind44 R1ind44_inst(.x({x[224], x[223], x[222], x[221], x[220]}), .y(y[44]));
  R1ind45 R1ind45_inst(.x({x[229], x[228], x[227], x[226], x[225]}), .y(y[45]));
  R1ind46 R1ind46_inst(.x({x[234], x[233], x[232], x[231], x[230]}), .y(y[46]));
  R1ind47 R1ind47_inst(.x({x[239], x[238], x[237], x[236], x[235]}), .y(y[47]));
  R1ind48 R1ind48_inst(.x({x[244], x[243], x[242], x[241], x[240]}), .y(y[48]));
  R1ind49 R1ind49_inst(.x({x[249], x[248], x[247], x[246], x[245]}), .y(y[49]));
  R1ind50 R1ind50_inst(.x({x[254], x[253], x[252], x[251], x[250]}), .y(y[50]));
  R1ind51 R1ind51_inst(.x({x[259], x[258], x[257], x[256], x[255]}), .y(y[51]));
  R1ind52 R1ind52_inst(.x({x[264], x[263], x[262], x[261], x[260]}), .y(y[52]));
  R1ind53 R1ind53_inst(.x({x[269], x[268], x[267], x[266], x[265]}), .y(y[53]));
  R1ind54 R1ind54_inst(.x({x[274], x[273], x[272], x[271], x[270]}), .y(y[54]));
  R1ind55 R1ind55_inst(.x({x[279], x[278], x[277], x[276], x[275]}), .y(y[55]));
  R1ind56 R1ind56_inst(.x({x[284], x[283], x[282], x[281], x[280]}), .y(y[56]));
  R1ind57 R1ind57_inst(.x({x[289], x[288], x[287], x[286], x[285]}), .y(y[57]));
  R1ind58 R1ind58_inst(.x({x[294], x[293], x[292], x[291], x[290]}), .y(y[58]));
  R1ind59 R1ind59_inst(.x({x[299], x[298], x[297], x[296], x[295]}), .y(y[59]));
  R1ind60 R1ind60_inst(.x({x[304], x[303], x[302], x[301], x[300]}), .y(y[60]));
  R1ind61 R1ind61_inst(.x({x[309], x[308], x[307], x[306], x[305]}), .y(y[61]));
  R1ind62 R1ind62_inst(.x({x[314], x[313], x[312], x[311], x[310]}), .y(y[62]));
  R1ind63 R1ind63_inst(.x({x[319], x[318], x[317], x[316], x[315]}), .y(y[63]));
  R1ind64 R1ind64_inst(.x({x[324], x[323], x[322], x[321], x[320]}), .y(y[64]));
  R1ind65 R1ind65_inst(.x({x[354], x[353], x[352], x[351], x[350], x[349], x[348], x[347], x[346], x[345], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[337], x[336], x[335], x[334], x[333], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[325]}), .y(y[65]));
  R1ind66 R1ind66_inst(.x({x[349], x[348], x[347], x[346], x[345], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[337], x[336], x[335], x[354], x[353], x[352], x[351], x[350], x[334], x[333], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[325], x[355]}), .y(y[66]));
  R1ind67 R1ind67_inst(.x({x[354], x[353], x[352], x[351], x[350], x[355]}), .y(y[67]));
  R1ind68 R1ind68_inst(.x({x[349], x[348], x[347], x[346], x[345], x[344], x[343], x[342], x[341], x[340], x[354], x[353], x[352], x[351], x[350], x[329], x[328], x[327], x[326], x[325], x[334], x[333], x[332], x[331], x[330], x[339], x[338], x[337], x[336], x[335], x[355]}), .y(y[68]));
  R1ind69 R1ind69_inst(.x({x[344], x[343], x[342], x[341], x[340], x[355]}), .y(y[69]));
  R1ind70 R1ind70_inst(.x({x[349], x[348], x[347], x[346], x[345], x[355]}), .y(y[70]));
  R1ind71 R1ind71_inst(.x({x[339], x[338], x[337], x[336], x[335], x[354], x[353], x[352], x[351], x[350], x[344], x[343], x[342], x[341], x[340], x[334], x[333], x[332], x[331], x[330], x[349], x[348], x[347], x[346], x[345], x[329], x[328], x[327], x[326], x[325], x[355]}), .y(y[71]));
  R1ind72 R1ind72_inst(.x({x[361], x[360], x[359], x[358], x[357], x[356], x[355]}), .y(y[72]));
  R1ind73 R1ind73_inst(.x({x[367], x[366], x[365], x[364], x[363], x[362], x[355]}), .y(y[73]));
  R1ind74 R1ind74_inst(.x({x[373], x[372], x[371], x[370], x[369], x[368], x[355]}), .y(y[74]));
  R1ind75 R1ind75_inst(.x({x[379], x[378], x[377], x[376], x[375], x[374], x[355]}), .y(y[75]));
  R1ind76 R1ind76_inst(.x({x[385], x[384], x[383], x[382], x[381], x[380], x[355]}), .y(y[76]));
  R1ind77 R1ind77_inst(.x({x[391], x[390], x[389], x[388], x[387], x[386], x[355]}), .y(y[77]));
  R1ind78 R1ind78_inst(.x({x[397], x[396], x[395], x[394], x[393], x[392], x[355]}), .y(y[78]));
  R1ind79 R1ind79_inst(.x({x[403], x[402], x[401], x[400], x[399], x[398], x[355]}), .y(y[79]));
  R1ind80 R1ind80_inst(.x({x[409], x[408], x[407], x[406], x[405], x[404], x[355]}), .y(y[80]));
  R1ind81 R1ind81_inst(.x({x[415], x[414], x[413], x[412], x[411], x[410], x[355]}), .y(y[81]));
  R1ind82 R1ind82_inst(.x({x[421], x[420], x[419], x[418], x[417], x[416], x[355]}), .y(y[82]));
  R1ind83 R1ind83_inst(.x({x[427], x[426], x[425], x[424], x[423], x[422], x[355]}), .y(y[83]));
  R1ind84 R1ind84_inst(.x({x[433], x[432], x[431], x[430], x[429], x[428], x[355]}), .y(y[84]));
  R1ind85 R1ind85_inst(.x({x[439], x[438], x[437], x[436], x[435], x[434], x[355]}), .y(y[85]));
  R1ind86 R1ind86_inst(.x({x[445], x[444], x[443], x[442], x[441], x[440], x[355]}), .y(y[86]));
  R1ind87 R1ind87_inst(.x({x[451], x[450], x[449], x[448], x[447], x[446], x[355]}), .y(y[87]));
  R1ind88 R1ind88_inst(.x({x[457], x[456], x[455], x[454], x[453], x[452], x[355]}), .y(y[88]));
  R1ind89 R1ind89_inst(.x({x[463], x[462], x[461], x[460], x[459], x[458], x[355]}), .y(y[89]));
  R1ind90 R1ind90_inst(.x({x[469], x[468], x[467], x[466], x[465], x[464], x[355]}), .y(y[90]));
  R1ind91 R1ind91_inst(.x({x[475], x[474], x[473], x[472], x[471], x[470], x[355]}), .y(y[91]));
  R1ind92 R1ind92_inst(.x({x[481], x[480], x[479], x[478], x[477], x[476], x[355]}), .y(y[92]));
  R1ind93 R1ind93_inst(.x({x[487], x[486], x[485], x[484], x[483], x[482], x[355]}), .y(y[93]));
  R1ind94 R1ind94_inst(.x({x[493], x[492], x[491], x[490], x[489], x[488], x[355]}), .y(y[94]));
  R1ind95 R1ind95_inst(.x({x[499], x[498], x[497], x[496], x[495], x[494], x[355]}), .y(y[95]));
  R1ind96 R1ind96_inst(.x({x[505], x[504], x[503], x[502], x[501], x[500], x[355]}), .y(y[96]));
  R1ind97 R1ind97_inst(.x({x[511], x[510], x[509], x[508], x[507], x[506], x[355]}), .y(y[97]));
  R1ind98 R1ind98_inst(.x({x[517], x[516], x[515], x[514], x[513], x[512], x[355]}), .y(y[98]));
  R1ind99 R1ind99_inst(.x({x[523], x[522], x[521], x[520], x[519], x[518], x[355]}), .y(y[99]));
  R1ind100 R1ind100_inst(.x({x[529], x[528], x[527], x[526], x[525], x[524], x[355]}), .y(y[100]));
  R1ind101 R1ind101_inst(.x({x[535], x[534], x[533], x[532], x[531], x[530], x[355]}), .y(y[101]));
  R1ind102 R1ind102_inst(.x({x[541], x[540], x[539], x[538], x[537], x[536], x[355]}), .y(y[102]));
  R1ind103 R1ind103_inst(.x({x[547], x[546], x[545], x[544], x[543], x[542], x[355]}), .y(y[103]));
  R1ind104 R1ind104_inst(.x({x[553], x[552], x[551], x[550], x[549], x[548], x[355]}), .y(y[104]));
  R1ind105 R1ind105_inst(.x({x[559], x[558], x[557], x[556], x[555], x[554], x[355]}), .y(y[105]));
  R1ind106 R1ind106_inst(.x({x[565], x[564], x[563], x[562], x[561], x[560], x[355]}), .y(y[106]));
  R1ind107 R1ind107_inst(.x({x[571], x[570], x[569], x[568], x[567], x[566], x[355]}), .y(y[107]));
  R1ind108 R1ind108_inst(.x({x[577], x[576], x[575], x[574], x[573], x[572], x[355]}), .y(y[108]));
  R1ind109 R1ind109_inst(.x({x[583], x[582], x[581], x[580], x[579], x[578], x[355]}), .y(y[109]));
  R1ind110 R1ind110_inst(.x({x[589], x[588], x[587], x[586], x[585], x[584], x[355]}), .y(y[110]));
  R1ind111 R1ind111_inst(.x({x[595], x[594], x[593], x[592], x[591], x[590], x[355]}), .y(y[111]));
  R1ind112 R1ind112_inst(.x({x[601], x[600], x[599], x[598], x[597], x[596], x[355]}), .y(y[112]));
  R1ind113 R1ind113_inst(.x({x[607], x[606], x[605], x[604], x[603], x[602], x[355]}), .y(y[113]));
  R1ind114 R1ind114_inst(.x({x[613], x[612], x[611], x[610], x[609], x[608], x[355]}), .y(y[114]));
  R1ind115 R1ind115_inst(.x({x[619], x[618], x[617], x[616], x[615], x[614], x[355]}), .y(y[115]));
  R1ind116 R1ind116_inst(.x({x[625], x[624], x[623], x[622], x[621], x[620], x[355]}), .y(y[116]));
  R1ind117 R1ind117_inst(.x({x[631], x[630], x[629], x[628], x[627], x[626], x[355]}), .y(y[117]));
  R1ind118 R1ind118_inst(.x({x[637], x[636], x[635], x[634], x[633], x[632], x[355]}), .y(y[118]));
  R1ind119 R1ind119_inst(.x({x[643], x[642], x[641], x[640], x[639], x[638], x[355]}), .y(y[119]));
  R1ind120 R1ind120_inst(.x({x[649], x[648], x[647], x[646], x[645], x[644], x[355]}), .y(y[120]));
  R1ind121 R1ind121_inst(.x({x[655], x[654], x[653], x[652], x[651], x[650], x[355]}), .y(y[121]));
  R1ind122 R1ind122_inst(.x({x[661], x[660], x[659], x[658], x[657], x[656], x[355]}), .y(y[122]));
  R1ind123 R1ind123_inst(.x({x[667], x[666], x[665], x[664], x[663], x[662], x[355]}), .y(y[123]));
  R1ind124 R1ind124_inst(.x({x[673], x[672], x[671], x[670], x[669], x[668], x[355]}), .y(y[124]));
  R1ind125 R1ind125_inst(.x({x[679], x[678], x[677], x[676], x[675], x[674], x[355]}), .y(y[125]));
  R1ind126 R1ind126_inst(.x({x[685], x[684], x[683], x[682], x[681], x[680], x[355]}), .y(y[126]));
  R1ind127 R1ind127_inst(.x({x[691], x[690], x[689], x[688], x[687], x[686], x[355]}), .y(y[127]));
  R1ind128 R1ind128_inst(.x({x[697], x[696], x[695], x[694], x[693], x[692], x[355]}), .y(y[128]));
  R1ind129 R1ind129_inst(.x({x[703], x[702], x[701], x[700], x[699], x[698], x[355]}), .y(y[129]));
  R1ind130 R1ind130_inst(.x({x[709], x[708], x[707], x[706], x[705], x[704], x[355]}), .y(y[130]));
  R1ind131 R1ind131_inst(.x({x[715], x[714], x[713], x[712], x[711], x[710], x[355]}), .y(y[131]));
  R1ind132 R1ind132_inst(.x({x[721], x[720], x[719], x[718], x[717], x[716], x[355]}), .y(y[132]));
  R1ind133 R1ind133_inst(.x({x[727], x[726], x[725], x[724], x[723], x[722], x[355]}), .y(y[133]));
  R1ind134 R1ind134_inst(.x({x[733], x[732], x[731], x[730], x[729], x[728], x[355]}), .y(y[134]));
  R1ind135 R1ind135_inst(.x({x[739], x[738], x[737], x[736], x[735], x[734], x[355]}), .y(y[135]));
  R1ind136 R1ind136_inst(.x({x[264], x[263], x[262], x[261], x[260], x[249], x[248], x[247], x[246], x[245], x[259], x[258], x[257], x[256], x[255], x[144], x[143], x[142], x[141], x[140], x[254], x[253], x[252], x[251], x[250], x[129], x[128], x[127], x[126], x[125], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[456], x[455], x[454], x[453], x[452], x[740], x[355]}), .y(y[136]));
  R1ind137 R1ind137_inst(.x({x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[256], x[255], x[249], x[248], x[247], x[246], x[245], x[144], x[143], x[142], x[141], x[140], x[254], x[253], x[252], x[251], x[250], x[139], x[138], x[137], x[136], x[135], x[129], x[128], x[127], x[126], x[125], x[134], x[133], x[132], x[131], x[130], x[462], x[461], x[460], x[459], x[458], x[741], x[355]}), .y(y[137]));
  R1ind138 R1ind138_inst(.x({x[254], x[253], x[252], x[251], x[250], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[256], x[255], x[134], x[133], x[132], x[131], x[130], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[468], x[467], x[466], x[465], x[464], x[742], x[355]}), .y(y[138]));
  R1ind139 R1ind139_inst(.x({x[264], x[263], x[262], x[261], x[260], x[254], x[253], x[252], x[251], x[250], x[259], x[258], x[257], x[256], x[255], x[249], x[248], x[247], x[246], x[245], x[144], x[143], x[142], x[141], x[140], x[134], x[133], x[132], x[131], x[130], x[139], x[138], x[137], x[136], x[135], x[129], x[128], x[127], x[126], x[125], x[474], x[473], x[472], x[471], x[470], x[743], x[355]}), .y(y[139]));
  R1ind140 R1ind140_inst(.x({x[284], x[283], x[282], x[281], x[280], x[269], x[268], x[267], x[266], x[265], x[279], x[278], x[277], x[276], x[275], x[164], x[163], x[162], x[161], x[160], x[274], x[273], x[272], x[271], x[270], x[149], x[148], x[147], x[146], x[145], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[480], x[479], x[478], x[477], x[476], x[744], x[355]}), .y(y[140]));
  R1ind141 R1ind141_inst(.x({x[284], x[283], x[282], x[281], x[280], x[164], x[163], x[162], x[161], x[160], x[279], x[278], x[277], x[276], x[275], x[269], x[268], x[267], x[266], x[265], x[274], x[273], x[272], x[271], x[270], x[159], x[158], x[157], x[156], x[155], x[149], x[148], x[147], x[146], x[145], x[154], x[153], x[152], x[151], x[150], x[486], x[485], x[484], x[483], x[482], x[745], x[355]}), .y(y[141]));
  R1ind142 R1ind142_inst(.x({x[274], x[273], x[272], x[271], x[270], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[277], x[276], x[275], x[154], x[153], x[152], x[151], x[150], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[155], x[492], x[491], x[490], x[489], x[488], x[746], x[355]}), .y(y[142]));
  R1ind143 R1ind143_inst(.x({x[284], x[283], x[282], x[281], x[280], x[274], x[273], x[272], x[271], x[270], x[279], x[278], x[277], x[276], x[275], x[269], x[268], x[267], x[266], x[265], x[164], x[163], x[162], x[161], x[160], x[154], x[153], x[152], x[151], x[150], x[159], x[158], x[157], x[156], x[155], x[149], x[148], x[147], x[146], x[145], x[498], x[497], x[496], x[495], x[494], x[747], x[355]}), .y(y[143]));
  R1ind144 R1ind144_inst(.x({x[304], x[303], x[302], x[301], x[300], x[289], x[288], x[287], x[286], x[285], x[299], x[298], x[297], x[296], x[295], x[104], x[103], x[102], x[101], x[100], x[294], x[293], x[292], x[291], x[290], x[89], x[88], x[87], x[86], x[85], x[99], x[98], x[97], x[96], x[95], x[94], x[93], x[92], x[91], x[90], x[504], x[503], x[502], x[501], x[500], x[748], x[355]}), .y(y[144]));
  R1ind145 R1ind145_inst(.x({x[304], x[303], x[302], x[301], x[300], x[299], x[298], x[297], x[296], x[295], x[289], x[288], x[287], x[286], x[285], x[104], x[103], x[102], x[101], x[100], x[294], x[293], x[292], x[291], x[290], x[99], x[98], x[97], x[96], x[95], x[89], x[88], x[87], x[86], x[85], x[94], x[93], x[92], x[91], x[90], x[510], x[509], x[508], x[507], x[506], x[749], x[355]}), .y(y[145]));
  R1ind146 R1ind146_inst(.x({x[294], x[293], x[292], x[291], x[290], x[304], x[303], x[302], x[301], x[300], x[299], x[298], x[297], x[296], x[295], x[94], x[93], x[92], x[91], x[90], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[516], x[515], x[514], x[513], x[512], x[750], x[355]}), .y(y[146]));
  R1ind147 R1ind147_inst(.x({x[304], x[303], x[302], x[301], x[300], x[294], x[293], x[292], x[291], x[290], x[299], x[298], x[297], x[296], x[295], x[289], x[288], x[287], x[286], x[285], x[104], x[103], x[102], x[101], x[100], x[94], x[93], x[92], x[91], x[90], x[99], x[98], x[97], x[96], x[95], x[89], x[88], x[87], x[86], x[85], x[522], x[521], x[520], x[519], x[518], x[751], x[355]}), .y(y[147]));
  R1ind148 R1ind148_inst(.x({x[324], x[323], x[322], x[321], x[320], x[309], x[308], x[307], x[306], x[305], x[319], x[318], x[317], x[316], x[315], x[314], x[313], x[312], x[311], x[310], x[124], x[123], x[122], x[121], x[120], x[109], x[108], x[107], x[106], x[105], x[119], x[118], x[117], x[116], x[115], x[354], x[353], x[352], x[351], x[350], x[114], x[113], x[112], x[111], x[110], x[528], x[527], x[526], x[525], x[524], x[752], x[355]}), .y(y[148]));
  R1ind149 R1ind149_inst(.x({x[324], x[323], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[309], x[308], x[307], x[306], x[305], x[314], x[313], x[312], x[311], x[310], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[109], x[108], x[107], x[106], x[105], x[339], x[338], x[337], x[336], x[335], x[114], x[113], x[112], x[111], x[110], x[534], x[533], x[532], x[531], x[530], x[753], x[355]}), .y(y[149]));
  R1ind150 R1ind150_inst(.x({x[314], x[313], x[312], x[311], x[310], x[324], x[323], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[114], x[113], x[112], x[111], x[110], x[344], x[343], x[342], x[341], x[340], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[540], x[539], x[538], x[537], x[536], x[754], x[355]}), .y(y[150]));
  R1ind151 R1ind151_inst(.x({x[324], x[323], x[322], x[321], x[320], x[314], x[313], x[312], x[311], x[310], x[319], x[318], x[317], x[316], x[315], x[309], x[308], x[307], x[306], x[305], x[124], x[123], x[122], x[121], x[120], x[114], x[113], x[112], x[111], x[110], x[119], x[118], x[117], x[116], x[115], x[109], x[108], x[107], x[106], x[105], x[349], x[348], x[347], x[346], x[345], x[546], x[545], x[544], x[543], x[542], x[755], x[355]}), .y(y[151]));
  R1ind152 R1ind152_inst(.x({x[204], x[203], x[202], x[201], x[200], x[189], x[188], x[187], x[186], x[185], x[199], x[198], x[197], x[196], x[195], x[144], x[143], x[142], x[141], x[140], x[194], x[193], x[192], x[191], x[190], x[129], x[128], x[127], x[126], x[125], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[384], x[383], x[382], x[381], x[380], x[756], x[355]}), .y(y[152]));
  R1ind153 R1ind153_inst(.x({x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[189], x[188], x[187], x[186], x[185], x[144], x[143], x[142], x[141], x[140], x[194], x[193], x[192], x[191], x[190], x[139], x[138], x[137], x[136], x[135], x[129], x[128], x[127], x[126], x[125], x[134], x[133], x[132], x[131], x[130], x[390], x[389], x[388], x[387], x[386], x[757], x[355]}), .y(y[153]));
  R1ind154 R1ind154_inst(.x({x[194], x[193], x[192], x[191], x[190], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[134], x[133], x[132], x[131], x[130], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[396], x[395], x[394], x[393], x[392], x[758], x[355]}), .y(y[154]));
  R1ind155 R1ind155_inst(.x({x[204], x[203], x[202], x[201], x[200], x[194], x[193], x[192], x[191], x[190], x[199], x[198], x[197], x[196], x[195], x[189], x[188], x[187], x[186], x[185], x[144], x[143], x[142], x[141], x[140], x[134], x[133], x[132], x[131], x[130], x[139], x[138], x[137], x[136], x[135], x[129], x[128], x[127], x[126], x[125], x[402], x[401], x[400], x[399], x[398], x[759], x[355]}), .y(y[155]));
  R1ind156 R1ind156_inst(.x({x[224], x[223], x[222], x[221], x[220], x[209], x[208], x[207], x[206], x[205], x[219], x[218], x[217], x[216], x[215], x[164], x[163], x[162], x[161], x[160], x[214], x[213], x[212], x[211], x[210], x[149], x[148], x[147], x[146], x[145], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[408], x[407], x[406], x[405], x[404], x[760], x[355]}), .y(y[156]));
  R1ind157 R1ind157_inst(.x({x[224], x[223], x[222], x[221], x[220], x[164], x[163], x[162], x[161], x[160], x[219], x[218], x[217], x[216], x[215], x[209], x[208], x[207], x[206], x[205], x[214], x[213], x[212], x[211], x[210], x[159], x[158], x[157], x[156], x[155], x[149], x[148], x[147], x[146], x[145], x[154], x[153], x[152], x[151], x[150], x[414], x[413], x[412], x[411], x[410], x[761], x[355]}), .y(y[157]));
  R1ind158 R1ind158_inst(.x({x[214], x[213], x[212], x[211], x[210], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[154], x[153], x[152], x[151], x[150], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[155], x[420], x[419], x[418], x[417], x[416], x[762], x[355]}), .y(y[158]));
  R1ind159 R1ind159_inst(.x({x[224], x[223], x[222], x[221], x[220], x[214], x[213], x[212], x[211], x[210], x[219], x[218], x[217], x[216], x[215], x[209], x[208], x[207], x[206], x[205], x[164], x[163], x[162], x[161], x[160], x[154], x[153], x[152], x[151], x[150], x[159], x[158], x[157], x[156], x[155], x[149], x[148], x[147], x[146], x[145], x[426], x[425], x[424], x[423], x[422], x[763], x[355]}), .y(y[159]));
  R1ind160 R1ind160_inst(.x({x[244], x[243], x[242], x[241], x[240], x[229], x[228], x[227], x[226], x[225], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[230], x[104], x[103], x[102], x[101], x[100], x[89], x[88], x[87], x[86], x[85], x[99], x[98], x[97], x[96], x[95], x[329], x[328], x[327], x[326], x[325], x[94], x[93], x[92], x[91], x[90], x[432], x[431], x[430], x[429], x[428], x[764], x[355]}), .y(y[160]));
  R1ind161 R1ind161_inst(.x({x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[235], x[229], x[228], x[227], x[226], x[225], x[234], x[233], x[232], x[231], x[230], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[89], x[88], x[87], x[86], x[85], x[334], x[333], x[332], x[331], x[330], x[94], x[93], x[92], x[91], x[90], x[438], x[437], x[436], x[435], x[434], x[765], x[355]}), .y(y[161]));
  R1ind162 R1ind162_inst(.x({x[234], x[233], x[232], x[231], x[230], x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[235], x[94], x[93], x[92], x[91], x[90], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[444], x[443], x[442], x[441], x[440], x[766], x[355]}), .y(y[162]));
  R1ind163 R1ind163_inst(.x({x[244], x[243], x[242], x[241], x[240], x[234], x[233], x[232], x[231], x[230], x[239], x[238], x[237], x[236], x[235], x[229], x[228], x[227], x[226], x[225], x[104], x[103], x[102], x[101], x[100], x[94], x[93], x[92], x[91], x[90], x[99], x[98], x[97], x[96], x[95], x[89], x[88], x[87], x[86], x[85], x[450], x[449], x[448], x[447], x[446], x[767], x[355]}), .y(y[163]));
  R1ind164 R1ind164_inst(.x({x[184], x[183], x[182], x[181], x[180], x[169], x[168], x[167], x[166], x[165], x[179], x[178], x[177], x[176], x[175], x[124], x[123], x[122], x[121], x[120], x[174], x[173], x[172], x[171], x[170], x[109], x[108], x[107], x[106], x[105], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[360], x[359], x[358], x[357], x[356], x[768], x[355]}), .y(y[164]));
  R1ind165 R1ind165_inst(.x({x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[169], x[168], x[167], x[166], x[165], x[124], x[123], x[122], x[121], x[120], x[174], x[173], x[172], x[171], x[170], x[119], x[118], x[117], x[116], x[115], x[109], x[108], x[107], x[106], x[105], x[114], x[113], x[112], x[111], x[110], x[366], x[365], x[364], x[363], x[362], x[769], x[355]}), .y(y[165]));
  R1ind166 R1ind166_inst(.x({x[174], x[173], x[172], x[171], x[170], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[114], x[113], x[112], x[111], x[110], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[372], x[371], x[370], x[369], x[368], x[770], x[355]}), .y(y[166]));
  R1ind167 R1ind167_inst(.x({x[184], x[183], x[182], x[181], x[180], x[174], x[173], x[172], x[171], x[170], x[179], x[178], x[177], x[176], x[175], x[169], x[168], x[167], x[166], x[165], x[124], x[123], x[122], x[121], x[120], x[114], x[113], x[112], x[111], x[110], x[119], x[118], x[117], x[116], x[115], x[109], x[108], x[107], x[106], x[105], x[378], x[377], x[376], x[375], x[374], x[771], x[355]}), .y(y[167]));
  R1ind168 R1ind168_inst(.x({x[264], x[263], x[262], x[261], x[260], x[249], x[248], x[247], x[246], x[245], x[259], x[258], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[456], x[455], x[454], x[453], x[452], x[772], x[355]}), .y(y[168]));
  R1ind169 R1ind169_inst(.x({x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[256], x[255], x[249], x[248], x[247], x[246], x[245], x[254], x[253], x[252], x[251], x[250], x[462], x[461], x[460], x[459], x[458], x[773], x[355]}), .y(y[169]));
  R1ind170 R1ind170_inst(.x({x[254], x[253], x[252], x[251], x[250], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[256], x[255], x[468], x[467], x[466], x[465], x[464], x[774], x[355]}), .y(y[170]));
  R1ind171 R1ind171_inst(.x({x[264], x[263], x[262], x[261], x[260], x[254], x[253], x[252], x[251], x[250], x[259], x[258], x[257], x[256], x[255], x[249], x[248], x[247], x[246], x[245], x[474], x[473], x[472], x[471], x[470], x[775], x[355]}), .y(y[171]));
  R1ind172 R1ind172_inst(.x({x[284], x[283], x[282], x[281], x[280], x[269], x[268], x[267], x[266], x[265], x[279], x[278], x[277], x[276], x[275], x[274], x[273], x[272], x[271], x[270], x[480], x[479], x[478], x[477], x[476], x[776], x[355]}), .y(y[172]));
  R1ind173 R1ind173_inst(.x({x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[277], x[276], x[275], x[269], x[268], x[267], x[266], x[265], x[274], x[273], x[272], x[271], x[270], x[486], x[485], x[484], x[483], x[482], x[777], x[355]}), .y(y[173]));
  R1ind174 R1ind174_inst(.x({x[274], x[273], x[272], x[271], x[270], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[277], x[276], x[275], x[492], x[491], x[490], x[489], x[488], x[778], x[355]}), .y(y[174]));
  R1ind175 R1ind175_inst(.x({x[284], x[283], x[282], x[281], x[280], x[274], x[273], x[272], x[271], x[270], x[279], x[278], x[277], x[276], x[275], x[269], x[268], x[267], x[266], x[265], x[498], x[497], x[496], x[495], x[494], x[779], x[355]}), .y(y[175]));
  R1ind176 R1ind176_inst(.x({x[304], x[303], x[302], x[301], x[300], x[289], x[288], x[287], x[286], x[285], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[292], x[291], x[290], x[504], x[503], x[502], x[501], x[500], x[780], x[355]}), .y(y[176]));
  R1ind177 R1ind177_inst(.x({x[304], x[303], x[302], x[301], x[300], x[299], x[298], x[297], x[296], x[295], x[289], x[288], x[287], x[286], x[285], x[294], x[293], x[292], x[291], x[290], x[510], x[509], x[508], x[507], x[506], x[781], x[355]}), .y(y[177]));
  R1ind178 R1ind178_inst(.x({x[294], x[293], x[292], x[291], x[290], x[304], x[303], x[302], x[301], x[300], x[299], x[298], x[297], x[296], x[295], x[516], x[515], x[514], x[513], x[512], x[782], x[355]}), .y(y[178]));
  R1ind179 R1ind179_inst(.x({x[304], x[303], x[302], x[301], x[300], x[294], x[293], x[292], x[291], x[290], x[299], x[298], x[297], x[296], x[295], x[289], x[288], x[287], x[286], x[285], x[522], x[521], x[520], x[519], x[518], x[783], x[355]}), .y(y[179]));
  R1ind180 R1ind180_inst(.x({x[324], x[323], x[322], x[321], x[320], x[309], x[308], x[307], x[306], x[305], x[319], x[318], x[317], x[316], x[315], x[314], x[313], x[312], x[311], x[310], x[354], x[353], x[352], x[351], x[350], x[528], x[527], x[526], x[525], x[524], x[784], x[355]}), .y(y[180]));
  R1ind181 R1ind181_inst(.x({x[324], x[323], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[309], x[308], x[307], x[306], x[305], x[314], x[313], x[312], x[311], x[310], x[339], x[338], x[337], x[336], x[335], x[534], x[533], x[532], x[531], x[530], x[785], x[355]}), .y(y[181]));
  R1ind182 R1ind182_inst(.x({x[314], x[313], x[312], x[311], x[310], x[324], x[323], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[344], x[343], x[342], x[341], x[340], x[540], x[539], x[538], x[537], x[536], x[786], x[355]}), .y(y[182]));
  R1ind183 R1ind183_inst(.x({x[324], x[323], x[322], x[321], x[320], x[314], x[313], x[312], x[311], x[310], x[319], x[318], x[317], x[316], x[315], x[309], x[308], x[307], x[306], x[305], x[349], x[348], x[347], x[346], x[345], x[546], x[545], x[544], x[543], x[542], x[787], x[355]}), .y(y[183]));
  R1ind184 R1ind184_inst(.x({x[264], x[263], x[262], x[261], x[260], x[84], x[83], x[82], x[81], x[80], x[144], x[143], x[142], x[141], x[140], x[249], x[248], x[247], x[246], x[245], x[259], x[258], x[257], x[256], x[255], x[69], x[68], x[67], x[66], x[65], x[79], x[78], x[77], x[76], x[75], x[129], x[128], x[127], x[126], x[125], x[139], x[138], x[137], x[136], x[135], x[254], x[253], x[252], x[251], x[250], x[74], x[73], x[72], x[71], x[70], x[134], x[133], x[132], x[131], x[130], x[456], x[455], x[454], x[453], x[452], x[788], x[355]}), .y(y[184]));
  R1ind185 R1ind185_inst(.x({x[264], x[263], x[262], x[261], x[260], x[84], x[83], x[82], x[81], x[80], x[144], x[143], x[142], x[141], x[140], x[259], x[258], x[257], x[256], x[255], x[249], x[248], x[247], x[246], x[245], x[79], x[78], x[77], x[76], x[75], x[69], x[68], x[67], x[66], x[65], x[139], x[138], x[137], x[136], x[135], x[129], x[128], x[127], x[126], x[125], x[254], x[253], x[252], x[251], x[250], x[74], x[73], x[72], x[71], x[70], x[134], x[133], x[132], x[131], x[130], x[462], x[461], x[460], x[459], x[458], x[789], x[355]}), .y(y[185]));
  R1ind186 R1ind186_inst(.x({x[254], x[253], x[252], x[251], x[250], x[74], x[73], x[72], x[71], x[70], x[134], x[133], x[132], x[131], x[130], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[256], x[255], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[468], x[467], x[466], x[465], x[464], x[790], x[355]}), .y(y[186]));
  R1ind187 R1ind187_inst(.x({x[264], x[263], x[262], x[261], x[260], x[84], x[83], x[82], x[81], x[80], x[144], x[143], x[142], x[141], x[140], x[254], x[253], x[252], x[251], x[250], x[259], x[258], x[257], x[256], x[255], x[249], x[248], x[247], x[246], x[245], x[74], x[73], x[72], x[71], x[70], x[79], x[78], x[77], x[76], x[75], x[69], x[68], x[67], x[66], x[65], x[134], x[133], x[132], x[131], x[130], x[139], x[138], x[137], x[136], x[135], x[129], x[128], x[127], x[126], x[125], x[474], x[473], x[472], x[471], x[470], x[791], x[355]}), .y(y[187]));
  R1ind188 R1ind188_inst(.x({x[284], x[283], x[282], x[281], x[280], x[24], x[23], x[22], x[21], x[20], x[164], x[163], x[162], x[161], x[160], x[269], x[268], x[267], x[266], x[265], x[279], x[278], x[277], x[276], x[275], x[9], x[8], x[7], x[6], x[5], x[19], x[18], x[17], x[16], x[15], x[149], x[148], x[147], x[146], x[145], x[159], x[158], x[157], x[156], x[155], x[274], x[273], x[272], x[271], x[270], x[14], x[13], x[12], x[11], x[10], x[154], x[153], x[152], x[151], x[150], x[480], x[479], x[478], x[477], x[476], x[792], x[355]}), .y(y[188]));
  R1ind189 R1ind189_inst(.x({x[164], x[163], x[162], x[161], x[160], x[284], x[283], x[282], x[281], x[280], x[24], x[23], x[22], x[21], x[20], x[159], x[158], x[157], x[156], x[155], x[149], x[148], x[147], x[146], x[145], x[279], x[278], x[277], x[276], x[275], x[269], x[268], x[267], x[266], x[265], x[19], x[18], x[17], x[16], x[15], x[9], x[8], x[7], x[6], x[5], x[154], x[153], x[152], x[151], x[150], x[274], x[273], x[272], x[271], x[270], x[14], x[13], x[12], x[11], x[10], x[486], x[485], x[484], x[483], x[482], x[793], x[355]}), .y(y[189]));
  R1ind190 R1ind190_inst(.x({x[274], x[273], x[272], x[271], x[270], x[14], x[13], x[12], x[11], x[10], x[154], x[153], x[152], x[151], x[150], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[277], x[276], x[275], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[155], x[492], x[491], x[490], x[489], x[488], x[794], x[355]}), .y(y[190]));
  R1ind191 R1ind191_inst(.x({x[284], x[283], x[282], x[281], x[280], x[24], x[23], x[22], x[21], x[20], x[164], x[163], x[162], x[161], x[160], x[274], x[273], x[272], x[271], x[270], x[279], x[278], x[277], x[276], x[275], x[269], x[268], x[267], x[266], x[265], x[14], x[13], x[12], x[11], x[10], x[19], x[18], x[17], x[16], x[15], x[9], x[8], x[7], x[6], x[5], x[154], x[153], x[152], x[151], x[150], x[159], x[158], x[157], x[156], x[155], x[149], x[148], x[147], x[146], x[145], x[498], x[497], x[496], x[495], x[494], x[795], x[355]}), .y(y[191]));
  R1ind192 R1ind192_inst(.x({x[304], x[303], x[302], x[301], x[300], x[44], x[43], x[42], x[41], x[40], x[104], x[103], x[102], x[101], x[100], x[289], x[288], x[287], x[286], x[285], x[299], x[298], x[297], x[296], x[295], x[29], x[28], x[27], x[26], x[25], x[39], x[38], x[37], x[36], x[35], x[89], x[88], x[87], x[86], x[85], x[99], x[98], x[97], x[96], x[95], x[294], x[293], x[292], x[291], x[290], x[34], x[33], x[32], x[31], x[30], x[94], x[93], x[92], x[91], x[90], x[504], x[503], x[502], x[501], x[500], x[796], x[355]}), .y(y[192]));
  R1ind193 R1ind193_inst(.x({x[304], x[303], x[302], x[301], x[300], x[44], x[43], x[42], x[41], x[40], x[104], x[103], x[102], x[101], x[100], x[299], x[298], x[297], x[296], x[295], x[289], x[288], x[287], x[286], x[285], x[39], x[38], x[37], x[36], x[35], x[29], x[28], x[27], x[26], x[25], x[99], x[98], x[97], x[96], x[95], x[89], x[88], x[87], x[86], x[85], x[294], x[293], x[292], x[291], x[290], x[34], x[33], x[32], x[31], x[30], x[94], x[93], x[92], x[91], x[90], x[510], x[509], x[508], x[507], x[506], x[797], x[355]}), .y(y[193]));
  R1ind194 R1ind194_inst(.x({x[294], x[293], x[292], x[291], x[290], x[34], x[33], x[32], x[31], x[30], x[94], x[93], x[92], x[91], x[90], x[304], x[303], x[302], x[301], x[300], x[299], x[298], x[297], x[296], x[295], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[516], x[515], x[514], x[513], x[512], x[798], x[355]}), .y(y[194]));
  R1ind195 R1ind195_inst(.x({x[304], x[303], x[302], x[301], x[300], x[44], x[43], x[42], x[41], x[40], x[104], x[103], x[102], x[101], x[100], x[294], x[293], x[292], x[291], x[290], x[299], x[298], x[297], x[296], x[295], x[289], x[288], x[287], x[286], x[285], x[34], x[33], x[32], x[31], x[30], x[39], x[38], x[37], x[36], x[35], x[29], x[28], x[27], x[26], x[25], x[94], x[93], x[92], x[91], x[90], x[99], x[98], x[97], x[96], x[95], x[89], x[88], x[87], x[86], x[85], x[522], x[521], x[520], x[519], x[518], x[799], x[355]}), .y(y[195]));
  R1ind196 R1ind196_inst(.x({x[324], x[323], x[322], x[321], x[320], x[309], x[308], x[307], x[306], x[305], x[319], x[318], x[317], x[316], x[315], x[64], x[63], x[62], x[61], x[60], x[124], x[123], x[122], x[121], x[120], x[314], x[313], x[312], x[311], x[310], x[49], x[48], x[47], x[46], x[45], x[59], x[58], x[57], x[56], x[55], x[109], x[108], x[107], x[106], x[105], x[119], x[118], x[117], x[116], x[115], x[54], x[53], x[52], x[51], x[50], x[114], x[113], x[112], x[111], x[110], x[354], x[353], x[352], x[351], x[350], x[528], x[527], x[526], x[525], x[524], x[800], x[355]}), .y(y[196]));
  R1ind197 R1ind197_inst(.x({x[324], x[323], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[309], x[308], x[307], x[306], x[305], x[64], x[63], x[62], x[61], x[60], x[124], x[123], x[122], x[121], x[120], x[314], x[313], x[312], x[311], x[310], x[59], x[58], x[57], x[56], x[55], x[49], x[48], x[47], x[46], x[45], x[119], x[118], x[117], x[116], x[115], x[109], x[108], x[107], x[106], x[105], x[54], x[53], x[52], x[51], x[50], x[114], x[113], x[112], x[111], x[110], x[339], x[338], x[337], x[336], x[335], x[534], x[533], x[532], x[531], x[530], x[801], x[355]}), .y(y[197]));
  R1ind198 R1ind198_inst(.x({x[314], x[313], x[312], x[311], x[310], x[324], x[323], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[54], x[53], x[52], x[51], x[50], x[114], x[113], x[112], x[111], x[110], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[344], x[343], x[342], x[341], x[340], x[540], x[539], x[538], x[537], x[536], x[802], x[355]}), .y(y[198]));
  R1ind199 R1ind199_inst(.x({x[324], x[323], x[322], x[321], x[320], x[314], x[313], x[312], x[311], x[310], x[319], x[318], x[317], x[316], x[315], x[309], x[308], x[307], x[306], x[305], x[64], x[63], x[62], x[61], x[60], x[124], x[123], x[122], x[121], x[120], x[54], x[53], x[52], x[51], x[50], x[59], x[58], x[57], x[56], x[55], x[49], x[48], x[47], x[46], x[45], x[114], x[113], x[112], x[111], x[110], x[119], x[118], x[117], x[116], x[115], x[109], x[108], x[107], x[106], x[105], x[349], x[348], x[347], x[346], x[345], x[546], x[545], x[544], x[543], x[542], x[803], x[355]}), .y(y[199]));
endmodule

module R2ind0(x, y);
 input [4:0] x;
 output y;

 wire [9:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (~t[2] & t[3] & t[4] & t[5]) | (t[2] & ~t[4] & ~t[5]) | (t[2] & ~t[3] & ~t[5]) | (t[2] & ~t[3] & ~t[4]);
  assign t[2] = t[6] ^ x[4];
  assign t[3] = t[7] ^ x[1];
  assign t[4] = t[8] ^ x[2];
  assign t[5] = t[9] ^ x[3];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign t[8] = (x[0]);
  assign t[9] = (x[0]);
  assign y = t[0];
endmodule

module R2ind1(x, y);
 input [4:0] x;
 output y;

 wire [9:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (t[2] & ~t[3] & t[4] & t[5]) | (t[3] & ~t[4] & ~t[5]) | (~t[2] & t[3] & ~t[5]) | (~t[2] & t[3] & ~t[4]);
  assign t[2] = t[6] ^ x[1];
  assign t[3] = t[7] ^ x[4];
  assign t[4] = t[8] ^ x[2];
  assign t[5] = t[9] ^ x[3];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign t[8] = (x[0]);
  assign t[9] = (x[0]);
  assign y = t[0];
endmodule

module R2ind2(x, y);
 input [4:0] x;
 output y;

 wire [9:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (t[2] & t[3] & ~t[4] & t[5]) | (~t[3] & t[4] & ~t[5]) | (~t[2] & t[4] & ~t[5]) | (~t[2] & ~t[3] & t[4]);
  assign t[2] = t[6] ^ x[1];
  assign t[3] = t[7] ^ x[2];
  assign t[4] = t[8] ^ x[4];
  assign t[5] = t[9] ^ x[3];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign t[8] = (x[0]);
  assign t[9] = (x[0]);
  assign y = t[0];
endmodule

module R2ind3(x, y);
 input [4:0] x;
 output y;

 wire [9:0] t;
  assign t[0] = t[1] ^ x[4];
  assign t[1] = (t[2] & t[3] & t[4] & ~t[5]) | (~t[3] & ~t[4] & t[5]) | (~t[2] & ~t[4] & t[5]) | (~t[2] & ~t[3] & t[5]);
  assign t[2] = t[6] ^ x[1];
  assign t[3] = t[7] ^ x[2];
  assign t[4] = t[8] ^ x[3];
  assign t[5] = t[9] ^ x[4];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign t[8] = (x[0]);
  assign t[9] = (x[0]);
  assign y = t[0];
endmodule

module R2ind4(x, y);
 input [29:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[4];
  assign t[13] = t[19] ^ x[9];
  assign t[14] = t[20] ^ x[14];
  assign t[15] = t[21] ^ x[19];
  assign t[16] = t[22] ^ x[24];
  assign t[17] = t[23] ^ x[29];
  assign t[18] = (~t[24] & t[25] & t[26] & t[27]) | (t[24] & ~t[26] & ~t[27]) | (t[24] & ~t[25] & ~t[27]) | (t[24] & ~t[25] & ~t[26]);
  assign t[19] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[21] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[22] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[23] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[24] = t[48] ^ x[4];
  assign t[25] = t[49] ^ x[1];
  assign t[26] = t[50] ^ x[2];
  assign t[27] = t[51] ^ x[3];
  assign t[28] = t[52] ^ x[9];
  assign t[29] = t[53] ^ x[6];
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[54] ^ x[7];
  assign t[31] = t[55] ^ x[8];
  assign t[32] = t[56] ^ x[14];
  assign t[33] = t[57] ^ x[11];
  assign t[34] = t[58] ^ x[12];
  assign t[35] = t[59] ^ x[13];
  assign t[36] = t[60] ^ x[19];
  assign t[37] = t[61] ^ x[16];
  assign t[38] = t[62] ^ x[17];
  assign t[39] = t[63] ^ x[18];
  assign t[3] = ~(t[8] | t[9]);
  assign t[40] = t[64] ^ x[24];
  assign t[41] = t[65] ^ x[21];
  assign t[42] = t[66] ^ x[22];
  assign t[43] = t[67] ^ x[23];
  assign t[44] = t[68] ^ x[29];
  assign t[45] = t[69] ^ x[26];
  assign t[46] = t[70] ^ x[27];
  assign t[47] = t[71] ^ x[28];
  assign t[48] = (x[0]);
  assign t[49] = (x[0]);
  assign t[4] = ~(t[10] | t[5]);
  assign t[50] = (x[0]);
  assign t[51] = (x[0]);
  assign t[52] = (x[5]);
  assign t[53] = (x[5]);
  assign t[54] = (x[5]);
  assign t[55] = (x[5]);
  assign t[56] = (x[10]);
  assign t[57] = (x[10]);
  assign t[58] = (x[10]);
  assign t[59] = (x[10]);
  assign t[5] = ~(t[11]);
  assign t[60] = (x[15]);
  assign t[61] = (x[15]);
  assign t[62] = (x[15]);
  assign t[63] = (x[15]);
  assign t[64] = (x[20]);
  assign t[65] = (x[20]);
  assign t[66] = (x[20]);
  assign t[67] = (x[20]);
  assign t[68] = (x[25]);
  assign t[69] = (x[25]);
  assign t[6] = (t[12]);
  assign t[70] = (x[25]);
  assign t[71] = (x[25]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind5(x, y);
 input [29:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[4];
  assign t[13] = t[19] ^ x[9];
  assign t[14] = t[20] ^ x[14];
  assign t[15] = t[21] ^ x[19];
  assign t[16] = t[22] ^ x[24];
  assign t[17] = t[23] ^ x[29];
  assign t[18] = (~t[24] & t[25] & t[26] & t[27]) | (t[24] & ~t[26] & ~t[27]) | (t[24] & ~t[25] & ~t[27]) | (t[24] & ~t[25] & ~t[26]);
  assign t[19] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[21] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[22] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[23] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[24] = t[48] ^ x[4];
  assign t[25] = t[49] ^ x[1];
  assign t[26] = t[50] ^ x[2];
  assign t[27] = t[51] ^ x[3];
  assign t[28] = t[52] ^ x[9];
  assign t[29] = t[53] ^ x[6];
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[54] ^ x[7];
  assign t[31] = t[55] ^ x[8];
  assign t[32] = t[56] ^ x[14];
  assign t[33] = t[57] ^ x[11];
  assign t[34] = t[58] ^ x[12];
  assign t[35] = t[59] ^ x[13];
  assign t[36] = t[60] ^ x[19];
  assign t[37] = t[61] ^ x[16];
  assign t[38] = t[62] ^ x[17];
  assign t[39] = t[63] ^ x[18];
  assign t[3] = ~(t[8] | t[9]);
  assign t[40] = t[64] ^ x[24];
  assign t[41] = t[65] ^ x[21];
  assign t[42] = t[66] ^ x[22];
  assign t[43] = t[67] ^ x[23];
  assign t[44] = t[68] ^ x[29];
  assign t[45] = t[69] ^ x[26];
  assign t[46] = t[70] ^ x[27];
  assign t[47] = t[71] ^ x[28];
  assign t[48] = (x[0]);
  assign t[49] = (x[0]);
  assign t[4] = ~(t[10] | t[5]);
  assign t[50] = (x[0]);
  assign t[51] = (x[0]);
  assign t[52] = (x[5]);
  assign t[53] = (x[5]);
  assign t[54] = (x[5]);
  assign t[55] = (x[5]);
  assign t[56] = (x[10]);
  assign t[57] = (x[10]);
  assign t[58] = (x[10]);
  assign t[59] = (x[10]);
  assign t[5] = ~(t[11]);
  assign t[60] = (x[15]);
  assign t[61] = (x[15]);
  assign t[62] = (x[15]);
  assign t[63] = (x[15]);
  assign t[64] = (x[20]);
  assign t[65] = (x[20]);
  assign t[66] = (x[20]);
  assign t[67] = (x[20]);
  assign t[68] = (x[25]);
  assign t[69] = (x[25]);
  assign t[6] = (t[12]);
  assign t[70] = (x[25]);
  assign t[71] = (x[25]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind6(x, y);
 input [29:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[4];
  assign t[13] = t[19] ^ x[9];
  assign t[14] = t[20] ^ x[14];
  assign t[15] = t[21] ^ x[19];
  assign t[16] = t[22] ^ x[24];
  assign t[17] = t[23] ^ x[29];
  assign t[18] = (~t[24] & t[25] & t[26] & t[27]) | (t[24] & ~t[26] & ~t[27]) | (t[24] & ~t[25] & ~t[27]) | (t[24] & ~t[25] & ~t[26]);
  assign t[19] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[21] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[22] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[23] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[24] = t[48] ^ x[4];
  assign t[25] = t[49] ^ x[1];
  assign t[26] = t[50] ^ x[2];
  assign t[27] = t[51] ^ x[3];
  assign t[28] = t[52] ^ x[9];
  assign t[29] = t[53] ^ x[6];
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[54] ^ x[7];
  assign t[31] = t[55] ^ x[8];
  assign t[32] = t[56] ^ x[14];
  assign t[33] = t[57] ^ x[11];
  assign t[34] = t[58] ^ x[12];
  assign t[35] = t[59] ^ x[13];
  assign t[36] = t[60] ^ x[19];
  assign t[37] = t[61] ^ x[16];
  assign t[38] = t[62] ^ x[17];
  assign t[39] = t[63] ^ x[18];
  assign t[3] = ~(t[8] | t[9]);
  assign t[40] = t[64] ^ x[24];
  assign t[41] = t[65] ^ x[21];
  assign t[42] = t[66] ^ x[22];
  assign t[43] = t[67] ^ x[23];
  assign t[44] = t[68] ^ x[29];
  assign t[45] = t[69] ^ x[26];
  assign t[46] = t[70] ^ x[27];
  assign t[47] = t[71] ^ x[28];
  assign t[48] = (x[0]);
  assign t[49] = (x[0]);
  assign t[4] = ~(t[10] | t[5]);
  assign t[50] = (x[0]);
  assign t[51] = (x[0]);
  assign t[52] = (x[5]);
  assign t[53] = (x[5]);
  assign t[54] = (x[5]);
  assign t[55] = (x[5]);
  assign t[56] = (x[10]);
  assign t[57] = (x[10]);
  assign t[58] = (x[10]);
  assign t[59] = (x[10]);
  assign t[5] = ~(t[11]);
  assign t[60] = (x[15]);
  assign t[61] = (x[15]);
  assign t[62] = (x[15]);
  assign t[63] = (x[15]);
  assign t[64] = (x[20]);
  assign t[65] = (x[20]);
  assign t[66] = (x[20]);
  assign t[67] = (x[20]);
  assign t[68] = (x[25]);
  assign t[69] = (x[25]);
  assign t[6] = (t[12]);
  assign t[70] = (x[25]);
  assign t[71] = (x[25]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind7(x, y);
 input [29:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[4];
  assign t[13] = t[19] ^ x[9];
  assign t[14] = t[20] ^ x[14];
  assign t[15] = t[21] ^ x[19];
  assign t[16] = t[22] ^ x[24];
  assign t[17] = t[23] ^ x[29];
  assign t[18] = (~t[24] & t[25] & t[26] & t[27]) | (t[24] & ~t[26] & ~t[27]) | (t[24] & ~t[25] & ~t[27]) | (t[24] & ~t[25] & ~t[26]);
  assign t[19] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[21] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[22] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[23] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[24] = t[48] ^ x[4];
  assign t[25] = t[49] ^ x[1];
  assign t[26] = t[50] ^ x[2];
  assign t[27] = t[51] ^ x[3];
  assign t[28] = t[52] ^ x[9];
  assign t[29] = t[53] ^ x[6];
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[54] ^ x[7];
  assign t[31] = t[55] ^ x[8];
  assign t[32] = t[56] ^ x[14];
  assign t[33] = t[57] ^ x[11];
  assign t[34] = t[58] ^ x[12];
  assign t[35] = t[59] ^ x[13];
  assign t[36] = t[60] ^ x[19];
  assign t[37] = t[61] ^ x[16];
  assign t[38] = t[62] ^ x[17];
  assign t[39] = t[63] ^ x[18];
  assign t[3] = ~(t[8] | t[9]);
  assign t[40] = t[64] ^ x[24];
  assign t[41] = t[65] ^ x[21];
  assign t[42] = t[66] ^ x[22];
  assign t[43] = t[67] ^ x[23];
  assign t[44] = t[68] ^ x[29];
  assign t[45] = t[69] ^ x[26];
  assign t[46] = t[70] ^ x[27];
  assign t[47] = t[71] ^ x[28];
  assign t[48] = (x[0]);
  assign t[49] = (x[0]);
  assign t[4] = ~(t[10] | t[5]);
  assign t[50] = (x[0]);
  assign t[51] = (x[0]);
  assign t[52] = (x[5]);
  assign t[53] = (x[5]);
  assign t[54] = (x[5]);
  assign t[55] = (x[5]);
  assign t[56] = (x[10]);
  assign t[57] = (x[10]);
  assign t[58] = (x[10]);
  assign t[59] = (x[10]);
  assign t[5] = ~(t[11]);
  assign t[60] = (x[15]);
  assign t[61] = (x[15]);
  assign t[62] = (x[15]);
  assign t[63] = (x[15]);
  assign t[64] = (x[20]);
  assign t[65] = (x[20]);
  assign t[66] = (x[20]);
  assign t[67] = (x[20]);
  assign t[68] = (x[25]);
  assign t[69] = (x[25]);
  assign t[6] = (t[12]);
  assign t[70] = (x[25]);
  assign t[71] = (x[25]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind8(x, y);
 input [30:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(~x[0] & ~t[1]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[5];
  assign t[13] = t[19] ^ x[10];
  assign t[14] = t[20] ^ x[15];
  assign t[15] = t[21] ^ x[20];
  assign t[16] = t[22] ^ x[25];
  assign t[17] = t[23] ^ x[30];
  assign t[18] = (~t[24] & t[25] & t[26] & t[27]) | (t[24] & ~t[26] & ~t[27]) | (t[24] & ~t[25] & ~t[27]) | (t[24] & ~t[25] & ~t[26]);
  assign t[19] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[1] = t[6] ? t[7] : t[2];
  assign t[20] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[21] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[22] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[23] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[24] = t[48] ^ x[5];
  assign t[25] = t[49] ^ x[2];
  assign t[26] = t[50] ^ x[3];
  assign t[27] = t[51] ^ x[4];
  assign t[28] = t[52] ^ x[10];
  assign t[29] = t[53] ^ x[7];
  assign t[2] = ~(t[7] & t[3]);
  assign t[30] = t[54] ^ x[8];
  assign t[31] = t[55] ^ x[9];
  assign t[32] = t[56] ^ x[15];
  assign t[33] = t[57] ^ x[12];
  assign t[34] = t[58] ^ x[13];
  assign t[35] = t[59] ^ x[14];
  assign t[36] = t[60] ^ x[20];
  assign t[37] = t[61] ^ x[17];
  assign t[38] = t[62] ^ x[18];
  assign t[39] = t[63] ^ x[19];
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = t[64] ^ x[25];
  assign t[41] = t[65] ^ x[22];
  assign t[42] = t[66] ^ x[23];
  assign t[43] = t[67] ^ x[24];
  assign t[44] = t[68] ^ x[30];
  assign t[45] = t[69] ^ x[27];
  assign t[46] = t[70] ^ x[28];
  assign t[47] = t[71] ^ x[29];
  assign t[48] = (x[1]);
  assign t[49] = (x[1]);
  assign t[4] = t[8] & t[9];
  assign t[50] = (x[1]);
  assign t[51] = (x[1]);
  assign t[52] = (x[6]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[6]);
  assign t[56] = (x[11]);
  assign t[57] = (x[11]);
  assign t[58] = (x[11]);
  assign t[59] = (x[11]);
  assign t[5] = ~(t[10] | t[11]);
  assign t[60] = (x[16]);
  assign t[61] = (x[16]);
  assign t[62] = (x[16]);
  assign t[63] = (x[16]);
  assign t[64] = (x[21]);
  assign t[65] = (x[21]);
  assign t[66] = (x[21]);
  assign t[67] = (x[21]);
  assign t[68] = (x[26]);
  assign t[69] = (x[26]);
  assign t[6] = (t[12]);
  assign t[70] = (x[26]);
  assign t[71] = (x[26]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind9(x, y);
 input [30:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(~x[0] & ~t[1]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[5];
  assign t[13] = t[19] ^ x[10];
  assign t[14] = t[20] ^ x[15];
  assign t[15] = t[21] ^ x[20];
  assign t[16] = t[22] ^ x[25];
  assign t[17] = t[23] ^ x[30];
  assign t[18] = (~t[24] & t[25] & t[26] & t[27]) | (t[24] & ~t[26] & ~t[27]) | (t[24] & ~t[25] & ~t[27]) | (t[24] & ~t[25] & ~t[26]);
  assign t[19] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[1] = t[6] ? t[7] : t[2];
  assign t[20] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[21] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[22] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[23] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[24] = t[48] ^ x[5];
  assign t[25] = t[49] ^ x[2];
  assign t[26] = t[50] ^ x[3];
  assign t[27] = t[51] ^ x[4];
  assign t[28] = t[52] ^ x[10];
  assign t[29] = t[53] ^ x[7];
  assign t[2] = ~(t[7] & t[3]);
  assign t[30] = t[54] ^ x[8];
  assign t[31] = t[55] ^ x[9];
  assign t[32] = t[56] ^ x[15];
  assign t[33] = t[57] ^ x[12];
  assign t[34] = t[58] ^ x[13];
  assign t[35] = t[59] ^ x[14];
  assign t[36] = t[60] ^ x[20];
  assign t[37] = t[61] ^ x[17];
  assign t[38] = t[62] ^ x[18];
  assign t[39] = t[63] ^ x[19];
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = t[64] ^ x[25];
  assign t[41] = t[65] ^ x[22];
  assign t[42] = t[66] ^ x[23];
  assign t[43] = t[67] ^ x[24];
  assign t[44] = t[68] ^ x[30];
  assign t[45] = t[69] ^ x[27];
  assign t[46] = t[70] ^ x[28];
  assign t[47] = t[71] ^ x[29];
  assign t[48] = (x[1]);
  assign t[49] = (x[1]);
  assign t[4] = t[8] & t[9];
  assign t[50] = (x[1]);
  assign t[51] = (x[1]);
  assign t[52] = (x[6]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[6]);
  assign t[56] = (x[11]);
  assign t[57] = (x[11]);
  assign t[58] = (x[11]);
  assign t[59] = (x[11]);
  assign t[5] = ~(t[10] | t[11]);
  assign t[60] = (x[16]);
  assign t[61] = (x[16]);
  assign t[62] = (x[16]);
  assign t[63] = (x[16]);
  assign t[64] = (x[21]);
  assign t[65] = (x[21]);
  assign t[66] = (x[21]);
  assign t[67] = (x[21]);
  assign t[68] = (x[26]);
  assign t[69] = (x[26]);
  assign t[6] = (t[12]);
  assign t[70] = (x[26]);
  assign t[71] = (x[26]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind10(x, y);
 input [30:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(~x[0] & ~t[1]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[5];
  assign t[13] = t[19] ^ x[10];
  assign t[14] = t[20] ^ x[15];
  assign t[15] = t[21] ^ x[20];
  assign t[16] = t[22] ^ x[25];
  assign t[17] = t[23] ^ x[30];
  assign t[18] = (~t[24] & t[25] & t[26] & t[27]) | (t[24] & ~t[26] & ~t[27]) | (t[24] & ~t[25] & ~t[27]) | (t[24] & ~t[25] & ~t[26]);
  assign t[19] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[1] = t[6] ? t[7] : t[2];
  assign t[20] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[21] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[22] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[23] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[24] = t[48] ^ x[5];
  assign t[25] = t[49] ^ x[2];
  assign t[26] = t[50] ^ x[3];
  assign t[27] = t[51] ^ x[4];
  assign t[28] = t[52] ^ x[10];
  assign t[29] = t[53] ^ x[7];
  assign t[2] = ~(t[7] & t[3]);
  assign t[30] = t[54] ^ x[8];
  assign t[31] = t[55] ^ x[9];
  assign t[32] = t[56] ^ x[15];
  assign t[33] = t[57] ^ x[12];
  assign t[34] = t[58] ^ x[13];
  assign t[35] = t[59] ^ x[14];
  assign t[36] = t[60] ^ x[20];
  assign t[37] = t[61] ^ x[17];
  assign t[38] = t[62] ^ x[18];
  assign t[39] = t[63] ^ x[19];
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = t[64] ^ x[25];
  assign t[41] = t[65] ^ x[22];
  assign t[42] = t[66] ^ x[23];
  assign t[43] = t[67] ^ x[24];
  assign t[44] = t[68] ^ x[30];
  assign t[45] = t[69] ^ x[27];
  assign t[46] = t[70] ^ x[28];
  assign t[47] = t[71] ^ x[29];
  assign t[48] = (x[1]);
  assign t[49] = (x[1]);
  assign t[4] = t[8] & t[9];
  assign t[50] = (x[1]);
  assign t[51] = (x[1]);
  assign t[52] = (x[6]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[6]);
  assign t[56] = (x[11]);
  assign t[57] = (x[11]);
  assign t[58] = (x[11]);
  assign t[59] = (x[11]);
  assign t[5] = ~(t[10] | t[11]);
  assign t[60] = (x[16]);
  assign t[61] = (x[16]);
  assign t[62] = (x[16]);
  assign t[63] = (x[16]);
  assign t[64] = (x[21]);
  assign t[65] = (x[21]);
  assign t[66] = (x[21]);
  assign t[67] = (x[21]);
  assign t[68] = (x[26]);
  assign t[69] = (x[26]);
  assign t[6] = (t[12]);
  assign t[70] = (x[26]);
  assign t[71] = (x[26]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind11(x, y);
 input [30:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(~x[0] & ~t[1]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[5];
  assign t[13] = t[19] ^ x[10];
  assign t[14] = t[20] ^ x[15];
  assign t[15] = t[21] ^ x[20];
  assign t[16] = t[22] ^ x[25];
  assign t[17] = t[23] ^ x[30];
  assign t[18] = (~t[24] & t[25] & t[26] & t[27]) | (t[24] & ~t[26] & ~t[27]) | (t[24] & ~t[25] & ~t[27]) | (t[24] & ~t[25] & ~t[26]);
  assign t[19] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[1] = t[6] ? t[7] : t[2];
  assign t[20] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[21] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[22] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[23] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[24] = t[48] ^ x[5];
  assign t[25] = t[49] ^ x[2];
  assign t[26] = t[50] ^ x[3];
  assign t[27] = t[51] ^ x[4];
  assign t[28] = t[52] ^ x[10];
  assign t[29] = t[53] ^ x[7];
  assign t[2] = ~(t[7] & t[3]);
  assign t[30] = t[54] ^ x[8];
  assign t[31] = t[55] ^ x[9];
  assign t[32] = t[56] ^ x[15];
  assign t[33] = t[57] ^ x[12];
  assign t[34] = t[58] ^ x[13];
  assign t[35] = t[59] ^ x[14];
  assign t[36] = t[60] ^ x[20];
  assign t[37] = t[61] ^ x[17];
  assign t[38] = t[62] ^ x[18];
  assign t[39] = t[63] ^ x[19];
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = t[64] ^ x[25];
  assign t[41] = t[65] ^ x[22];
  assign t[42] = t[66] ^ x[23];
  assign t[43] = t[67] ^ x[24];
  assign t[44] = t[68] ^ x[30];
  assign t[45] = t[69] ^ x[27];
  assign t[46] = t[70] ^ x[28];
  assign t[47] = t[71] ^ x[29];
  assign t[48] = (x[1]);
  assign t[49] = (x[1]);
  assign t[4] = t[8] & t[9];
  assign t[50] = (x[1]);
  assign t[51] = (x[1]);
  assign t[52] = (x[6]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[6]);
  assign t[56] = (x[11]);
  assign t[57] = (x[11]);
  assign t[58] = (x[11]);
  assign t[59] = (x[11]);
  assign t[5] = ~(t[10] | t[11]);
  assign t[60] = (x[16]);
  assign t[61] = (x[16]);
  assign t[62] = (x[16]);
  assign t[63] = (x[16]);
  assign t[64] = (x[21]);
  assign t[65] = (x[21]);
  assign t[66] = (x[21]);
  assign t[67] = (x[21]);
  assign t[68] = (x[26]);
  assign t[69] = (x[26]);
  assign t[6] = (t[12]);
  assign t[70] = (x[26]);
  assign t[71] = (x[26]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind12(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind13(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind14(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind15(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind16(x, y);
 input [30:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[5];
  assign t[13] = t[19] ^ x[10];
  assign t[14] = t[20] ^ x[15];
  assign t[15] = t[21] ^ x[20];
  assign t[16] = t[22] ^ x[25];
  assign t[17] = t[23] ^ x[30];
  assign t[18] = (~t[24] & t[25] & t[26] & t[27]) | (t[24] & ~t[26] & ~t[27]) | (t[24] & ~t[25] & ~t[27]) | (t[24] & ~t[25] & ~t[26]);
  assign t[19] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[1] = t[2] & t[6];
  assign t[20] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[21] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[22] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[23] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[24] = t[48] ^ x[5];
  assign t[25] = t[49] ^ x[2];
  assign t[26] = t[50] ^ x[3];
  assign t[27] = t[51] ^ x[4];
  assign t[28] = t[52] ^ x[10];
  assign t[29] = t[53] ^ x[7];
  assign t[2] = ~(t[3] & t[7]);
  assign t[30] = t[54] ^ x[8];
  assign t[31] = t[55] ^ x[9];
  assign t[32] = t[56] ^ x[15];
  assign t[33] = t[57] ^ x[12];
  assign t[34] = t[58] ^ x[13];
  assign t[35] = t[59] ^ x[14];
  assign t[36] = t[60] ^ x[20];
  assign t[37] = t[61] ^ x[17];
  assign t[38] = t[62] ^ x[18];
  assign t[39] = t[63] ^ x[19];
  assign t[3] = ~(t[8] | t[4]);
  assign t[40] = t[64] ^ x[25];
  assign t[41] = t[65] ^ x[22];
  assign t[42] = t[66] ^ x[23];
  assign t[43] = t[67] ^ x[24];
  assign t[44] = t[68] ^ x[30];
  assign t[45] = t[69] ^ x[27];
  assign t[46] = t[70] ^ x[28];
  assign t[47] = t[71] ^ x[29];
  assign t[48] = (x[1]);
  assign t[49] = (x[1]);
  assign t[4] = ~(t[9] & t[5]);
  assign t[50] = (x[1]);
  assign t[51] = (x[1]);
  assign t[52] = (x[6]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[6]);
  assign t[56] = (x[11]);
  assign t[57] = (x[11]);
  assign t[58] = (x[11]);
  assign t[59] = (x[11]);
  assign t[5] = ~(t[10] | t[11]);
  assign t[60] = (x[16]);
  assign t[61] = (x[16]);
  assign t[62] = (x[16]);
  assign t[63] = (x[16]);
  assign t[64] = (x[21]);
  assign t[65] = (x[21]);
  assign t[66] = (x[21]);
  assign t[67] = (x[21]);
  assign t[68] = (x[26]);
  assign t[69] = (x[26]);
  assign t[6] = (t[12]);
  assign t[70] = (x[26]);
  assign t[71] = (x[26]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind17(x, y);
 input [30:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[5];
  assign t[13] = t[19] ^ x[10];
  assign t[14] = t[20] ^ x[15];
  assign t[15] = t[21] ^ x[20];
  assign t[16] = t[22] ^ x[25];
  assign t[17] = t[23] ^ x[30];
  assign t[18] = (~t[24] & t[25] & t[26] & t[27]) | (t[24] & ~t[26] & ~t[27]) | (t[24] & ~t[25] & ~t[27]) | (t[24] & ~t[25] & ~t[26]);
  assign t[19] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[1] = t[2] & t[6];
  assign t[20] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[21] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[22] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[23] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[24] = t[48] ^ x[5];
  assign t[25] = t[49] ^ x[2];
  assign t[26] = t[50] ^ x[3];
  assign t[27] = t[51] ^ x[4];
  assign t[28] = t[52] ^ x[10];
  assign t[29] = t[53] ^ x[7];
  assign t[2] = ~(t[3] & t[7]);
  assign t[30] = t[54] ^ x[8];
  assign t[31] = t[55] ^ x[9];
  assign t[32] = t[56] ^ x[15];
  assign t[33] = t[57] ^ x[12];
  assign t[34] = t[58] ^ x[13];
  assign t[35] = t[59] ^ x[14];
  assign t[36] = t[60] ^ x[20];
  assign t[37] = t[61] ^ x[17];
  assign t[38] = t[62] ^ x[18];
  assign t[39] = t[63] ^ x[19];
  assign t[3] = ~(t[8] | t[4]);
  assign t[40] = t[64] ^ x[25];
  assign t[41] = t[65] ^ x[22];
  assign t[42] = t[66] ^ x[23];
  assign t[43] = t[67] ^ x[24];
  assign t[44] = t[68] ^ x[30];
  assign t[45] = t[69] ^ x[27];
  assign t[46] = t[70] ^ x[28];
  assign t[47] = t[71] ^ x[29];
  assign t[48] = (x[1]);
  assign t[49] = (x[1]);
  assign t[4] = ~(t[9] & t[5]);
  assign t[50] = (x[1]);
  assign t[51] = (x[1]);
  assign t[52] = (x[6]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[6]);
  assign t[56] = (x[11]);
  assign t[57] = (x[11]);
  assign t[58] = (x[11]);
  assign t[59] = (x[11]);
  assign t[5] = ~(t[10] | t[11]);
  assign t[60] = (x[16]);
  assign t[61] = (x[16]);
  assign t[62] = (x[16]);
  assign t[63] = (x[16]);
  assign t[64] = (x[21]);
  assign t[65] = (x[21]);
  assign t[66] = (x[21]);
  assign t[67] = (x[21]);
  assign t[68] = (x[26]);
  assign t[69] = (x[26]);
  assign t[6] = (t[12]);
  assign t[70] = (x[26]);
  assign t[71] = (x[26]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind18(x, y);
 input [30:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[5];
  assign t[13] = t[19] ^ x[10];
  assign t[14] = t[20] ^ x[15];
  assign t[15] = t[21] ^ x[20];
  assign t[16] = t[22] ^ x[25];
  assign t[17] = t[23] ^ x[30];
  assign t[18] = (~t[24] & t[25] & t[26] & t[27]) | (t[24] & ~t[26] & ~t[27]) | (t[24] & ~t[25] & ~t[27]) | (t[24] & ~t[25] & ~t[26]);
  assign t[19] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[1] = t[2] & t[6];
  assign t[20] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[21] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[22] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[23] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[24] = t[48] ^ x[5];
  assign t[25] = t[49] ^ x[2];
  assign t[26] = t[50] ^ x[3];
  assign t[27] = t[51] ^ x[4];
  assign t[28] = t[52] ^ x[10];
  assign t[29] = t[53] ^ x[7];
  assign t[2] = ~(t[3] & t[7]);
  assign t[30] = t[54] ^ x[8];
  assign t[31] = t[55] ^ x[9];
  assign t[32] = t[56] ^ x[15];
  assign t[33] = t[57] ^ x[12];
  assign t[34] = t[58] ^ x[13];
  assign t[35] = t[59] ^ x[14];
  assign t[36] = t[60] ^ x[20];
  assign t[37] = t[61] ^ x[17];
  assign t[38] = t[62] ^ x[18];
  assign t[39] = t[63] ^ x[19];
  assign t[3] = ~(t[8] | t[4]);
  assign t[40] = t[64] ^ x[25];
  assign t[41] = t[65] ^ x[22];
  assign t[42] = t[66] ^ x[23];
  assign t[43] = t[67] ^ x[24];
  assign t[44] = t[68] ^ x[30];
  assign t[45] = t[69] ^ x[27];
  assign t[46] = t[70] ^ x[28];
  assign t[47] = t[71] ^ x[29];
  assign t[48] = (x[1]);
  assign t[49] = (x[1]);
  assign t[4] = ~(t[9] & t[5]);
  assign t[50] = (x[1]);
  assign t[51] = (x[1]);
  assign t[52] = (x[6]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[6]);
  assign t[56] = (x[11]);
  assign t[57] = (x[11]);
  assign t[58] = (x[11]);
  assign t[59] = (x[11]);
  assign t[5] = ~(t[10] | t[11]);
  assign t[60] = (x[16]);
  assign t[61] = (x[16]);
  assign t[62] = (x[16]);
  assign t[63] = (x[16]);
  assign t[64] = (x[21]);
  assign t[65] = (x[21]);
  assign t[66] = (x[21]);
  assign t[67] = (x[21]);
  assign t[68] = (x[26]);
  assign t[69] = (x[26]);
  assign t[6] = (t[12]);
  assign t[70] = (x[26]);
  assign t[71] = (x[26]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind19(x, y);
 input [30:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[5];
  assign t[13] = t[19] ^ x[10];
  assign t[14] = t[20] ^ x[15];
  assign t[15] = t[21] ^ x[20];
  assign t[16] = t[22] ^ x[25];
  assign t[17] = t[23] ^ x[30];
  assign t[18] = (~t[24] & t[25] & t[26] & t[27]) | (t[24] & ~t[26] & ~t[27]) | (t[24] & ~t[25] & ~t[27]) | (t[24] & ~t[25] & ~t[26]);
  assign t[19] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[1] = t[2] & t[6];
  assign t[20] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[21] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[22] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[23] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[24] = t[48] ^ x[5];
  assign t[25] = t[49] ^ x[2];
  assign t[26] = t[50] ^ x[3];
  assign t[27] = t[51] ^ x[4];
  assign t[28] = t[52] ^ x[10];
  assign t[29] = t[53] ^ x[7];
  assign t[2] = ~(t[3] & t[7]);
  assign t[30] = t[54] ^ x[8];
  assign t[31] = t[55] ^ x[9];
  assign t[32] = t[56] ^ x[15];
  assign t[33] = t[57] ^ x[12];
  assign t[34] = t[58] ^ x[13];
  assign t[35] = t[59] ^ x[14];
  assign t[36] = t[60] ^ x[20];
  assign t[37] = t[61] ^ x[17];
  assign t[38] = t[62] ^ x[18];
  assign t[39] = t[63] ^ x[19];
  assign t[3] = ~(t[8] | t[4]);
  assign t[40] = t[64] ^ x[25];
  assign t[41] = t[65] ^ x[22];
  assign t[42] = t[66] ^ x[23];
  assign t[43] = t[67] ^ x[24];
  assign t[44] = t[68] ^ x[30];
  assign t[45] = t[69] ^ x[27];
  assign t[46] = t[70] ^ x[28];
  assign t[47] = t[71] ^ x[29];
  assign t[48] = (x[1]);
  assign t[49] = (x[1]);
  assign t[4] = ~(t[9] & t[5]);
  assign t[50] = (x[1]);
  assign t[51] = (x[1]);
  assign t[52] = (x[6]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[6]);
  assign t[56] = (x[11]);
  assign t[57] = (x[11]);
  assign t[58] = (x[11]);
  assign t[59] = (x[11]);
  assign t[5] = ~(t[10] | t[11]);
  assign t[60] = (x[16]);
  assign t[61] = (x[16]);
  assign t[62] = (x[16]);
  assign t[63] = (x[16]);
  assign t[64] = (x[21]);
  assign t[65] = (x[21]);
  assign t[66] = (x[21]);
  assign t[67] = (x[21]);
  assign t[68] = (x[26]);
  assign t[69] = (x[26]);
  assign t[6] = (t[12]);
  assign t[70] = (x[26]);
  assign t[71] = (x[26]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind20(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind21(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind22(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind23(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind24(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind25(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind26(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind27(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind28(x, y);
 input [30:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[5];
  assign t[13] = t[19] ^ x[10];
  assign t[14] = t[20] ^ x[15];
  assign t[15] = t[21] ^ x[20];
  assign t[16] = t[22] ^ x[25];
  assign t[17] = t[23] ^ x[30];
  assign t[18] = (~t[24] & t[25] & t[26] & t[27]) | (t[24] & ~t[26] & ~t[27]) | (t[24] & ~t[25] & ~t[27]) | (t[24] & ~t[25] & ~t[26]);
  assign t[19] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[1] = t[6] | t[2];
  assign t[20] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[21] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[22] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[23] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[24] = t[48] ^ x[5];
  assign t[25] = t[49] ^ x[2];
  assign t[26] = t[50] ^ x[3];
  assign t[27] = t[51] ^ x[4];
  assign t[28] = t[52] ^ x[10];
  assign t[29] = t[53] ^ x[7];
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = t[54] ^ x[8];
  assign t[31] = t[55] ^ x[9];
  assign t[32] = t[56] ^ x[15];
  assign t[33] = t[57] ^ x[12];
  assign t[34] = t[58] ^ x[13];
  assign t[35] = t[59] ^ x[14];
  assign t[36] = t[60] ^ x[20];
  assign t[37] = t[61] ^ x[17];
  assign t[38] = t[62] ^ x[18];
  assign t[39] = t[63] ^ x[19];
  assign t[3] = ~(t[8] & t[4]);
  assign t[40] = t[64] ^ x[25];
  assign t[41] = t[65] ^ x[22];
  assign t[42] = t[66] ^ x[23];
  assign t[43] = t[67] ^ x[24];
  assign t[44] = t[68] ^ x[30];
  assign t[45] = t[69] ^ x[27];
  assign t[46] = t[70] ^ x[28];
  assign t[47] = t[71] ^ x[29];
  assign t[48] = (x[1]);
  assign t[49] = (x[1]);
  assign t[4] = ~(t[9] | t[5]);
  assign t[50] = (x[1]);
  assign t[51] = (x[1]);
  assign t[52] = (x[6]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[6]);
  assign t[56] = (x[11]);
  assign t[57] = (x[11]);
  assign t[58] = (x[11]);
  assign t[59] = (x[11]);
  assign t[5] = ~(t[10] & t[11]);
  assign t[60] = (x[16]);
  assign t[61] = (x[16]);
  assign t[62] = (x[16]);
  assign t[63] = (x[16]);
  assign t[64] = (x[21]);
  assign t[65] = (x[21]);
  assign t[66] = (x[21]);
  assign t[67] = (x[21]);
  assign t[68] = (x[26]);
  assign t[69] = (x[26]);
  assign t[6] = (t[12]);
  assign t[70] = (x[26]);
  assign t[71] = (x[26]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind29(x, y);
 input [30:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[5];
  assign t[13] = t[19] ^ x[10];
  assign t[14] = t[20] ^ x[15];
  assign t[15] = t[21] ^ x[20];
  assign t[16] = t[22] ^ x[25];
  assign t[17] = t[23] ^ x[30];
  assign t[18] = (~t[24] & t[25] & t[26] & t[27]) | (t[24] & ~t[26] & ~t[27]) | (t[24] & ~t[25] & ~t[27]) | (t[24] & ~t[25] & ~t[26]);
  assign t[19] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[1] = t[6] | t[2];
  assign t[20] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[21] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[22] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[23] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[24] = t[48] ^ x[5];
  assign t[25] = t[49] ^ x[2];
  assign t[26] = t[50] ^ x[3];
  assign t[27] = t[51] ^ x[4];
  assign t[28] = t[52] ^ x[10];
  assign t[29] = t[53] ^ x[7];
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = t[54] ^ x[8];
  assign t[31] = t[55] ^ x[9];
  assign t[32] = t[56] ^ x[15];
  assign t[33] = t[57] ^ x[12];
  assign t[34] = t[58] ^ x[13];
  assign t[35] = t[59] ^ x[14];
  assign t[36] = t[60] ^ x[20];
  assign t[37] = t[61] ^ x[17];
  assign t[38] = t[62] ^ x[18];
  assign t[39] = t[63] ^ x[19];
  assign t[3] = ~(t[8] & t[4]);
  assign t[40] = t[64] ^ x[25];
  assign t[41] = t[65] ^ x[22];
  assign t[42] = t[66] ^ x[23];
  assign t[43] = t[67] ^ x[24];
  assign t[44] = t[68] ^ x[30];
  assign t[45] = t[69] ^ x[27];
  assign t[46] = t[70] ^ x[28];
  assign t[47] = t[71] ^ x[29];
  assign t[48] = (x[1]);
  assign t[49] = (x[1]);
  assign t[4] = ~(t[9] | t[5]);
  assign t[50] = (x[1]);
  assign t[51] = (x[1]);
  assign t[52] = (x[6]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[6]);
  assign t[56] = (x[11]);
  assign t[57] = (x[11]);
  assign t[58] = (x[11]);
  assign t[59] = (x[11]);
  assign t[5] = ~(t[10] & t[11]);
  assign t[60] = (x[16]);
  assign t[61] = (x[16]);
  assign t[62] = (x[16]);
  assign t[63] = (x[16]);
  assign t[64] = (x[21]);
  assign t[65] = (x[21]);
  assign t[66] = (x[21]);
  assign t[67] = (x[21]);
  assign t[68] = (x[26]);
  assign t[69] = (x[26]);
  assign t[6] = (t[12]);
  assign t[70] = (x[26]);
  assign t[71] = (x[26]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind30(x, y);
 input [30:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[5];
  assign t[13] = t[19] ^ x[10];
  assign t[14] = t[20] ^ x[15];
  assign t[15] = t[21] ^ x[20];
  assign t[16] = t[22] ^ x[25];
  assign t[17] = t[23] ^ x[30];
  assign t[18] = (~t[24] & t[25] & t[26] & t[27]) | (t[24] & ~t[26] & ~t[27]) | (t[24] & ~t[25] & ~t[27]) | (t[24] & ~t[25] & ~t[26]);
  assign t[19] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[1] = t[6] | t[2];
  assign t[20] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[21] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[22] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[23] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[24] = t[48] ^ x[5];
  assign t[25] = t[49] ^ x[2];
  assign t[26] = t[50] ^ x[3];
  assign t[27] = t[51] ^ x[4];
  assign t[28] = t[52] ^ x[10];
  assign t[29] = t[53] ^ x[7];
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = t[54] ^ x[8];
  assign t[31] = t[55] ^ x[9];
  assign t[32] = t[56] ^ x[15];
  assign t[33] = t[57] ^ x[12];
  assign t[34] = t[58] ^ x[13];
  assign t[35] = t[59] ^ x[14];
  assign t[36] = t[60] ^ x[20];
  assign t[37] = t[61] ^ x[17];
  assign t[38] = t[62] ^ x[18];
  assign t[39] = t[63] ^ x[19];
  assign t[3] = ~(t[8] & t[4]);
  assign t[40] = t[64] ^ x[25];
  assign t[41] = t[65] ^ x[22];
  assign t[42] = t[66] ^ x[23];
  assign t[43] = t[67] ^ x[24];
  assign t[44] = t[68] ^ x[30];
  assign t[45] = t[69] ^ x[27];
  assign t[46] = t[70] ^ x[28];
  assign t[47] = t[71] ^ x[29];
  assign t[48] = (x[1]);
  assign t[49] = (x[1]);
  assign t[4] = ~(t[9] | t[5]);
  assign t[50] = (x[1]);
  assign t[51] = (x[1]);
  assign t[52] = (x[6]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[6]);
  assign t[56] = (x[11]);
  assign t[57] = (x[11]);
  assign t[58] = (x[11]);
  assign t[59] = (x[11]);
  assign t[5] = ~(t[10] & t[11]);
  assign t[60] = (x[16]);
  assign t[61] = (x[16]);
  assign t[62] = (x[16]);
  assign t[63] = (x[16]);
  assign t[64] = (x[21]);
  assign t[65] = (x[21]);
  assign t[66] = (x[21]);
  assign t[67] = (x[21]);
  assign t[68] = (x[26]);
  assign t[69] = (x[26]);
  assign t[6] = (t[12]);
  assign t[70] = (x[26]);
  assign t[71] = (x[26]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind31(x, y);
 input [30:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[5];
  assign t[13] = t[19] ^ x[10];
  assign t[14] = t[20] ^ x[15];
  assign t[15] = t[21] ^ x[20];
  assign t[16] = t[22] ^ x[25];
  assign t[17] = t[23] ^ x[30];
  assign t[18] = (~t[24] & t[25] & t[26] & t[27]) | (t[24] & ~t[26] & ~t[27]) | (t[24] & ~t[25] & ~t[27]) | (t[24] & ~t[25] & ~t[26]);
  assign t[19] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[1] = t[6] | t[2];
  assign t[20] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[21] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[22] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[23] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[24] = t[48] ^ x[5];
  assign t[25] = t[49] ^ x[2];
  assign t[26] = t[50] ^ x[3];
  assign t[27] = t[51] ^ x[4];
  assign t[28] = t[52] ^ x[10];
  assign t[29] = t[53] ^ x[7];
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = t[54] ^ x[8];
  assign t[31] = t[55] ^ x[9];
  assign t[32] = t[56] ^ x[15];
  assign t[33] = t[57] ^ x[12];
  assign t[34] = t[58] ^ x[13];
  assign t[35] = t[59] ^ x[14];
  assign t[36] = t[60] ^ x[20];
  assign t[37] = t[61] ^ x[17];
  assign t[38] = t[62] ^ x[18];
  assign t[39] = t[63] ^ x[19];
  assign t[3] = ~(t[8] & t[4]);
  assign t[40] = t[64] ^ x[25];
  assign t[41] = t[65] ^ x[22];
  assign t[42] = t[66] ^ x[23];
  assign t[43] = t[67] ^ x[24];
  assign t[44] = t[68] ^ x[30];
  assign t[45] = t[69] ^ x[27];
  assign t[46] = t[70] ^ x[28];
  assign t[47] = t[71] ^ x[29];
  assign t[48] = (x[1]);
  assign t[49] = (x[1]);
  assign t[4] = ~(t[9] | t[5]);
  assign t[50] = (x[1]);
  assign t[51] = (x[1]);
  assign t[52] = (x[6]);
  assign t[53] = (x[6]);
  assign t[54] = (x[6]);
  assign t[55] = (x[6]);
  assign t[56] = (x[11]);
  assign t[57] = (x[11]);
  assign t[58] = (x[11]);
  assign t[59] = (x[11]);
  assign t[5] = ~(t[10] & t[11]);
  assign t[60] = (x[16]);
  assign t[61] = (x[16]);
  assign t[62] = (x[16]);
  assign t[63] = (x[16]);
  assign t[64] = (x[21]);
  assign t[65] = (x[21]);
  assign t[66] = (x[21]);
  assign t[67] = (x[21]);
  assign t[68] = (x[26]);
  assign t[69] = (x[26]);
  assign t[6] = (t[12]);
  assign t[70] = (x[26]);
  assign t[71] = (x[26]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind32(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind33(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind34(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind35(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind36(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[38] ^ t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind37(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[38] ^ t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind38(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[38] ^ t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind39(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[38] ^ t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind40(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind41(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind42(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind43(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind44(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind45(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind46(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind47(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind48(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind49(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind50(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind51(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind52(x, y);
 input [46:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[136] ^ x[45];
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[2]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[7]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[17];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[12]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[17]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[18] & t[19];
  assign t[120] = (x[22]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[27]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[32]);
  assign t[129] = (x[37]);
  assign t[12] = t[20] ^ t[11];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[37]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[136] = (x[42]);
  assign t[13] = t[39] ^ t[18];
  assign t[14] = t[21] ^ t[22];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[40] ^ t[41];
  assign t[17] = t[18] & t[25];
  assign t[18] = ~(t[41]);
  assign t[19] = ~(t[39] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[39] & t[26];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[42] ^ t[29];
  assign t[25] = t[39] ^ t[32];
  assign t[26] = t[33] ^ t[17];
  assign t[27] = t[43] ^ t[44];
  assign t[28] = t[29] & t[34];
  assign t[29] = ~(t[44]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[42] ^ t[29]);
  assign t[31] = t[42] & t[35];
  assign t[32] = t[41] ^ t[45];
  assign t[33] = t[39] ^ t[16];
  assign t[34] = t[42] ^ t[36];
  assign t[35] = t[37] ^ t[28];
  assign t[36] = t[44] ^ t[46];
  assign t[37] = t[42] ^ t[27];
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = (t[55]);
  assign t[47] = t[56] ^ x[6];
  assign t[48] = t[57] ^ x[11];
  assign t[49] = t[58] ^ x[16];
  assign t[4] = ~(t[6] ^ t[38]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[26];
  assign t[52] = t[61] ^ x[31];
  assign t[53] = t[62] ^ x[36];
  assign t[54] = t[63] ^ x[41];
  assign t[55] = t[64] ^ x[46];
  assign t[56] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[57] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[58] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[59] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[60] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[61] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[62] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[63] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[64] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[65] = t[101] ^ x[6];
  assign t[66] = t[102] ^ x[3];
  assign t[67] = t[103] ^ x[4];
  assign t[68] = t[104] ^ x[5];
  assign t[69] = t[105] ^ x[11];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[8];
  assign t[71] = t[107] ^ x[9];
  assign t[72] = t[108] ^ x[10];
  assign t[73] = t[109] ^ x[16];
  assign t[74] = t[110] ^ x[13];
  assign t[75] = t[111] ^ x[14];
  assign t[76] = t[112] ^ x[15];
  assign t[77] = t[113] ^ x[21];
  assign t[78] = t[114] ^ x[18];
  assign t[79] = t[115] ^ x[19];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[20];
  assign t[81] = t[117] ^ x[26];
  assign t[82] = t[118] ^ x[23];
  assign t[83] = t[119] ^ x[24];
  assign t[84] = t[120] ^ x[25];
  assign t[85] = t[121] ^ x[31];
  assign t[86] = t[122] ^ x[28];
  assign t[87] = t[123] ^ x[29];
  assign t[88] = t[124] ^ x[30];
  assign t[89] = t[125] ^ x[36];
  assign t[8] = t[12] ^ t[13];
  assign t[90] = t[126] ^ x[33];
  assign t[91] = t[127] ^ x[34];
  assign t[92] = t[128] ^ x[35];
  assign t[93] = t[129] ^ x[41];
  assign t[94] = t[130] ^ x[38];
  assign t[95] = t[131] ^ x[39];
  assign t[96] = t[132] ^ x[40];
  assign t[97] = t[133] ^ x[46];
  assign t[98] = t[134] ^ x[43];
  assign t[99] = t[135] ^ x[44];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = (t[0]);
endmodule

module R2ind53(x, y);
 input [46:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[136] ^ x[45];
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[2]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[7]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[17];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[12]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[17]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[18] & t[19];
  assign t[120] = (x[22]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[27]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[32]);
  assign t[129] = (x[37]);
  assign t[12] = t[20] ^ t[11];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[37]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[136] = (x[42]);
  assign t[13] = t[39] ^ t[18];
  assign t[14] = t[21] ^ t[22];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[40] ^ t[41];
  assign t[17] = t[18] & t[25];
  assign t[18] = ~(t[41]);
  assign t[19] = ~(t[39] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[39] & t[26];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[42] ^ t[29];
  assign t[25] = t[39] ^ t[32];
  assign t[26] = t[33] ^ t[17];
  assign t[27] = t[43] ^ t[44];
  assign t[28] = t[29] & t[34];
  assign t[29] = ~(t[44]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[42] ^ t[29]);
  assign t[31] = t[42] & t[35];
  assign t[32] = t[41] ^ t[45];
  assign t[33] = t[39] ^ t[16];
  assign t[34] = t[42] ^ t[36];
  assign t[35] = t[37] ^ t[28];
  assign t[36] = t[44] ^ t[46];
  assign t[37] = t[42] ^ t[27];
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = (t[55]);
  assign t[47] = t[56] ^ x[6];
  assign t[48] = t[57] ^ x[11];
  assign t[49] = t[58] ^ x[16];
  assign t[4] = ~(t[6] ^ t[38]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[26];
  assign t[52] = t[61] ^ x[31];
  assign t[53] = t[62] ^ x[36];
  assign t[54] = t[63] ^ x[41];
  assign t[55] = t[64] ^ x[46];
  assign t[56] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[57] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[58] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[59] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[60] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[61] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[62] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[63] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[64] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[65] = t[101] ^ x[6];
  assign t[66] = t[102] ^ x[3];
  assign t[67] = t[103] ^ x[4];
  assign t[68] = t[104] ^ x[5];
  assign t[69] = t[105] ^ x[11];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[8];
  assign t[71] = t[107] ^ x[9];
  assign t[72] = t[108] ^ x[10];
  assign t[73] = t[109] ^ x[16];
  assign t[74] = t[110] ^ x[13];
  assign t[75] = t[111] ^ x[14];
  assign t[76] = t[112] ^ x[15];
  assign t[77] = t[113] ^ x[21];
  assign t[78] = t[114] ^ x[18];
  assign t[79] = t[115] ^ x[19];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[20];
  assign t[81] = t[117] ^ x[26];
  assign t[82] = t[118] ^ x[23];
  assign t[83] = t[119] ^ x[24];
  assign t[84] = t[120] ^ x[25];
  assign t[85] = t[121] ^ x[31];
  assign t[86] = t[122] ^ x[28];
  assign t[87] = t[123] ^ x[29];
  assign t[88] = t[124] ^ x[30];
  assign t[89] = t[125] ^ x[36];
  assign t[8] = t[12] ^ t[13];
  assign t[90] = t[126] ^ x[33];
  assign t[91] = t[127] ^ x[34];
  assign t[92] = t[128] ^ x[35];
  assign t[93] = t[129] ^ x[41];
  assign t[94] = t[130] ^ x[38];
  assign t[95] = t[131] ^ x[39];
  assign t[96] = t[132] ^ x[40];
  assign t[97] = t[133] ^ x[46];
  assign t[98] = t[134] ^ x[43];
  assign t[99] = t[135] ^ x[44];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = (t[0]);
endmodule

module R2ind54(x, y);
 input [46:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[136] ^ x[45];
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[2]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[7]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[17];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[12]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[17]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[18] & t[19];
  assign t[120] = (x[22]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[27]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[32]);
  assign t[129] = (x[37]);
  assign t[12] = t[20] ^ t[11];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[37]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[136] = (x[42]);
  assign t[13] = t[39] ^ t[18];
  assign t[14] = t[21] ^ t[22];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[40] ^ t[41];
  assign t[17] = t[18] & t[25];
  assign t[18] = ~(t[41]);
  assign t[19] = ~(t[39] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[39] & t[26];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[42] ^ t[29];
  assign t[25] = t[39] ^ t[32];
  assign t[26] = t[33] ^ t[17];
  assign t[27] = t[43] ^ t[44];
  assign t[28] = t[29] & t[34];
  assign t[29] = ~(t[44]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[42] ^ t[29]);
  assign t[31] = t[42] & t[35];
  assign t[32] = t[41] ^ t[45];
  assign t[33] = t[39] ^ t[16];
  assign t[34] = t[42] ^ t[36];
  assign t[35] = t[37] ^ t[28];
  assign t[36] = t[44] ^ t[46];
  assign t[37] = t[42] ^ t[27];
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = (t[55]);
  assign t[47] = t[56] ^ x[6];
  assign t[48] = t[57] ^ x[11];
  assign t[49] = t[58] ^ x[16];
  assign t[4] = ~(t[6] ^ t[38]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[26];
  assign t[52] = t[61] ^ x[31];
  assign t[53] = t[62] ^ x[36];
  assign t[54] = t[63] ^ x[41];
  assign t[55] = t[64] ^ x[46];
  assign t[56] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[57] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[58] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[59] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[60] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[61] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[62] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[63] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[64] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[65] = t[101] ^ x[6];
  assign t[66] = t[102] ^ x[3];
  assign t[67] = t[103] ^ x[4];
  assign t[68] = t[104] ^ x[5];
  assign t[69] = t[105] ^ x[11];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[8];
  assign t[71] = t[107] ^ x[9];
  assign t[72] = t[108] ^ x[10];
  assign t[73] = t[109] ^ x[16];
  assign t[74] = t[110] ^ x[13];
  assign t[75] = t[111] ^ x[14];
  assign t[76] = t[112] ^ x[15];
  assign t[77] = t[113] ^ x[21];
  assign t[78] = t[114] ^ x[18];
  assign t[79] = t[115] ^ x[19];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[20];
  assign t[81] = t[117] ^ x[26];
  assign t[82] = t[118] ^ x[23];
  assign t[83] = t[119] ^ x[24];
  assign t[84] = t[120] ^ x[25];
  assign t[85] = t[121] ^ x[31];
  assign t[86] = t[122] ^ x[28];
  assign t[87] = t[123] ^ x[29];
  assign t[88] = t[124] ^ x[30];
  assign t[89] = t[125] ^ x[36];
  assign t[8] = t[12] ^ t[13];
  assign t[90] = t[126] ^ x[33];
  assign t[91] = t[127] ^ x[34];
  assign t[92] = t[128] ^ x[35];
  assign t[93] = t[129] ^ x[41];
  assign t[94] = t[130] ^ x[38];
  assign t[95] = t[131] ^ x[39];
  assign t[96] = t[132] ^ x[40];
  assign t[97] = t[133] ^ x[46];
  assign t[98] = t[134] ^ x[43];
  assign t[99] = t[135] ^ x[44];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = (t[0]);
endmodule

module R2ind55(x, y);
 input [46:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[136] ^ x[45];
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[2]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[7]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[17];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[12]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[17]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[18] & t[19];
  assign t[120] = (x[22]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[27]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[32]);
  assign t[129] = (x[37]);
  assign t[12] = t[20] ^ t[11];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[37]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[136] = (x[42]);
  assign t[13] = t[39] ^ t[18];
  assign t[14] = t[21] ^ t[22];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[40] ^ t[41];
  assign t[17] = t[18] & t[25];
  assign t[18] = ~(t[41]);
  assign t[19] = ~(t[39] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[39] & t[26];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[42] ^ t[29];
  assign t[25] = t[39] ^ t[32];
  assign t[26] = t[33] ^ t[17];
  assign t[27] = t[43] ^ t[44];
  assign t[28] = t[29] & t[34];
  assign t[29] = ~(t[44]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[42] ^ t[29]);
  assign t[31] = t[42] & t[35];
  assign t[32] = t[41] ^ t[45];
  assign t[33] = t[39] ^ t[16];
  assign t[34] = t[42] ^ t[36];
  assign t[35] = t[37] ^ t[28];
  assign t[36] = t[44] ^ t[46];
  assign t[37] = t[42] ^ t[27];
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = (t[55]);
  assign t[47] = t[56] ^ x[6];
  assign t[48] = t[57] ^ x[11];
  assign t[49] = t[58] ^ x[16];
  assign t[4] = ~(t[6] ^ t[38]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[26];
  assign t[52] = t[61] ^ x[31];
  assign t[53] = t[62] ^ x[36];
  assign t[54] = t[63] ^ x[41];
  assign t[55] = t[64] ^ x[46];
  assign t[56] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[57] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[58] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[59] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[60] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[61] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[62] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[63] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[64] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[65] = t[101] ^ x[6];
  assign t[66] = t[102] ^ x[3];
  assign t[67] = t[103] ^ x[4];
  assign t[68] = t[104] ^ x[5];
  assign t[69] = t[105] ^ x[11];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[8];
  assign t[71] = t[107] ^ x[9];
  assign t[72] = t[108] ^ x[10];
  assign t[73] = t[109] ^ x[16];
  assign t[74] = t[110] ^ x[13];
  assign t[75] = t[111] ^ x[14];
  assign t[76] = t[112] ^ x[15];
  assign t[77] = t[113] ^ x[21];
  assign t[78] = t[114] ^ x[18];
  assign t[79] = t[115] ^ x[19];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[20];
  assign t[81] = t[117] ^ x[26];
  assign t[82] = t[118] ^ x[23];
  assign t[83] = t[119] ^ x[24];
  assign t[84] = t[120] ^ x[25];
  assign t[85] = t[121] ^ x[31];
  assign t[86] = t[122] ^ x[28];
  assign t[87] = t[123] ^ x[29];
  assign t[88] = t[124] ^ x[30];
  assign t[89] = t[125] ^ x[36];
  assign t[8] = t[12] ^ t[13];
  assign t[90] = t[126] ^ x[33];
  assign t[91] = t[127] ^ x[34];
  assign t[92] = t[128] ^ x[35];
  assign t[93] = t[129] ^ x[41];
  assign t[94] = t[130] ^ x[38];
  assign t[95] = t[131] ^ x[39];
  assign t[96] = t[132] ^ x[40];
  assign t[97] = t[133] ^ x[46];
  assign t[98] = t[134] ^ x[43];
  assign t[99] = t[135] ^ x[44];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = (t[0]);
endmodule

module R2ind56(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind57(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind58(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind59(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind60(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind61(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind62(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind63(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind64(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind65(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind66(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind67(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind68(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[38] ^ t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind69(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[38] ^ t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind70(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[38] ^ t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind71(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[38] ^ t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind72(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind73(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind74(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind75(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind76(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind77(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind78(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind79(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind80(x, y);
 input [51:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ^ x[40];
  assign t[101] = t[141] ^ x[46];
  assign t[102] = t[142] ^ x[43];
  assign t[103] = t[143] ^ x[44];
  assign t[104] = t[144] ^ x[45];
  assign t[105] = t[145] ^ x[51];
  assign t[106] = t[146] ^ x[48];
  assign t[107] = t[147] ^ x[49];
  assign t[108] = t[148] ^ x[50];
  assign t[109] = (x[2]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[2]);
  assign t[111] = (x[2]);
  assign t[112] = (x[2]);
  assign t[113] = (x[7]);
  assign t[114] = (x[7]);
  assign t[115] = (x[7]);
  assign t[116] = (x[7]);
  assign t[117] = (x[12]);
  assign t[118] = (x[12]);
  assign t[119] = (x[12]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[12]);
  assign t[121] = (x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[17]);
  assign t[124] = (x[17]);
  assign t[125] = (x[22]);
  assign t[126] = (x[22]);
  assign t[127] = (x[22]);
  assign t[128] = (x[22]);
  assign t[129] = (x[27]);
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[130] = (x[27]);
  assign t[131] = (x[27]);
  assign t[132] = (x[27]);
  assign t[133] = (x[32]);
  assign t[134] = (x[32]);
  assign t[135] = (x[32]);
  assign t[136] = (x[32]);
  assign t[137] = (x[37]);
  assign t[138] = (x[37]);
  assign t[139] = (x[37]);
  assign t[13] = t[19] ^ t[20];
  assign t[140] = (x[37]);
  assign t[141] = (x[42]);
  assign t[142] = (x[42]);
  assign t[143] = (x[42]);
  assign t[144] = (x[42]);
  assign t[145] = (x[47]);
  assign t[146] = (x[47]);
  assign t[147] = (x[47]);
  assign t[148] = (x[47]);
  assign t[14] = ~(t[42]);
  assign t[15] = ~(t[40] ^ t[14]);
  assign t[16] = t[43] ^ t[42];
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[18] = ~t[22];
  assign t[19] = t[40] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[40] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[42] ^ t[44];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[45] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[45] ^ t[31]);
  assign t[33] = t[47] ^ t[46];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[45] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[45] ^ t[38];
  assign t[38] = t[46] ^ t[48];
  assign t[39] = (t[49]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[6];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[11];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[21];
  assign t[53] = t[63] ^ x[26];
  assign t[54] = t[64] ^ x[31];
  assign t[55] = t[65] ^ x[36];
  assign t[56] = t[66] ^ x[41];
  assign t[57] = t[67] ^ x[46];
  assign t[58] = t[68] ^ x[51];
  assign t[59] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[61] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[62] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[63] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[64] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[65] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[66] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[67] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[68] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[69] = t[109] ^ x[6];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[110] ^ x[3];
  assign t[71] = t[111] ^ x[4];
  assign t[72] = t[112] ^ x[5];
  assign t[73] = t[113] ^ x[11];
  assign t[74] = t[114] ^ x[8];
  assign t[75] = t[115] ^ x[9];
  assign t[76] = t[116] ^ x[10];
  assign t[77] = t[117] ^ x[16];
  assign t[78] = t[118] ^ x[13];
  assign t[79] = t[119] ^ x[14];
  assign t[7] = ~t[12];
  assign t[80] = t[120] ^ x[15];
  assign t[81] = t[121] ^ x[21];
  assign t[82] = t[122] ^ x[18];
  assign t[83] = t[123] ^ x[19];
  assign t[84] = t[124] ^ x[20];
  assign t[85] = t[125] ^ x[26];
  assign t[86] = t[126] ^ x[23];
  assign t[87] = t[127] ^ x[24];
  assign t[88] = t[128] ^ x[25];
  assign t[89] = t[129] ^ x[31];
  assign t[8] = t[40] & t[13];
  assign t[90] = t[130] ^ x[28];
  assign t[91] = t[131] ^ x[29];
  assign t[92] = t[132] ^ x[30];
  assign t[93] = t[133] ^ x[36];
  assign t[94] = t[134] ^ x[33];
  assign t[95] = t[135] ^ x[34];
  assign t[96] = t[136] ^ x[35];
  assign t[97] = t[137] ^ x[41];
  assign t[98] = t[138] ^ x[38];
  assign t[99] = t[139] ^ x[39];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind81(x, y);
 input [51:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ^ x[40];
  assign t[101] = t[141] ^ x[46];
  assign t[102] = t[142] ^ x[43];
  assign t[103] = t[143] ^ x[44];
  assign t[104] = t[144] ^ x[45];
  assign t[105] = t[145] ^ x[51];
  assign t[106] = t[146] ^ x[48];
  assign t[107] = t[147] ^ x[49];
  assign t[108] = t[148] ^ x[50];
  assign t[109] = (x[2]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[2]);
  assign t[111] = (x[2]);
  assign t[112] = (x[2]);
  assign t[113] = (x[7]);
  assign t[114] = (x[7]);
  assign t[115] = (x[7]);
  assign t[116] = (x[7]);
  assign t[117] = (x[12]);
  assign t[118] = (x[12]);
  assign t[119] = (x[12]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[12]);
  assign t[121] = (x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[17]);
  assign t[124] = (x[17]);
  assign t[125] = (x[22]);
  assign t[126] = (x[22]);
  assign t[127] = (x[22]);
  assign t[128] = (x[22]);
  assign t[129] = (x[27]);
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[130] = (x[27]);
  assign t[131] = (x[27]);
  assign t[132] = (x[27]);
  assign t[133] = (x[32]);
  assign t[134] = (x[32]);
  assign t[135] = (x[32]);
  assign t[136] = (x[32]);
  assign t[137] = (x[37]);
  assign t[138] = (x[37]);
  assign t[139] = (x[37]);
  assign t[13] = t[19] ^ t[20];
  assign t[140] = (x[37]);
  assign t[141] = (x[42]);
  assign t[142] = (x[42]);
  assign t[143] = (x[42]);
  assign t[144] = (x[42]);
  assign t[145] = (x[47]);
  assign t[146] = (x[47]);
  assign t[147] = (x[47]);
  assign t[148] = (x[47]);
  assign t[14] = ~(t[42]);
  assign t[15] = ~(t[40] ^ t[14]);
  assign t[16] = t[43] ^ t[42];
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[18] = ~t[22];
  assign t[19] = t[40] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[40] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[42] ^ t[44];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[45] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[45] ^ t[31]);
  assign t[33] = t[47] ^ t[46];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[45] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[45] ^ t[38];
  assign t[38] = t[46] ^ t[48];
  assign t[39] = (t[49]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[6];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[11];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[21];
  assign t[53] = t[63] ^ x[26];
  assign t[54] = t[64] ^ x[31];
  assign t[55] = t[65] ^ x[36];
  assign t[56] = t[66] ^ x[41];
  assign t[57] = t[67] ^ x[46];
  assign t[58] = t[68] ^ x[51];
  assign t[59] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[61] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[62] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[63] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[64] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[65] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[66] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[67] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[68] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[69] = t[109] ^ x[6];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[110] ^ x[3];
  assign t[71] = t[111] ^ x[4];
  assign t[72] = t[112] ^ x[5];
  assign t[73] = t[113] ^ x[11];
  assign t[74] = t[114] ^ x[8];
  assign t[75] = t[115] ^ x[9];
  assign t[76] = t[116] ^ x[10];
  assign t[77] = t[117] ^ x[16];
  assign t[78] = t[118] ^ x[13];
  assign t[79] = t[119] ^ x[14];
  assign t[7] = ~t[12];
  assign t[80] = t[120] ^ x[15];
  assign t[81] = t[121] ^ x[21];
  assign t[82] = t[122] ^ x[18];
  assign t[83] = t[123] ^ x[19];
  assign t[84] = t[124] ^ x[20];
  assign t[85] = t[125] ^ x[26];
  assign t[86] = t[126] ^ x[23];
  assign t[87] = t[127] ^ x[24];
  assign t[88] = t[128] ^ x[25];
  assign t[89] = t[129] ^ x[31];
  assign t[8] = t[40] & t[13];
  assign t[90] = t[130] ^ x[28];
  assign t[91] = t[131] ^ x[29];
  assign t[92] = t[132] ^ x[30];
  assign t[93] = t[133] ^ x[36];
  assign t[94] = t[134] ^ x[33];
  assign t[95] = t[135] ^ x[34];
  assign t[96] = t[136] ^ x[35];
  assign t[97] = t[137] ^ x[41];
  assign t[98] = t[138] ^ x[38];
  assign t[99] = t[139] ^ x[39];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind82(x, y);
 input [51:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ^ x[40];
  assign t[101] = t[141] ^ x[46];
  assign t[102] = t[142] ^ x[43];
  assign t[103] = t[143] ^ x[44];
  assign t[104] = t[144] ^ x[45];
  assign t[105] = t[145] ^ x[51];
  assign t[106] = t[146] ^ x[48];
  assign t[107] = t[147] ^ x[49];
  assign t[108] = t[148] ^ x[50];
  assign t[109] = (x[2]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[2]);
  assign t[111] = (x[2]);
  assign t[112] = (x[2]);
  assign t[113] = (x[7]);
  assign t[114] = (x[7]);
  assign t[115] = (x[7]);
  assign t[116] = (x[7]);
  assign t[117] = (x[12]);
  assign t[118] = (x[12]);
  assign t[119] = (x[12]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[12]);
  assign t[121] = (x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[17]);
  assign t[124] = (x[17]);
  assign t[125] = (x[22]);
  assign t[126] = (x[22]);
  assign t[127] = (x[22]);
  assign t[128] = (x[22]);
  assign t[129] = (x[27]);
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[130] = (x[27]);
  assign t[131] = (x[27]);
  assign t[132] = (x[27]);
  assign t[133] = (x[32]);
  assign t[134] = (x[32]);
  assign t[135] = (x[32]);
  assign t[136] = (x[32]);
  assign t[137] = (x[37]);
  assign t[138] = (x[37]);
  assign t[139] = (x[37]);
  assign t[13] = t[19] ^ t[20];
  assign t[140] = (x[37]);
  assign t[141] = (x[42]);
  assign t[142] = (x[42]);
  assign t[143] = (x[42]);
  assign t[144] = (x[42]);
  assign t[145] = (x[47]);
  assign t[146] = (x[47]);
  assign t[147] = (x[47]);
  assign t[148] = (x[47]);
  assign t[14] = ~(t[42]);
  assign t[15] = ~(t[40] ^ t[14]);
  assign t[16] = t[43] ^ t[42];
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[18] = ~t[22];
  assign t[19] = t[40] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[40] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[42] ^ t[44];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[45] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[45] ^ t[31]);
  assign t[33] = t[47] ^ t[46];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[45] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[45] ^ t[38];
  assign t[38] = t[46] ^ t[48];
  assign t[39] = (t[49]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[6];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[11];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[21];
  assign t[53] = t[63] ^ x[26];
  assign t[54] = t[64] ^ x[31];
  assign t[55] = t[65] ^ x[36];
  assign t[56] = t[66] ^ x[41];
  assign t[57] = t[67] ^ x[46];
  assign t[58] = t[68] ^ x[51];
  assign t[59] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[61] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[62] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[63] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[64] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[65] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[66] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[67] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[68] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[69] = t[109] ^ x[6];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[110] ^ x[3];
  assign t[71] = t[111] ^ x[4];
  assign t[72] = t[112] ^ x[5];
  assign t[73] = t[113] ^ x[11];
  assign t[74] = t[114] ^ x[8];
  assign t[75] = t[115] ^ x[9];
  assign t[76] = t[116] ^ x[10];
  assign t[77] = t[117] ^ x[16];
  assign t[78] = t[118] ^ x[13];
  assign t[79] = t[119] ^ x[14];
  assign t[7] = ~t[12];
  assign t[80] = t[120] ^ x[15];
  assign t[81] = t[121] ^ x[21];
  assign t[82] = t[122] ^ x[18];
  assign t[83] = t[123] ^ x[19];
  assign t[84] = t[124] ^ x[20];
  assign t[85] = t[125] ^ x[26];
  assign t[86] = t[126] ^ x[23];
  assign t[87] = t[127] ^ x[24];
  assign t[88] = t[128] ^ x[25];
  assign t[89] = t[129] ^ x[31];
  assign t[8] = t[40] & t[13];
  assign t[90] = t[130] ^ x[28];
  assign t[91] = t[131] ^ x[29];
  assign t[92] = t[132] ^ x[30];
  assign t[93] = t[133] ^ x[36];
  assign t[94] = t[134] ^ x[33];
  assign t[95] = t[135] ^ x[34];
  assign t[96] = t[136] ^ x[35];
  assign t[97] = t[137] ^ x[41];
  assign t[98] = t[138] ^ x[38];
  assign t[99] = t[139] ^ x[39];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind83(x, y);
 input [51:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ^ x[40];
  assign t[101] = t[141] ^ x[46];
  assign t[102] = t[142] ^ x[43];
  assign t[103] = t[143] ^ x[44];
  assign t[104] = t[144] ^ x[45];
  assign t[105] = t[145] ^ x[51];
  assign t[106] = t[146] ^ x[48];
  assign t[107] = t[147] ^ x[49];
  assign t[108] = t[148] ^ x[50];
  assign t[109] = (x[2]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[2]);
  assign t[111] = (x[2]);
  assign t[112] = (x[2]);
  assign t[113] = (x[7]);
  assign t[114] = (x[7]);
  assign t[115] = (x[7]);
  assign t[116] = (x[7]);
  assign t[117] = (x[12]);
  assign t[118] = (x[12]);
  assign t[119] = (x[12]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[12]);
  assign t[121] = (x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[17]);
  assign t[124] = (x[17]);
  assign t[125] = (x[22]);
  assign t[126] = (x[22]);
  assign t[127] = (x[22]);
  assign t[128] = (x[22]);
  assign t[129] = (x[27]);
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[130] = (x[27]);
  assign t[131] = (x[27]);
  assign t[132] = (x[27]);
  assign t[133] = (x[32]);
  assign t[134] = (x[32]);
  assign t[135] = (x[32]);
  assign t[136] = (x[32]);
  assign t[137] = (x[37]);
  assign t[138] = (x[37]);
  assign t[139] = (x[37]);
  assign t[13] = t[19] ^ t[20];
  assign t[140] = (x[37]);
  assign t[141] = (x[42]);
  assign t[142] = (x[42]);
  assign t[143] = (x[42]);
  assign t[144] = (x[42]);
  assign t[145] = (x[47]);
  assign t[146] = (x[47]);
  assign t[147] = (x[47]);
  assign t[148] = (x[47]);
  assign t[14] = ~(t[42]);
  assign t[15] = ~(t[40] ^ t[14]);
  assign t[16] = t[43] ^ t[42];
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[18] = ~t[22];
  assign t[19] = t[40] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[40] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[42] ^ t[44];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[45] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[45] ^ t[31]);
  assign t[33] = t[47] ^ t[46];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[45] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[45] ^ t[38];
  assign t[38] = t[46] ^ t[48];
  assign t[39] = (t[49]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[6];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[11];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[21];
  assign t[53] = t[63] ^ x[26];
  assign t[54] = t[64] ^ x[31];
  assign t[55] = t[65] ^ x[36];
  assign t[56] = t[66] ^ x[41];
  assign t[57] = t[67] ^ x[46];
  assign t[58] = t[68] ^ x[51];
  assign t[59] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[61] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[62] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[63] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[64] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[65] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[66] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[67] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[68] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[69] = t[109] ^ x[6];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[110] ^ x[3];
  assign t[71] = t[111] ^ x[4];
  assign t[72] = t[112] ^ x[5];
  assign t[73] = t[113] ^ x[11];
  assign t[74] = t[114] ^ x[8];
  assign t[75] = t[115] ^ x[9];
  assign t[76] = t[116] ^ x[10];
  assign t[77] = t[117] ^ x[16];
  assign t[78] = t[118] ^ x[13];
  assign t[79] = t[119] ^ x[14];
  assign t[7] = ~t[12];
  assign t[80] = t[120] ^ x[15];
  assign t[81] = t[121] ^ x[21];
  assign t[82] = t[122] ^ x[18];
  assign t[83] = t[123] ^ x[19];
  assign t[84] = t[124] ^ x[20];
  assign t[85] = t[125] ^ x[26];
  assign t[86] = t[126] ^ x[23];
  assign t[87] = t[127] ^ x[24];
  assign t[88] = t[128] ^ x[25];
  assign t[89] = t[129] ^ x[31];
  assign t[8] = t[40] & t[13];
  assign t[90] = t[130] ^ x[28];
  assign t[91] = t[131] ^ x[29];
  assign t[92] = t[132] ^ x[30];
  assign t[93] = t[133] ^ x[36];
  assign t[94] = t[134] ^ x[33];
  assign t[95] = t[135] ^ x[34];
  assign t[96] = t[136] ^ x[35];
  assign t[97] = t[137] ^ x[41];
  assign t[98] = t[138] ^ x[38];
  assign t[99] = t[139] ^ x[39];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind84(x, y);
 input [51:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ^ x[40];
  assign t[101] = t[141] ^ x[46];
  assign t[102] = t[142] ^ x[43];
  assign t[103] = t[143] ^ x[44];
  assign t[104] = t[144] ^ x[45];
  assign t[105] = t[145] ^ x[51];
  assign t[106] = t[146] ^ x[48];
  assign t[107] = t[147] ^ x[49];
  assign t[108] = t[148] ^ x[50];
  assign t[109] = (x[2]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[2]);
  assign t[111] = (x[2]);
  assign t[112] = (x[2]);
  assign t[113] = (x[7]);
  assign t[114] = (x[7]);
  assign t[115] = (x[7]);
  assign t[116] = (x[7]);
  assign t[117] = (x[12]);
  assign t[118] = (x[12]);
  assign t[119] = (x[12]);
  assign t[11] = t[40] ^ t[15];
  assign t[120] = (x[12]);
  assign t[121] = (x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[17]);
  assign t[124] = (x[17]);
  assign t[125] = (x[22]);
  assign t[126] = (x[22]);
  assign t[127] = (x[22]);
  assign t[128] = (x[22]);
  assign t[129] = (x[27]);
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[130] = (x[27]);
  assign t[131] = (x[27]);
  assign t[132] = (x[27]);
  assign t[133] = (x[32]);
  assign t[134] = (x[32]);
  assign t[135] = (x[32]);
  assign t[136] = (x[32]);
  assign t[137] = (x[37]);
  assign t[138] = (x[37]);
  assign t[139] = (x[37]);
  assign t[13] = t[42] ^ t[43];
  assign t[140] = (x[37]);
  assign t[141] = (x[42]);
  assign t[142] = (x[42]);
  assign t[143] = (x[42]);
  assign t[144] = (x[42]);
  assign t[145] = (x[47]);
  assign t[146] = (x[47]);
  assign t[147] = (x[47]);
  assign t[148] = (x[47]);
  assign t[14] = t[15] & t[19];
  assign t[15] = ~(t[43]);
  assign t[16] = ~(t[40] ^ t[15]);
  assign t[17] = t[40] & t[20];
  assign t[18] = ~t[21];
  assign t[19] = t[40] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] ^ t[14];
  assign t[21] = ~(t[24] ^ t[25]);
  assign t[22] = t[43] ^ t[44];
  assign t[23] = t[40] ^ t[13];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[34] ^ t[27];
  assign t[29] = t[45] ^ t[32];
  assign t[2] = ~t[4];
  assign t[30] = t[46] ^ t[47];
  assign t[31] = t[32] & t[35];
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[45] ^ t[32]);
  assign t[34] = t[45] & t[36];
  assign t[35] = t[45] ^ t[37];
  assign t[36] = t[38] ^ t[31];
  assign t[37] = t[47] ^ t[48];
  assign t[38] = t[45] ^ t[30];
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[6];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[11];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[21];
  assign t[53] = t[63] ^ x[26];
  assign t[54] = t[64] ^ x[31];
  assign t[55] = t[65] ^ x[36];
  assign t[56] = t[66] ^ x[41];
  assign t[57] = t[67] ^ x[46];
  assign t[58] = t[68] ^ x[51];
  assign t[59] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[61] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[62] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[63] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[64] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[65] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[66] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[67] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[68] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[69] = t[109] ^ x[6];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[110] ^ x[3];
  assign t[71] = t[111] ^ x[4];
  assign t[72] = t[112] ^ x[5];
  assign t[73] = t[113] ^ x[11];
  assign t[74] = t[114] ^ x[8];
  assign t[75] = t[115] ^ x[9];
  assign t[76] = t[116] ^ x[10];
  assign t[77] = t[117] ^ x[16];
  assign t[78] = t[118] ^ x[13];
  assign t[79] = t[119] ^ x[14];
  assign t[7] = ~t[12];
  assign t[80] = t[120] ^ x[15];
  assign t[81] = t[121] ^ x[21];
  assign t[82] = t[122] ^ x[18];
  assign t[83] = t[123] ^ x[19];
  assign t[84] = t[124] ^ x[20];
  assign t[85] = t[125] ^ x[26];
  assign t[86] = t[126] ^ x[23];
  assign t[87] = t[127] ^ x[24];
  assign t[88] = t[128] ^ x[25];
  assign t[89] = t[129] ^ x[31];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[130] ^ x[28];
  assign t[91] = t[131] ^ x[29];
  assign t[92] = t[132] ^ x[30];
  assign t[93] = t[133] ^ x[36];
  assign t[94] = t[134] ^ x[33];
  assign t[95] = t[135] ^ x[34];
  assign t[96] = t[136] ^ x[35];
  assign t[97] = t[137] ^ x[41];
  assign t[98] = t[138] ^ x[38];
  assign t[99] = t[139] ^ x[39];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind85(x, y);
 input [51:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ^ x[40];
  assign t[101] = t[141] ^ x[46];
  assign t[102] = t[142] ^ x[43];
  assign t[103] = t[143] ^ x[44];
  assign t[104] = t[144] ^ x[45];
  assign t[105] = t[145] ^ x[51];
  assign t[106] = t[146] ^ x[48];
  assign t[107] = t[147] ^ x[49];
  assign t[108] = t[148] ^ x[50];
  assign t[109] = (x[2]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[2]);
  assign t[111] = (x[2]);
  assign t[112] = (x[2]);
  assign t[113] = (x[7]);
  assign t[114] = (x[7]);
  assign t[115] = (x[7]);
  assign t[116] = (x[7]);
  assign t[117] = (x[12]);
  assign t[118] = (x[12]);
  assign t[119] = (x[12]);
  assign t[11] = t[40] ^ t[15];
  assign t[120] = (x[12]);
  assign t[121] = (x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[17]);
  assign t[124] = (x[17]);
  assign t[125] = (x[22]);
  assign t[126] = (x[22]);
  assign t[127] = (x[22]);
  assign t[128] = (x[22]);
  assign t[129] = (x[27]);
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[130] = (x[27]);
  assign t[131] = (x[27]);
  assign t[132] = (x[27]);
  assign t[133] = (x[32]);
  assign t[134] = (x[32]);
  assign t[135] = (x[32]);
  assign t[136] = (x[32]);
  assign t[137] = (x[37]);
  assign t[138] = (x[37]);
  assign t[139] = (x[37]);
  assign t[13] = t[42] ^ t[43];
  assign t[140] = (x[37]);
  assign t[141] = (x[42]);
  assign t[142] = (x[42]);
  assign t[143] = (x[42]);
  assign t[144] = (x[42]);
  assign t[145] = (x[47]);
  assign t[146] = (x[47]);
  assign t[147] = (x[47]);
  assign t[148] = (x[47]);
  assign t[14] = t[15] & t[19];
  assign t[15] = ~(t[43]);
  assign t[16] = ~(t[40] ^ t[15]);
  assign t[17] = t[40] & t[20];
  assign t[18] = ~t[21];
  assign t[19] = t[40] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] ^ t[14];
  assign t[21] = ~(t[24] ^ t[25]);
  assign t[22] = t[43] ^ t[44];
  assign t[23] = t[40] ^ t[13];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[34] ^ t[27];
  assign t[29] = t[45] ^ t[32];
  assign t[2] = ~t[4];
  assign t[30] = t[46] ^ t[47];
  assign t[31] = t[32] & t[35];
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[45] ^ t[32]);
  assign t[34] = t[45] & t[36];
  assign t[35] = t[45] ^ t[37];
  assign t[36] = t[38] ^ t[31];
  assign t[37] = t[47] ^ t[48];
  assign t[38] = t[45] ^ t[30];
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[6];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[11];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[21];
  assign t[53] = t[63] ^ x[26];
  assign t[54] = t[64] ^ x[31];
  assign t[55] = t[65] ^ x[36];
  assign t[56] = t[66] ^ x[41];
  assign t[57] = t[67] ^ x[46];
  assign t[58] = t[68] ^ x[51];
  assign t[59] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[61] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[62] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[63] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[64] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[65] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[66] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[67] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[68] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[69] = t[109] ^ x[6];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[110] ^ x[3];
  assign t[71] = t[111] ^ x[4];
  assign t[72] = t[112] ^ x[5];
  assign t[73] = t[113] ^ x[11];
  assign t[74] = t[114] ^ x[8];
  assign t[75] = t[115] ^ x[9];
  assign t[76] = t[116] ^ x[10];
  assign t[77] = t[117] ^ x[16];
  assign t[78] = t[118] ^ x[13];
  assign t[79] = t[119] ^ x[14];
  assign t[7] = ~t[12];
  assign t[80] = t[120] ^ x[15];
  assign t[81] = t[121] ^ x[21];
  assign t[82] = t[122] ^ x[18];
  assign t[83] = t[123] ^ x[19];
  assign t[84] = t[124] ^ x[20];
  assign t[85] = t[125] ^ x[26];
  assign t[86] = t[126] ^ x[23];
  assign t[87] = t[127] ^ x[24];
  assign t[88] = t[128] ^ x[25];
  assign t[89] = t[129] ^ x[31];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[130] ^ x[28];
  assign t[91] = t[131] ^ x[29];
  assign t[92] = t[132] ^ x[30];
  assign t[93] = t[133] ^ x[36];
  assign t[94] = t[134] ^ x[33];
  assign t[95] = t[135] ^ x[34];
  assign t[96] = t[136] ^ x[35];
  assign t[97] = t[137] ^ x[41];
  assign t[98] = t[138] ^ x[38];
  assign t[99] = t[139] ^ x[39];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind86(x, y);
 input [51:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ^ x[40];
  assign t[101] = t[141] ^ x[46];
  assign t[102] = t[142] ^ x[43];
  assign t[103] = t[143] ^ x[44];
  assign t[104] = t[144] ^ x[45];
  assign t[105] = t[145] ^ x[51];
  assign t[106] = t[146] ^ x[48];
  assign t[107] = t[147] ^ x[49];
  assign t[108] = t[148] ^ x[50];
  assign t[109] = (x[2]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[2]);
  assign t[111] = (x[2]);
  assign t[112] = (x[2]);
  assign t[113] = (x[7]);
  assign t[114] = (x[7]);
  assign t[115] = (x[7]);
  assign t[116] = (x[7]);
  assign t[117] = (x[12]);
  assign t[118] = (x[12]);
  assign t[119] = (x[12]);
  assign t[11] = t[40] ^ t[15];
  assign t[120] = (x[12]);
  assign t[121] = (x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[17]);
  assign t[124] = (x[17]);
  assign t[125] = (x[22]);
  assign t[126] = (x[22]);
  assign t[127] = (x[22]);
  assign t[128] = (x[22]);
  assign t[129] = (x[27]);
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[130] = (x[27]);
  assign t[131] = (x[27]);
  assign t[132] = (x[27]);
  assign t[133] = (x[32]);
  assign t[134] = (x[32]);
  assign t[135] = (x[32]);
  assign t[136] = (x[32]);
  assign t[137] = (x[37]);
  assign t[138] = (x[37]);
  assign t[139] = (x[37]);
  assign t[13] = t[42] ^ t[43];
  assign t[140] = (x[37]);
  assign t[141] = (x[42]);
  assign t[142] = (x[42]);
  assign t[143] = (x[42]);
  assign t[144] = (x[42]);
  assign t[145] = (x[47]);
  assign t[146] = (x[47]);
  assign t[147] = (x[47]);
  assign t[148] = (x[47]);
  assign t[14] = t[15] & t[19];
  assign t[15] = ~(t[43]);
  assign t[16] = ~(t[40] ^ t[15]);
  assign t[17] = t[40] & t[20];
  assign t[18] = ~t[21];
  assign t[19] = t[40] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] ^ t[14];
  assign t[21] = ~(t[24] ^ t[25]);
  assign t[22] = t[43] ^ t[44];
  assign t[23] = t[40] ^ t[13];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[34] ^ t[27];
  assign t[29] = t[45] ^ t[32];
  assign t[2] = ~t[4];
  assign t[30] = t[46] ^ t[47];
  assign t[31] = t[32] & t[35];
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[45] ^ t[32]);
  assign t[34] = t[45] & t[36];
  assign t[35] = t[45] ^ t[37];
  assign t[36] = t[38] ^ t[31];
  assign t[37] = t[47] ^ t[48];
  assign t[38] = t[45] ^ t[30];
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[6];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[11];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[21];
  assign t[53] = t[63] ^ x[26];
  assign t[54] = t[64] ^ x[31];
  assign t[55] = t[65] ^ x[36];
  assign t[56] = t[66] ^ x[41];
  assign t[57] = t[67] ^ x[46];
  assign t[58] = t[68] ^ x[51];
  assign t[59] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[61] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[62] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[63] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[64] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[65] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[66] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[67] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[68] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[69] = t[109] ^ x[6];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[110] ^ x[3];
  assign t[71] = t[111] ^ x[4];
  assign t[72] = t[112] ^ x[5];
  assign t[73] = t[113] ^ x[11];
  assign t[74] = t[114] ^ x[8];
  assign t[75] = t[115] ^ x[9];
  assign t[76] = t[116] ^ x[10];
  assign t[77] = t[117] ^ x[16];
  assign t[78] = t[118] ^ x[13];
  assign t[79] = t[119] ^ x[14];
  assign t[7] = ~t[12];
  assign t[80] = t[120] ^ x[15];
  assign t[81] = t[121] ^ x[21];
  assign t[82] = t[122] ^ x[18];
  assign t[83] = t[123] ^ x[19];
  assign t[84] = t[124] ^ x[20];
  assign t[85] = t[125] ^ x[26];
  assign t[86] = t[126] ^ x[23];
  assign t[87] = t[127] ^ x[24];
  assign t[88] = t[128] ^ x[25];
  assign t[89] = t[129] ^ x[31];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[130] ^ x[28];
  assign t[91] = t[131] ^ x[29];
  assign t[92] = t[132] ^ x[30];
  assign t[93] = t[133] ^ x[36];
  assign t[94] = t[134] ^ x[33];
  assign t[95] = t[135] ^ x[34];
  assign t[96] = t[136] ^ x[35];
  assign t[97] = t[137] ^ x[41];
  assign t[98] = t[138] ^ x[38];
  assign t[99] = t[139] ^ x[39];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind87(x, y);
 input [51:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ^ x[40];
  assign t[101] = t[141] ^ x[46];
  assign t[102] = t[142] ^ x[43];
  assign t[103] = t[143] ^ x[44];
  assign t[104] = t[144] ^ x[45];
  assign t[105] = t[145] ^ x[51];
  assign t[106] = t[146] ^ x[48];
  assign t[107] = t[147] ^ x[49];
  assign t[108] = t[148] ^ x[50];
  assign t[109] = (x[2]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[2]);
  assign t[111] = (x[2]);
  assign t[112] = (x[2]);
  assign t[113] = (x[7]);
  assign t[114] = (x[7]);
  assign t[115] = (x[7]);
  assign t[116] = (x[7]);
  assign t[117] = (x[12]);
  assign t[118] = (x[12]);
  assign t[119] = (x[12]);
  assign t[11] = t[40] ^ t[15];
  assign t[120] = (x[12]);
  assign t[121] = (x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[17]);
  assign t[124] = (x[17]);
  assign t[125] = (x[22]);
  assign t[126] = (x[22]);
  assign t[127] = (x[22]);
  assign t[128] = (x[22]);
  assign t[129] = (x[27]);
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[130] = (x[27]);
  assign t[131] = (x[27]);
  assign t[132] = (x[27]);
  assign t[133] = (x[32]);
  assign t[134] = (x[32]);
  assign t[135] = (x[32]);
  assign t[136] = (x[32]);
  assign t[137] = (x[37]);
  assign t[138] = (x[37]);
  assign t[139] = (x[37]);
  assign t[13] = t[42] ^ t[43];
  assign t[140] = (x[37]);
  assign t[141] = (x[42]);
  assign t[142] = (x[42]);
  assign t[143] = (x[42]);
  assign t[144] = (x[42]);
  assign t[145] = (x[47]);
  assign t[146] = (x[47]);
  assign t[147] = (x[47]);
  assign t[148] = (x[47]);
  assign t[14] = t[15] & t[19];
  assign t[15] = ~(t[43]);
  assign t[16] = ~(t[40] ^ t[15]);
  assign t[17] = t[40] & t[20];
  assign t[18] = ~t[21];
  assign t[19] = t[40] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] ^ t[14];
  assign t[21] = ~(t[24] ^ t[25]);
  assign t[22] = t[43] ^ t[44];
  assign t[23] = t[40] ^ t[13];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[34] ^ t[27];
  assign t[29] = t[45] ^ t[32];
  assign t[2] = ~t[4];
  assign t[30] = t[46] ^ t[47];
  assign t[31] = t[32] & t[35];
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[45] ^ t[32]);
  assign t[34] = t[45] & t[36];
  assign t[35] = t[45] ^ t[37];
  assign t[36] = t[38] ^ t[31];
  assign t[37] = t[47] ^ t[48];
  assign t[38] = t[45] ^ t[30];
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[6];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[11];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[21];
  assign t[53] = t[63] ^ x[26];
  assign t[54] = t[64] ^ x[31];
  assign t[55] = t[65] ^ x[36];
  assign t[56] = t[66] ^ x[41];
  assign t[57] = t[67] ^ x[46];
  assign t[58] = t[68] ^ x[51];
  assign t[59] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[61] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[62] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[63] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[64] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[65] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[66] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[67] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[68] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[69] = t[109] ^ x[6];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[110] ^ x[3];
  assign t[71] = t[111] ^ x[4];
  assign t[72] = t[112] ^ x[5];
  assign t[73] = t[113] ^ x[11];
  assign t[74] = t[114] ^ x[8];
  assign t[75] = t[115] ^ x[9];
  assign t[76] = t[116] ^ x[10];
  assign t[77] = t[117] ^ x[16];
  assign t[78] = t[118] ^ x[13];
  assign t[79] = t[119] ^ x[14];
  assign t[7] = ~t[12];
  assign t[80] = t[120] ^ x[15];
  assign t[81] = t[121] ^ x[21];
  assign t[82] = t[122] ^ x[18];
  assign t[83] = t[123] ^ x[19];
  assign t[84] = t[124] ^ x[20];
  assign t[85] = t[125] ^ x[26];
  assign t[86] = t[126] ^ x[23];
  assign t[87] = t[127] ^ x[24];
  assign t[88] = t[128] ^ x[25];
  assign t[89] = t[129] ^ x[31];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[130] ^ x[28];
  assign t[91] = t[131] ^ x[29];
  assign t[92] = t[132] ^ x[30];
  assign t[93] = t[133] ^ x[36];
  assign t[94] = t[134] ^ x[33];
  assign t[95] = t[135] ^ x[34];
  assign t[96] = t[136] ^ x[35];
  assign t[97] = t[137] ^ x[41];
  assign t[98] = t[138] ^ x[38];
  assign t[99] = t[139] ^ x[39];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind88(x, y);
 input [41:0] x;
 output y;

 wire [106:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[32]);
  assign t[101] = (x[32]);
  assign t[102] = (x[32]);
  assign t[103] = (x[37]);
  assign t[104] = (x[37]);
  assign t[105] = (x[37]);
  assign t[106] = (x[37]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[23] ^ t[10]);
  assign t[12] = ~t[13];
  assign t[13] = ~(t[14]);
  assign t[14] = t[15] ^ t[16];
  assign t[15] = t[24] ^ t[25];
  assign t[16] = t[17] & t[18];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[26] ^ t[17]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = (t[30]);
  assign t[23] = (t[31]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = t[35] ^ x[6];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = t[37] ^ x[16];
  assign t[2] = ~t[4];
  assign t[30] = t[38] ^ x[21];
  assign t[31] = t[39] ^ x[26];
  assign t[32] = t[40] ^ x[31];
  assign t[33] = t[41] ^ x[36];
  assign t[34] = t[42] ^ x[41];
  assign t[35] = (~t[43] & t[44] & t[45] & t[46]) | (t[43] & ~t[45] & ~t[46]) | (t[43] & ~t[44] & ~t[46]) | (t[43] & ~t[44] & ~t[45]);
  assign t[36] = (~t[47] & t[48] & t[49] & t[50]) | (t[47] & ~t[49] & ~t[50]) | (t[47] & ~t[48] & ~t[50]) | (t[47] & ~t[48] & ~t[49]);
  assign t[37] = (~t[51] & t[52] & t[53] & t[54]) | (t[51] & ~t[53] & ~t[54]) | (t[51] & ~t[52] & ~t[54]) | (t[51] & ~t[52] & ~t[53]);
  assign t[38] = (~t[55] & t[56] & t[57] & t[58]) | (t[55] & ~t[57] & ~t[58]) | (t[55] & ~t[56] & ~t[58]) | (t[55] & ~t[56] & ~t[57]);
  assign t[39] = (~t[59] & t[60] & t[61] & t[62]) | (t[59] & ~t[61] & ~t[62]) | (t[59] & ~t[60] & ~t[62]) | (t[59] & ~t[60] & ~t[61]);
  assign t[3] = ~(t[5]);
  assign t[40] = (~t[63] & t[64] & t[65] & t[66]) | (t[63] & ~t[65] & ~t[66]) | (t[63] & ~t[64] & ~t[66]) | (t[63] & ~t[64] & ~t[65]);
  assign t[41] = (~t[67] & t[68] & t[69] & t[70]) | (t[67] & ~t[69] & ~t[70]) | (t[67] & ~t[68] & ~t[70]) | (t[67] & ~t[68] & ~t[69]);
  assign t[42] = (~t[71] & t[72] & t[73] & t[74]) | (t[71] & ~t[73] & ~t[74]) | (t[71] & ~t[72] & ~t[74]) | (t[71] & ~t[72] & ~t[73]);
  assign t[43] = t[75] ^ x[6];
  assign t[44] = t[76] ^ x[3];
  assign t[45] = t[77] ^ x[4];
  assign t[46] = t[78] ^ x[5];
  assign t[47] = t[79] ^ x[11];
  assign t[48] = t[80] ^ x[8];
  assign t[49] = t[81] ^ x[9];
  assign t[4] = ~(t[6] ^ t[19]);
  assign t[50] = t[82] ^ x[10];
  assign t[51] = t[83] ^ x[16];
  assign t[52] = t[84] ^ x[13];
  assign t[53] = t[85] ^ x[14];
  assign t[54] = t[86] ^ x[15];
  assign t[55] = t[87] ^ x[21];
  assign t[56] = t[88] ^ x[18];
  assign t[57] = t[89] ^ x[19];
  assign t[58] = t[90] ^ x[20];
  assign t[59] = t[91] ^ x[26];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[92] ^ x[23];
  assign t[61] = t[93] ^ x[24];
  assign t[62] = t[94] ^ x[25];
  assign t[63] = t[95] ^ x[31];
  assign t[64] = t[96] ^ x[28];
  assign t[65] = t[97] ^ x[29];
  assign t[66] = t[98] ^ x[30];
  assign t[67] = t[99] ^ x[36];
  assign t[68] = t[100] ^ x[33];
  assign t[69] = t[101] ^ x[34];
  assign t[6] = ~t[9];
  assign t[70] = t[102] ^ x[35];
  assign t[71] = t[103] ^ x[41];
  assign t[72] = t[104] ^ x[38];
  assign t[73] = t[105] ^ x[39];
  assign t[74] = t[106] ^ x[40];
  assign t[75] = (x[2]);
  assign t[76] = (x[2]);
  assign t[77] = (x[2]);
  assign t[78] = (x[2]);
  assign t[79] = (x[7]);
  assign t[7] = t[20] ^ t[21];
  assign t[80] = (x[7]);
  assign t[81] = (x[7]);
  assign t[82] = (x[7]);
  assign t[83] = (x[12]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[12]);
  assign t[87] = (x[17]);
  assign t[88] = (x[17]);
  assign t[89] = (x[17]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[17]);
  assign t[91] = (x[22]);
  assign t[92] = (x[22]);
  assign t[93] = (x[22]);
  assign t[94] = (x[22]);
  assign t[95] = (x[27]);
  assign t[96] = (x[27]);
  assign t[97] = (x[27]);
  assign t[98] = (x[27]);
  assign t[99] = (x[32]);
  assign t[9] = ~(t[12] ^ t[22]);
  assign y = (t[0]);
endmodule

module R2ind89(x, y);
 input [41:0] x;
 output y;

 wire [106:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[32]);
  assign t[101] = (x[32]);
  assign t[102] = (x[32]);
  assign t[103] = (x[37]);
  assign t[104] = (x[37]);
  assign t[105] = (x[37]);
  assign t[106] = (x[37]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[23] ^ t[10]);
  assign t[12] = ~t[13];
  assign t[13] = ~(t[14]);
  assign t[14] = t[15] ^ t[16];
  assign t[15] = t[24] ^ t[25];
  assign t[16] = t[17] & t[18];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[26] ^ t[17]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = (t[30]);
  assign t[23] = (t[31]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = t[35] ^ x[6];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = t[37] ^ x[16];
  assign t[2] = ~t[4];
  assign t[30] = t[38] ^ x[21];
  assign t[31] = t[39] ^ x[26];
  assign t[32] = t[40] ^ x[31];
  assign t[33] = t[41] ^ x[36];
  assign t[34] = t[42] ^ x[41];
  assign t[35] = (~t[43] & t[44] & t[45] & t[46]) | (t[43] & ~t[45] & ~t[46]) | (t[43] & ~t[44] & ~t[46]) | (t[43] & ~t[44] & ~t[45]);
  assign t[36] = (~t[47] & t[48] & t[49] & t[50]) | (t[47] & ~t[49] & ~t[50]) | (t[47] & ~t[48] & ~t[50]) | (t[47] & ~t[48] & ~t[49]);
  assign t[37] = (~t[51] & t[52] & t[53] & t[54]) | (t[51] & ~t[53] & ~t[54]) | (t[51] & ~t[52] & ~t[54]) | (t[51] & ~t[52] & ~t[53]);
  assign t[38] = (~t[55] & t[56] & t[57] & t[58]) | (t[55] & ~t[57] & ~t[58]) | (t[55] & ~t[56] & ~t[58]) | (t[55] & ~t[56] & ~t[57]);
  assign t[39] = (~t[59] & t[60] & t[61] & t[62]) | (t[59] & ~t[61] & ~t[62]) | (t[59] & ~t[60] & ~t[62]) | (t[59] & ~t[60] & ~t[61]);
  assign t[3] = ~(t[5]);
  assign t[40] = (~t[63] & t[64] & t[65] & t[66]) | (t[63] & ~t[65] & ~t[66]) | (t[63] & ~t[64] & ~t[66]) | (t[63] & ~t[64] & ~t[65]);
  assign t[41] = (~t[67] & t[68] & t[69] & t[70]) | (t[67] & ~t[69] & ~t[70]) | (t[67] & ~t[68] & ~t[70]) | (t[67] & ~t[68] & ~t[69]);
  assign t[42] = (~t[71] & t[72] & t[73] & t[74]) | (t[71] & ~t[73] & ~t[74]) | (t[71] & ~t[72] & ~t[74]) | (t[71] & ~t[72] & ~t[73]);
  assign t[43] = t[75] ^ x[6];
  assign t[44] = t[76] ^ x[3];
  assign t[45] = t[77] ^ x[4];
  assign t[46] = t[78] ^ x[5];
  assign t[47] = t[79] ^ x[11];
  assign t[48] = t[80] ^ x[8];
  assign t[49] = t[81] ^ x[9];
  assign t[4] = ~(t[6] ^ t[19]);
  assign t[50] = t[82] ^ x[10];
  assign t[51] = t[83] ^ x[16];
  assign t[52] = t[84] ^ x[13];
  assign t[53] = t[85] ^ x[14];
  assign t[54] = t[86] ^ x[15];
  assign t[55] = t[87] ^ x[21];
  assign t[56] = t[88] ^ x[18];
  assign t[57] = t[89] ^ x[19];
  assign t[58] = t[90] ^ x[20];
  assign t[59] = t[91] ^ x[26];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[92] ^ x[23];
  assign t[61] = t[93] ^ x[24];
  assign t[62] = t[94] ^ x[25];
  assign t[63] = t[95] ^ x[31];
  assign t[64] = t[96] ^ x[28];
  assign t[65] = t[97] ^ x[29];
  assign t[66] = t[98] ^ x[30];
  assign t[67] = t[99] ^ x[36];
  assign t[68] = t[100] ^ x[33];
  assign t[69] = t[101] ^ x[34];
  assign t[6] = ~t[9];
  assign t[70] = t[102] ^ x[35];
  assign t[71] = t[103] ^ x[41];
  assign t[72] = t[104] ^ x[38];
  assign t[73] = t[105] ^ x[39];
  assign t[74] = t[106] ^ x[40];
  assign t[75] = (x[2]);
  assign t[76] = (x[2]);
  assign t[77] = (x[2]);
  assign t[78] = (x[2]);
  assign t[79] = (x[7]);
  assign t[7] = t[20] ^ t[21];
  assign t[80] = (x[7]);
  assign t[81] = (x[7]);
  assign t[82] = (x[7]);
  assign t[83] = (x[12]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[12]);
  assign t[87] = (x[17]);
  assign t[88] = (x[17]);
  assign t[89] = (x[17]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[17]);
  assign t[91] = (x[22]);
  assign t[92] = (x[22]);
  assign t[93] = (x[22]);
  assign t[94] = (x[22]);
  assign t[95] = (x[27]);
  assign t[96] = (x[27]);
  assign t[97] = (x[27]);
  assign t[98] = (x[27]);
  assign t[99] = (x[32]);
  assign t[9] = ~(t[12] ^ t[22]);
  assign y = (t[0]);
endmodule

module R2ind90(x, y);
 input [41:0] x;
 output y;

 wire [106:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[32]);
  assign t[101] = (x[32]);
  assign t[102] = (x[32]);
  assign t[103] = (x[37]);
  assign t[104] = (x[37]);
  assign t[105] = (x[37]);
  assign t[106] = (x[37]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[23] ^ t[10]);
  assign t[12] = ~t[13];
  assign t[13] = ~(t[14]);
  assign t[14] = t[15] ^ t[16];
  assign t[15] = t[24] ^ t[25];
  assign t[16] = t[17] & t[18];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[26] ^ t[17]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = (t[30]);
  assign t[23] = (t[31]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = t[35] ^ x[6];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = t[37] ^ x[16];
  assign t[2] = ~t[4];
  assign t[30] = t[38] ^ x[21];
  assign t[31] = t[39] ^ x[26];
  assign t[32] = t[40] ^ x[31];
  assign t[33] = t[41] ^ x[36];
  assign t[34] = t[42] ^ x[41];
  assign t[35] = (~t[43] & t[44] & t[45] & t[46]) | (t[43] & ~t[45] & ~t[46]) | (t[43] & ~t[44] & ~t[46]) | (t[43] & ~t[44] & ~t[45]);
  assign t[36] = (~t[47] & t[48] & t[49] & t[50]) | (t[47] & ~t[49] & ~t[50]) | (t[47] & ~t[48] & ~t[50]) | (t[47] & ~t[48] & ~t[49]);
  assign t[37] = (~t[51] & t[52] & t[53] & t[54]) | (t[51] & ~t[53] & ~t[54]) | (t[51] & ~t[52] & ~t[54]) | (t[51] & ~t[52] & ~t[53]);
  assign t[38] = (~t[55] & t[56] & t[57] & t[58]) | (t[55] & ~t[57] & ~t[58]) | (t[55] & ~t[56] & ~t[58]) | (t[55] & ~t[56] & ~t[57]);
  assign t[39] = (~t[59] & t[60] & t[61] & t[62]) | (t[59] & ~t[61] & ~t[62]) | (t[59] & ~t[60] & ~t[62]) | (t[59] & ~t[60] & ~t[61]);
  assign t[3] = ~(t[5]);
  assign t[40] = (~t[63] & t[64] & t[65] & t[66]) | (t[63] & ~t[65] & ~t[66]) | (t[63] & ~t[64] & ~t[66]) | (t[63] & ~t[64] & ~t[65]);
  assign t[41] = (~t[67] & t[68] & t[69] & t[70]) | (t[67] & ~t[69] & ~t[70]) | (t[67] & ~t[68] & ~t[70]) | (t[67] & ~t[68] & ~t[69]);
  assign t[42] = (~t[71] & t[72] & t[73] & t[74]) | (t[71] & ~t[73] & ~t[74]) | (t[71] & ~t[72] & ~t[74]) | (t[71] & ~t[72] & ~t[73]);
  assign t[43] = t[75] ^ x[6];
  assign t[44] = t[76] ^ x[3];
  assign t[45] = t[77] ^ x[4];
  assign t[46] = t[78] ^ x[5];
  assign t[47] = t[79] ^ x[11];
  assign t[48] = t[80] ^ x[8];
  assign t[49] = t[81] ^ x[9];
  assign t[4] = ~(t[6] ^ t[19]);
  assign t[50] = t[82] ^ x[10];
  assign t[51] = t[83] ^ x[16];
  assign t[52] = t[84] ^ x[13];
  assign t[53] = t[85] ^ x[14];
  assign t[54] = t[86] ^ x[15];
  assign t[55] = t[87] ^ x[21];
  assign t[56] = t[88] ^ x[18];
  assign t[57] = t[89] ^ x[19];
  assign t[58] = t[90] ^ x[20];
  assign t[59] = t[91] ^ x[26];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[92] ^ x[23];
  assign t[61] = t[93] ^ x[24];
  assign t[62] = t[94] ^ x[25];
  assign t[63] = t[95] ^ x[31];
  assign t[64] = t[96] ^ x[28];
  assign t[65] = t[97] ^ x[29];
  assign t[66] = t[98] ^ x[30];
  assign t[67] = t[99] ^ x[36];
  assign t[68] = t[100] ^ x[33];
  assign t[69] = t[101] ^ x[34];
  assign t[6] = ~t[9];
  assign t[70] = t[102] ^ x[35];
  assign t[71] = t[103] ^ x[41];
  assign t[72] = t[104] ^ x[38];
  assign t[73] = t[105] ^ x[39];
  assign t[74] = t[106] ^ x[40];
  assign t[75] = (x[2]);
  assign t[76] = (x[2]);
  assign t[77] = (x[2]);
  assign t[78] = (x[2]);
  assign t[79] = (x[7]);
  assign t[7] = t[20] ^ t[21];
  assign t[80] = (x[7]);
  assign t[81] = (x[7]);
  assign t[82] = (x[7]);
  assign t[83] = (x[12]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[12]);
  assign t[87] = (x[17]);
  assign t[88] = (x[17]);
  assign t[89] = (x[17]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[17]);
  assign t[91] = (x[22]);
  assign t[92] = (x[22]);
  assign t[93] = (x[22]);
  assign t[94] = (x[22]);
  assign t[95] = (x[27]);
  assign t[96] = (x[27]);
  assign t[97] = (x[27]);
  assign t[98] = (x[27]);
  assign t[99] = (x[32]);
  assign t[9] = ~(t[12] ^ t[22]);
  assign y = (t[0]);
endmodule

module R2ind91(x, y);
 input [41:0] x;
 output y;

 wire [106:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[32]);
  assign t[101] = (x[32]);
  assign t[102] = (x[32]);
  assign t[103] = (x[37]);
  assign t[104] = (x[37]);
  assign t[105] = (x[37]);
  assign t[106] = (x[37]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[23] ^ t[10]);
  assign t[12] = ~t[13];
  assign t[13] = ~(t[14]);
  assign t[14] = t[15] ^ t[16];
  assign t[15] = t[24] ^ t[25];
  assign t[16] = t[17] & t[18];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[26] ^ t[17]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = (t[30]);
  assign t[23] = (t[31]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = t[35] ^ x[6];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = t[37] ^ x[16];
  assign t[2] = ~t[4];
  assign t[30] = t[38] ^ x[21];
  assign t[31] = t[39] ^ x[26];
  assign t[32] = t[40] ^ x[31];
  assign t[33] = t[41] ^ x[36];
  assign t[34] = t[42] ^ x[41];
  assign t[35] = (~t[43] & t[44] & t[45] & t[46]) | (t[43] & ~t[45] & ~t[46]) | (t[43] & ~t[44] & ~t[46]) | (t[43] & ~t[44] & ~t[45]);
  assign t[36] = (~t[47] & t[48] & t[49] & t[50]) | (t[47] & ~t[49] & ~t[50]) | (t[47] & ~t[48] & ~t[50]) | (t[47] & ~t[48] & ~t[49]);
  assign t[37] = (~t[51] & t[52] & t[53] & t[54]) | (t[51] & ~t[53] & ~t[54]) | (t[51] & ~t[52] & ~t[54]) | (t[51] & ~t[52] & ~t[53]);
  assign t[38] = (~t[55] & t[56] & t[57] & t[58]) | (t[55] & ~t[57] & ~t[58]) | (t[55] & ~t[56] & ~t[58]) | (t[55] & ~t[56] & ~t[57]);
  assign t[39] = (~t[59] & t[60] & t[61] & t[62]) | (t[59] & ~t[61] & ~t[62]) | (t[59] & ~t[60] & ~t[62]) | (t[59] & ~t[60] & ~t[61]);
  assign t[3] = ~(t[5]);
  assign t[40] = (~t[63] & t[64] & t[65] & t[66]) | (t[63] & ~t[65] & ~t[66]) | (t[63] & ~t[64] & ~t[66]) | (t[63] & ~t[64] & ~t[65]);
  assign t[41] = (~t[67] & t[68] & t[69] & t[70]) | (t[67] & ~t[69] & ~t[70]) | (t[67] & ~t[68] & ~t[70]) | (t[67] & ~t[68] & ~t[69]);
  assign t[42] = (~t[71] & t[72] & t[73] & t[74]) | (t[71] & ~t[73] & ~t[74]) | (t[71] & ~t[72] & ~t[74]) | (t[71] & ~t[72] & ~t[73]);
  assign t[43] = t[75] ^ x[6];
  assign t[44] = t[76] ^ x[3];
  assign t[45] = t[77] ^ x[4];
  assign t[46] = t[78] ^ x[5];
  assign t[47] = t[79] ^ x[11];
  assign t[48] = t[80] ^ x[8];
  assign t[49] = t[81] ^ x[9];
  assign t[4] = ~(t[6] ^ t[19]);
  assign t[50] = t[82] ^ x[10];
  assign t[51] = t[83] ^ x[16];
  assign t[52] = t[84] ^ x[13];
  assign t[53] = t[85] ^ x[14];
  assign t[54] = t[86] ^ x[15];
  assign t[55] = t[87] ^ x[21];
  assign t[56] = t[88] ^ x[18];
  assign t[57] = t[89] ^ x[19];
  assign t[58] = t[90] ^ x[20];
  assign t[59] = t[91] ^ x[26];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[92] ^ x[23];
  assign t[61] = t[93] ^ x[24];
  assign t[62] = t[94] ^ x[25];
  assign t[63] = t[95] ^ x[31];
  assign t[64] = t[96] ^ x[28];
  assign t[65] = t[97] ^ x[29];
  assign t[66] = t[98] ^ x[30];
  assign t[67] = t[99] ^ x[36];
  assign t[68] = t[100] ^ x[33];
  assign t[69] = t[101] ^ x[34];
  assign t[6] = ~t[9];
  assign t[70] = t[102] ^ x[35];
  assign t[71] = t[103] ^ x[41];
  assign t[72] = t[104] ^ x[38];
  assign t[73] = t[105] ^ x[39];
  assign t[74] = t[106] ^ x[40];
  assign t[75] = (x[2]);
  assign t[76] = (x[2]);
  assign t[77] = (x[2]);
  assign t[78] = (x[2]);
  assign t[79] = (x[7]);
  assign t[7] = t[20] ^ t[21];
  assign t[80] = (x[7]);
  assign t[81] = (x[7]);
  assign t[82] = (x[7]);
  assign t[83] = (x[12]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[12]);
  assign t[87] = (x[17]);
  assign t[88] = (x[17]);
  assign t[89] = (x[17]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[17]);
  assign t[91] = (x[22]);
  assign t[92] = (x[22]);
  assign t[93] = (x[22]);
  assign t[94] = (x[22]);
  assign t[95] = (x[27]);
  assign t[96] = (x[27]);
  assign t[97] = (x[27]);
  assign t[98] = (x[27]);
  assign t[99] = (x[32]);
  assign t[9] = ~(t[12] ^ t[22]);
  assign y = (t[0]);
endmodule

module R2ind92(x, y);
 input [51:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[7]);
  assign t[102] = (x[7]);
  assign t[103] = (x[7]);
  assign t[104] = (x[7]);
  assign t[105] = (x[12]);
  assign t[106] = (x[12]);
  assign t[107] = (x[12]);
  assign t[108] = (x[12]);
  assign t[109] = (x[17]);
  assign t[10] = t[29] ^ t[30];
  assign t[110] = (x[17]);
  assign t[111] = (x[17]);
  assign t[112] = (x[17]);
  assign t[113] = (x[22]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[22]);
  assign t[117] = (x[27]);
  assign t[118] = (x[27]);
  assign t[119] = (x[27]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[32]);
  assign t[122] = (x[32]);
  assign t[123] = (x[32]);
  assign t[124] = (x[32]);
  assign t[125] = (x[37]);
  assign t[126] = (x[37]);
  assign t[127] = (x[37]);
  assign t[128] = (x[37]);
  assign t[129] = (x[42]);
  assign t[12] = ~(t[30]);
  assign t[130] = (x[42]);
  assign t[131] = (x[42]);
  assign t[132] = (x[42]);
  assign t[133] = (x[47]);
  assign t[134] = (x[47]);
  assign t[135] = (x[47]);
  assign t[136] = (x[47]);
  assign t[13] = ~(t[31] ^ t[12]);
  assign t[14] = ~t[16];
  assign t[15] = t[31] ^ t[17];
  assign t[16] = ~(t[18]);
  assign t[17] = t[30] ^ t[32];
  assign t[18] = t[19] ^ t[20];
  assign t[19] = t[21] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] & t[24];
  assign t[21] = t[33] ^ t[34];
  assign t[22] = t[23] & t[25];
  assign t[23] = ~(t[34]);
  assign t[24] = ~(t[35] ^ t[23]);
  assign t[25] = t[35] ^ t[26];
  assign t[26] = t[34] ^ t[36];
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~t[4];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = t[47] ^ x[6];
  assign t[38] = t[48] ^ x[11];
  assign t[39] = t[49] ^ x[16];
  assign t[3] = ~(t[5]);
  assign t[40] = t[50] ^ x[21];
  assign t[41] = t[51] ^ x[26];
  assign t[42] = t[52] ^ x[31];
  assign t[43] = t[53] ^ x[36];
  assign t[44] = t[54] ^ x[41];
  assign t[45] = t[55] ^ x[46];
  assign t[46] = t[56] ^ x[51];
  assign t[47] = (~t[57] & t[58] & t[59] & t[60]) | (t[57] & ~t[59] & ~t[60]) | (t[57] & ~t[58] & ~t[60]) | (t[57] & ~t[58] & ~t[59]);
  assign t[48] = (~t[61] & t[62] & t[63] & t[64]) | (t[61] & ~t[63] & ~t[64]) | (t[61] & ~t[62] & ~t[64]) | (t[61] & ~t[62] & ~t[63]);
  assign t[49] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[4] = ~(t[6] ^ t[27]);
  assign t[50] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[51] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[52] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[53] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[54] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[55] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[56] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[57] = t[97] ^ x[6];
  assign t[58] = t[98] ^ x[3];
  assign t[59] = t[99] ^ x[4];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[100] ^ x[5];
  assign t[61] = t[101] ^ x[11];
  assign t[62] = t[102] ^ x[8];
  assign t[63] = t[103] ^ x[9];
  assign t[64] = t[104] ^ x[10];
  assign t[65] = t[105] ^ x[16];
  assign t[66] = t[106] ^ x[13];
  assign t[67] = t[107] ^ x[14];
  assign t[68] = t[108] ^ x[15];
  assign t[69] = t[109] ^ x[21];
  assign t[6] = ~t[9];
  assign t[70] = t[110] ^ x[18];
  assign t[71] = t[111] ^ x[19];
  assign t[72] = t[112] ^ x[20];
  assign t[73] = t[113] ^ x[26];
  assign t[74] = t[114] ^ x[23];
  assign t[75] = t[115] ^ x[24];
  assign t[76] = t[116] ^ x[25];
  assign t[77] = t[117] ^ x[31];
  assign t[78] = t[118] ^ x[28];
  assign t[79] = t[119] ^ x[29];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[120] ^ x[30];
  assign t[81] = t[121] ^ x[36];
  assign t[82] = t[122] ^ x[33];
  assign t[83] = t[123] ^ x[34];
  assign t[84] = t[124] ^ x[35];
  assign t[85] = t[125] ^ x[41];
  assign t[86] = t[126] ^ x[38];
  assign t[87] = t[127] ^ x[39];
  assign t[88] = t[128] ^ x[40];
  assign t[89] = t[129] ^ x[46];
  assign t[8] = t[12] & t[13];
  assign t[90] = t[130] ^ x[43];
  assign t[91] = t[131] ^ x[44];
  assign t[92] = t[132] ^ x[45];
  assign t[93] = t[133] ^ x[51];
  assign t[94] = t[134] ^ x[48];
  assign t[95] = t[135] ^ x[49];
  assign t[96] = t[136] ^ x[50];
  assign t[97] = (x[2]);
  assign t[98] = (x[2]);
  assign t[99] = (x[2]);
  assign t[9] = ~(t[14] ^ t[28]);
  assign y = (t[0]);
endmodule

module R2ind93(x, y);
 input [51:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[7]);
  assign t[102] = (x[7]);
  assign t[103] = (x[7]);
  assign t[104] = (x[7]);
  assign t[105] = (x[12]);
  assign t[106] = (x[12]);
  assign t[107] = (x[12]);
  assign t[108] = (x[12]);
  assign t[109] = (x[17]);
  assign t[10] = t[29] ^ t[30];
  assign t[110] = (x[17]);
  assign t[111] = (x[17]);
  assign t[112] = (x[17]);
  assign t[113] = (x[22]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[22]);
  assign t[117] = (x[27]);
  assign t[118] = (x[27]);
  assign t[119] = (x[27]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[32]);
  assign t[122] = (x[32]);
  assign t[123] = (x[32]);
  assign t[124] = (x[32]);
  assign t[125] = (x[37]);
  assign t[126] = (x[37]);
  assign t[127] = (x[37]);
  assign t[128] = (x[37]);
  assign t[129] = (x[42]);
  assign t[12] = ~(t[30]);
  assign t[130] = (x[42]);
  assign t[131] = (x[42]);
  assign t[132] = (x[42]);
  assign t[133] = (x[47]);
  assign t[134] = (x[47]);
  assign t[135] = (x[47]);
  assign t[136] = (x[47]);
  assign t[13] = ~(t[31] ^ t[12]);
  assign t[14] = ~t[16];
  assign t[15] = t[31] ^ t[17];
  assign t[16] = ~(t[18]);
  assign t[17] = t[30] ^ t[32];
  assign t[18] = t[19] ^ t[20];
  assign t[19] = t[21] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] & t[24];
  assign t[21] = t[33] ^ t[34];
  assign t[22] = t[23] & t[25];
  assign t[23] = ~(t[34]);
  assign t[24] = ~(t[35] ^ t[23]);
  assign t[25] = t[35] ^ t[26];
  assign t[26] = t[34] ^ t[36];
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~t[4];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = t[47] ^ x[6];
  assign t[38] = t[48] ^ x[11];
  assign t[39] = t[49] ^ x[16];
  assign t[3] = ~(t[5]);
  assign t[40] = t[50] ^ x[21];
  assign t[41] = t[51] ^ x[26];
  assign t[42] = t[52] ^ x[31];
  assign t[43] = t[53] ^ x[36];
  assign t[44] = t[54] ^ x[41];
  assign t[45] = t[55] ^ x[46];
  assign t[46] = t[56] ^ x[51];
  assign t[47] = (~t[57] & t[58] & t[59] & t[60]) | (t[57] & ~t[59] & ~t[60]) | (t[57] & ~t[58] & ~t[60]) | (t[57] & ~t[58] & ~t[59]);
  assign t[48] = (~t[61] & t[62] & t[63] & t[64]) | (t[61] & ~t[63] & ~t[64]) | (t[61] & ~t[62] & ~t[64]) | (t[61] & ~t[62] & ~t[63]);
  assign t[49] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[4] = ~(t[6] ^ t[27]);
  assign t[50] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[51] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[52] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[53] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[54] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[55] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[56] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[57] = t[97] ^ x[6];
  assign t[58] = t[98] ^ x[3];
  assign t[59] = t[99] ^ x[4];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[100] ^ x[5];
  assign t[61] = t[101] ^ x[11];
  assign t[62] = t[102] ^ x[8];
  assign t[63] = t[103] ^ x[9];
  assign t[64] = t[104] ^ x[10];
  assign t[65] = t[105] ^ x[16];
  assign t[66] = t[106] ^ x[13];
  assign t[67] = t[107] ^ x[14];
  assign t[68] = t[108] ^ x[15];
  assign t[69] = t[109] ^ x[21];
  assign t[6] = ~t[9];
  assign t[70] = t[110] ^ x[18];
  assign t[71] = t[111] ^ x[19];
  assign t[72] = t[112] ^ x[20];
  assign t[73] = t[113] ^ x[26];
  assign t[74] = t[114] ^ x[23];
  assign t[75] = t[115] ^ x[24];
  assign t[76] = t[116] ^ x[25];
  assign t[77] = t[117] ^ x[31];
  assign t[78] = t[118] ^ x[28];
  assign t[79] = t[119] ^ x[29];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[120] ^ x[30];
  assign t[81] = t[121] ^ x[36];
  assign t[82] = t[122] ^ x[33];
  assign t[83] = t[123] ^ x[34];
  assign t[84] = t[124] ^ x[35];
  assign t[85] = t[125] ^ x[41];
  assign t[86] = t[126] ^ x[38];
  assign t[87] = t[127] ^ x[39];
  assign t[88] = t[128] ^ x[40];
  assign t[89] = t[129] ^ x[46];
  assign t[8] = t[12] & t[13];
  assign t[90] = t[130] ^ x[43];
  assign t[91] = t[131] ^ x[44];
  assign t[92] = t[132] ^ x[45];
  assign t[93] = t[133] ^ x[51];
  assign t[94] = t[134] ^ x[48];
  assign t[95] = t[135] ^ x[49];
  assign t[96] = t[136] ^ x[50];
  assign t[97] = (x[2]);
  assign t[98] = (x[2]);
  assign t[99] = (x[2]);
  assign t[9] = ~(t[14] ^ t[28]);
  assign y = (t[0]);
endmodule

module R2ind94(x, y);
 input [51:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[7]);
  assign t[102] = (x[7]);
  assign t[103] = (x[7]);
  assign t[104] = (x[7]);
  assign t[105] = (x[12]);
  assign t[106] = (x[12]);
  assign t[107] = (x[12]);
  assign t[108] = (x[12]);
  assign t[109] = (x[17]);
  assign t[10] = t[29] ^ t[30];
  assign t[110] = (x[17]);
  assign t[111] = (x[17]);
  assign t[112] = (x[17]);
  assign t[113] = (x[22]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[22]);
  assign t[117] = (x[27]);
  assign t[118] = (x[27]);
  assign t[119] = (x[27]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[32]);
  assign t[122] = (x[32]);
  assign t[123] = (x[32]);
  assign t[124] = (x[32]);
  assign t[125] = (x[37]);
  assign t[126] = (x[37]);
  assign t[127] = (x[37]);
  assign t[128] = (x[37]);
  assign t[129] = (x[42]);
  assign t[12] = ~(t[30]);
  assign t[130] = (x[42]);
  assign t[131] = (x[42]);
  assign t[132] = (x[42]);
  assign t[133] = (x[47]);
  assign t[134] = (x[47]);
  assign t[135] = (x[47]);
  assign t[136] = (x[47]);
  assign t[13] = ~(t[31] ^ t[12]);
  assign t[14] = ~t[16];
  assign t[15] = t[31] ^ t[17];
  assign t[16] = ~(t[18]);
  assign t[17] = t[30] ^ t[32];
  assign t[18] = t[19] ^ t[20];
  assign t[19] = t[21] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] & t[24];
  assign t[21] = t[33] ^ t[34];
  assign t[22] = t[23] & t[25];
  assign t[23] = ~(t[34]);
  assign t[24] = ~(t[35] ^ t[23]);
  assign t[25] = t[35] ^ t[26];
  assign t[26] = t[34] ^ t[36];
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~t[4];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = t[47] ^ x[6];
  assign t[38] = t[48] ^ x[11];
  assign t[39] = t[49] ^ x[16];
  assign t[3] = ~(t[5]);
  assign t[40] = t[50] ^ x[21];
  assign t[41] = t[51] ^ x[26];
  assign t[42] = t[52] ^ x[31];
  assign t[43] = t[53] ^ x[36];
  assign t[44] = t[54] ^ x[41];
  assign t[45] = t[55] ^ x[46];
  assign t[46] = t[56] ^ x[51];
  assign t[47] = (~t[57] & t[58] & t[59] & t[60]) | (t[57] & ~t[59] & ~t[60]) | (t[57] & ~t[58] & ~t[60]) | (t[57] & ~t[58] & ~t[59]);
  assign t[48] = (~t[61] & t[62] & t[63] & t[64]) | (t[61] & ~t[63] & ~t[64]) | (t[61] & ~t[62] & ~t[64]) | (t[61] & ~t[62] & ~t[63]);
  assign t[49] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[4] = ~(t[6] ^ t[27]);
  assign t[50] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[51] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[52] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[53] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[54] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[55] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[56] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[57] = t[97] ^ x[6];
  assign t[58] = t[98] ^ x[3];
  assign t[59] = t[99] ^ x[4];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[100] ^ x[5];
  assign t[61] = t[101] ^ x[11];
  assign t[62] = t[102] ^ x[8];
  assign t[63] = t[103] ^ x[9];
  assign t[64] = t[104] ^ x[10];
  assign t[65] = t[105] ^ x[16];
  assign t[66] = t[106] ^ x[13];
  assign t[67] = t[107] ^ x[14];
  assign t[68] = t[108] ^ x[15];
  assign t[69] = t[109] ^ x[21];
  assign t[6] = ~t[9];
  assign t[70] = t[110] ^ x[18];
  assign t[71] = t[111] ^ x[19];
  assign t[72] = t[112] ^ x[20];
  assign t[73] = t[113] ^ x[26];
  assign t[74] = t[114] ^ x[23];
  assign t[75] = t[115] ^ x[24];
  assign t[76] = t[116] ^ x[25];
  assign t[77] = t[117] ^ x[31];
  assign t[78] = t[118] ^ x[28];
  assign t[79] = t[119] ^ x[29];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[120] ^ x[30];
  assign t[81] = t[121] ^ x[36];
  assign t[82] = t[122] ^ x[33];
  assign t[83] = t[123] ^ x[34];
  assign t[84] = t[124] ^ x[35];
  assign t[85] = t[125] ^ x[41];
  assign t[86] = t[126] ^ x[38];
  assign t[87] = t[127] ^ x[39];
  assign t[88] = t[128] ^ x[40];
  assign t[89] = t[129] ^ x[46];
  assign t[8] = t[12] & t[13];
  assign t[90] = t[130] ^ x[43];
  assign t[91] = t[131] ^ x[44];
  assign t[92] = t[132] ^ x[45];
  assign t[93] = t[133] ^ x[51];
  assign t[94] = t[134] ^ x[48];
  assign t[95] = t[135] ^ x[49];
  assign t[96] = t[136] ^ x[50];
  assign t[97] = (x[2]);
  assign t[98] = (x[2]);
  assign t[99] = (x[2]);
  assign t[9] = ~(t[14] ^ t[28]);
  assign y = (t[0]);
endmodule

module R2ind95(x, y);
 input [51:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[7]);
  assign t[102] = (x[7]);
  assign t[103] = (x[7]);
  assign t[104] = (x[7]);
  assign t[105] = (x[12]);
  assign t[106] = (x[12]);
  assign t[107] = (x[12]);
  assign t[108] = (x[12]);
  assign t[109] = (x[17]);
  assign t[10] = t[29] ^ t[30];
  assign t[110] = (x[17]);
  assign t[111] = (x[17]);
  assign t[112] = (x[17]);
  assign t[113] = (x[22]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[22]);
  assign t[117] = (x[27]);
  assign t[118] = (x[27]);
  assign t[119] = (x[27]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[32]);
  assign t[122] = (x[32]);
  assign t[123] = (x[32]);
  assign t[124] = (x[32]);
  assign t[125] = (x[37]);
  assign t[126] = (x[37]);
  assign t[127] = (x[37]);
  assign t[128] = (x[37]);
  assign t[129] = (x[42]);
  assign t[12] = ~(t[30]);
  assign t[130] = (x[42]);
  assign t[131] = (x[42]);
  assign t[132] = (x[42]);
  assign t[133] = (x[47]);
  assign t[134] = (x[47]);
  assign t[135] = (x[47]);
  assign t[136] = (x[47]);
  assign t[13] = ~(t[31] ^ t[12]);
  assign t[14] = ~t[16];
  assign t[15] = t[31] ^ t[17];
  assign t[16] = ~(t[18]);
  assign t[17] = t[30] ^ t[32];
  assign t[18] = t[19] ^ t[20];
  assign t[19] = t[21] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] & t[24];
  assign t[21] = t[33] ^ t[34];
  assign t[22] = t[23] & t[25];
  assign t[23] = ~(t[34]);
  assign t[24] = ~(t[35] ^ t[23]);
  assign t[25] = t[35] ^ t[26];
  assign t[26] = t[34] ^ t[36];
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~t[4];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = t[47] ^ x[6];
  assign t[38] = t[48] ^ x[11];
  assign t[39] = t[49] ^ x[16];
  assign t[3] = ~(t[5]);
  assign t[40] = t[50] ^ x[21];
  assign t[41] = t[51] ^ x[26];
  assign t[42] = t[52] ^ x[31];
  assign t[43] = t[53] ^ x[36];
  assign t[44] = t[54] ^ x[41];
  assign t[45] = t[55] ^ x[46];
  assign t[46] = t[56] ^ x[51];
  assign t[47] = (~t[57] & t[58] & t[59] & t[60]) | (t[57] & ~t[59] & ~t[60]) | (t[57] & ~t[58] & ~t[60]) | (t[57] & ~t[58] & ~t[59]);
  assign t[48] = (~t[61] & t[62] & t[63] & t[64]) | (t[61] & ~t[63] & ~t[64]) | (t[61] & ~t[62] & ~t[64]) | (t[61] & ~t[62] & ~t[63]);
  assign t[49] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[4] = ~(t[6] ^ t[27]);
  assign t[50] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[51] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[52] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[53] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[54] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[55] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[56] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[57] = t[97] ^ x[6];
  assign t[58] = t[98] ^ x[3];
  assign t[59] = t[99] ^ x[4];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[100] ^ x[5];
  assign t[61] = t[101] ^ x[11];
  assign t[62] = t[102] ^ x[8];
  assign t[63] = t[103] ^ x[9];
  assign t[64] = t[104] ^ x[10];
  assign t[65] = t[105] ^ x[16];
  assign t[66] = t[106] ^ x[13];
  assign t[67] = t[107] ^ x[14];
  assign t[68] = t[108] ^ x[15];
  assign t[69] = t[109] ^ x[21];
  assign t[6] = ~t[9];
  assign t[70] = t[110] ^ x[18];
  assign t[71] = t[111] ^ x[19];
  assign t[72] = t[112] ^ x[20];
  assign t[73] = t[113] ^ x[26];
  assign t[74] = t[114] ^ x[23];
  assign t[75] = t[115] ^ x[24];
  assign t[76] = t[116] ^ x[25];
  assign t[77] = t[117] ^ x[31];
  assign t[78] = t[118] ^ x[28];
  assign t[79] = t[119] ^ x[29];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[120] ^ x[30];
  assign t[81] = t[121] ^ x[36];
  assign t[82] = t[122] ^ x[33];
  assign t[83] = t[123] ^ x[34];
  assign t[84] = t[124] ^ x[35];
  assign t[85] = t[125] ^ x[41];
  assign t[86] = t[126] ^ x[38];
  assign t[87] = t[127] ^ x[39];
  assign t[88] = t[128] ^ x[40];
  assign t[89] = t[129] ^ x[46];
  assign t[8] = t[12] & t[13];
  assign t[90] = t[130] ^ x[43];
  assign t[91] = t[131] ^ x[44];
  assign t[92] = t[132] ^ x[45];
  assign t[93] = t[133] ^ x[51];
  assign t[94] = t[134] ^ x[48];
  assign t[95] = t[135] ^ x[49];
  assign t[96] = t[136] ^ x[50];
  assign t[97] = (x[2]);
  assign t[98] = (x[2]);
  assign t[99] = (x[2]);
  assign t[9] = ~(t[14] ^ t[28]);
  assign y = (t[0]);
endmodule

module R2ind96(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind97(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind98(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind99(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind100(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[38] ^ t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind101(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[38] ^ t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind102(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[38] ^ t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind103(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[38] ^ t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind104(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind105(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind106(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind107(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind108(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind109(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind110(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind111(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind112(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind113(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind114(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind115(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind116(x, y);
 input [46:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[136] ^ x[45];
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[2]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[7]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[17];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[12]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[17]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[18] & t[19];
  assign t[120] = (x[22]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[27]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[32]);
  assign t[129] = (x[37]);
  assign t[12] = t[20] ^ t[11];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[37]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[136] = (x[42]);
  assign t[13] = t[39] ^ t[18];
  assign t[14] = t[21] ^ t[22];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[40] ^ t[41];
  assign t[17] = t[18] & t[25];
  assign t[18] = ~(t[41]);
  assign t[19] = ~(t[39] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[39] & t[26];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[42] ^ t[29];
  assign t[25] = t[39] ^ t[32];
  assign t[26] = t[33] ^ t[17];
  assign t[27] = t[43] ^ t[44];
  assign t[28] = t[29] & t[34];
  assign t[29] = ~(t[44]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[42] ^ t[29]);
  assign t[31] = t[42] & t[35];
  assign t[32] = t[41] ^ t[45];
  assign t[33] = t[39] ^ t[16];
  assign t[34] = t[42] ^ t[36];
  assign t[35] = t[37] ^ t[28];
  assign t[36] = t[44] ^ t[46];
  assign t[37] = t[42] ^ t[27];
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = (t[55]);
  assign t[47] = t[56] ^ x[6];
  assign t[48] = t[57] ^ x[11];
  assign t[49] = t[58] ^ x[16];
  assign t[4] = ~(t[6] ^ t[38]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[26];
  assign t[52] = t[61] ^ x[31];
  assign t[53] = t[62] ^ x[36];
  assign t[54] = t[63] ^ x[41];
  assign t[55] = t[64] ^ x[46];
  assign t[56] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[57] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[58] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[59] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[60] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[61] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[62] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[63] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[64] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[65] = t[101] ^ x[6];
  assign t[66] = t[102] ^ x[3];
  assign t[67] = t[103] ^ x[4];
  assign t[68] = t[104] ^ x[5];
  assign t[69] = t[105] ^ x[11];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[8];
  assign t[71] = t[107] ^ x[9];
  assign t[72] = t[108] ^ x[10];
  assign t[73] = t[109] ^ x[16];
  assign t[74] = t[110] ^ x[13];
  assign t[75] = t[111] ^ x[14];
  assign t[76] = t[112] ^ x[15];
  assign t[77] = t[113] ^ x[21];
  assign t[78] = t[114] ^ x[18];
  assign t[79] = t[115] ^ x[19];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[20];
  assign t[81] = t[117] ^ x[26];
  assign t[82] = t[118] ^ x[23];
  assign t[83] = t[119] ^ x[24];
  assign t[84] = t[120] ^ x[25];
  assign t[85] = t[121] ^ x[31];
  assign t[86] = t[122] ^ x[28];
  assign t[87] = t[123] ^ x[29];
  assign t[88] = t[124] ^ x[30];
  assign t[89] = t[125] ^ x[36];
  assign t[8] = t[12] ^ t[13];
  assign t[90] = t[126] ^ x[33];
  assign t[91] = t[127] ^ x[34];
  assign t[92] = t[128] ^ x[35];
  assign t[93] = t[129] ^ x[41];
  assign t[94] = t[130] ^ x[38];
  assign t[95] = t[131] ^ x[39];
  assign t[96] = t[132] ^ x[40];
  assign t[97] = t[133] ^ x[46];
  assign t[98] = t[134] ^ x[43];
  assign t[99] = t[135] ^ x[44];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = (t[0]);
endmodule

module R2ind117(x, y);
 input [46:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[136] ^ x[45];
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[2]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[7]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[17];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[12]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[17]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[18] & t[19];
  assign t[120] = (x[22]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[27]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[32]);
  assign t[129] = (x[37]);
  assign t[12] = t[20] ^ t[11];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[37]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[136] = (x[42]);
  assign t[13] = t[39] ^ t[18];
  assign t[14] = t[21] ^ t[22];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[40] ^ t[41];
  assign t[17] = t[18] & t[25];
  assign t[18] = ~(t[41]);
  assign t[19] = ~(t[39] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[39] & t[26];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[42] ^ t[29];
  assign t[25] = t[39] ^ t[32];
  assign t[26] = t[33] ^ t[17];
  assign t[27] = t[43] ^ t[44];
  assign t[28] = t[29] & t[34];
  assign t[29] = ~(t[44]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[42] ^ t[29]);
  assign t[31] = t[42] & t[35];
  assign t[32] = t[41] ^ t[45];
  assign t[33] = t[39] ^ t[16];
  assign t[34] = t[42] ^ t[36];
  assign t[35] = t[37] ^ t[28];
  assign t[36] = t[44] ^ t[46];
  assign t[37] = t[42] ^ t[27];
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = (t[55]);
  assign t[47] = t[56] ^ x[6];
  assign t[48] = t[57] ^ x[11];
  assign t[49] = t[58] ^ x[16];
  assign t[4] = ~(t[6] ^ t[38]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[26];
  assign t[52] = t[61] ^ x[31];
  assign t[53] = t[62] ^ x[36];
  assign t[54] = t[63] ^ x[41];
  assign t[55] = t[64] ^ x[46];
  assign t[56] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[57] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[58] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[59] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[60] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[61] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[62] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[63] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[64] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[65] = t[101] ^ x[6];
  assign t[66] = t[102] ^ x[3];
  assign t[67] = t[103] ^ x[4];
  assign t[68] = t[104] ^ x[5];
  assign t[69] = t[105] ^ x[11];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[8];
  assign t[71] = t[107] ^ x[9];
  assign t[72] = t[108] ^ x[10];
  assign t[73] = t[109] ^ x[16];
  assign t[74] = t[110] ^ x[13];
  assign t[75] = t[111] ^ x[14];
  assign t[76] = t[112] ^ x[15];
  assign t[77] = t[113] ^ x[21];
  assign t[78] = t[114] ^ x[18];
  assign t[79] = t[115] ^ x[19];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[20];
  assign t[81] = t[117] ^ x[26];
  assign t[82] = t[118] ^ x[23];
  assign t[83] = t[119] ^ x[24];
  assign t[84] = t[120] ^ x[25];
  assign t[85] = t[121] ^ x[31];
  assign t[86] = t[122] ^ x[28];
  assign t[87] = t[123] ^ x[29];
  assign t[88] = t[124] ^ x[30];
  assign t[89] = t[125] ^ x[36];
  assign t[8] = t[12] ^ t[13];
  assign t[90] = t[126] ^ x[33];
  assign t[91] = t[127] ^ x[34];
  assign t[92] = t[128] ^ x[35];
  assign t[93] = t[129] ^ x[41];
  assign t[94] = t[130] ^ x[38];
  assign t[95] = t[131] ^ x[39];
  assign t[96] = t[132] ^ x[40];
  assign t[97] = t[133] ^ x[46];
  assign t[98] = t[134] ^ x[43];
  assign t[99] = t[135] ^ x[44];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = (t[0]);
endmodule

module R2ind118(x, y);
 input [46:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[136] ^ x[45];
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[2]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[7]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[17];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[12]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[17]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[18] & t[19];
  assign t[120] = (x[22]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[27]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[32]);
  assign t[129] = (x[37]);
  assign t[12] = t[20] ^ t[11];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[37]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[136] = (x[42]);
  assign t[13] = t[39] ^ t[18];
  assign t[14] = t[21] ^ t[22];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[40] ^ t[41];
  assign t[17] = t[18] & t[25];
  assign t[18] = ~(t[41]);
  assign t[19] = ~(t[39] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[39] & t[26];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[42] ^ t[29];
  assign t[25] = t[39] ^ t[32];
  assign t[26] = t[33] ^ t[17];
  assign t[27] = t[43] ^ t[44];
  assign t[28] = t[29] & t[34];
  assign t[29] = ~(t[44]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[42] ^ t[29]);
  assign t[31] = t[42] & t[35];
  assign t[32] = t[41] ^ t[45];
  assign t[33] = t[39] ^ t[16];
  assign t[34] = t[42] ^ t[36];
  assign t[35] = t[37] ^ t[28];
  assign t[36] = t[44] ^ t[46];
  assign t[37] = t[42] ^ t[27];
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = (t[55]);
  assign t[47] = t[56] ^ x[6];
  assign t[48] = t[57] ^ x[11];
  assign t[49] = t[58] ^ x[16];
  assign t[4] = ~(t[6] ^ t[38]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[26];
  assign t[52] = t[61] ^ x[31];
  assign t[53] = t[62] ^ x[36];
  assign t[54] = t[63] ^ x[41];
  assign t[55] = t[64] ^ x[46];
  assign t[56] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[57] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[58] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[59] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[60] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[61] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[62] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[63] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[64] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[65] = t[101] ^ x[6];
  assign t[66] = t[102] ^ x[3];
  assign t[67] = t[103] ^ x[4];
  assign t[68] = t[104] ^ x[5];
  assign t[69] = t[105] ^ x[11];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[8];
  assign t[71] = t[107] ^ x[9];
  assign t[72] = t[108] ^ x[10];
  assign t[73] = t[109] ^ x[16];
  assign t[74] = t[110] ^ x[13];
  assign t[75] = t[111] ^ x[14];
  assign t[76] = t[112] ^ x[15];
  assign t[77] = t[113] ^ x[21];
  assign t[78] = t[114] ^ x[18];
  assign t[79] = t[115] ^ x[19];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[20];
  assign t[81] = t[117] ^ x[26];
  assign t[82] = t[118] ^ x[23];
  assign t[83] = t[119] ^ x[24];
  assign t[84] = t[120] ^ x[25];
  assign t[85] = t[121] ^ x[31];
  assign t[86] = t[122] ^ x[28];
  assign t[87] = t[123] ^ x[29];
  assign t[88] = t[124] ^ x[30];
  assign t[89] = t[125] ^ x[36];
  assign t[8] = t[12] ^ t[13];
  assign t[90] = t[126] ^ x[33];
  assign t[91] = t[127] ^ x[34];
  assign t[92] = t[128] ^ x[35];
  assign t[93] = t[129] ^ x[41];
  assign t[94] = t[130] ^ x[38];
  assign t[95] = t[131] ^ x[39];
  assign t[96] = t[132] ^ x[40];
  assign t[97] = t[133] ^ x[46];
  assign t[98] = t[134] ^ x[43];
  assign t[99] = t[135] ^ x[44];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = (t[0]);
endmodule

module R2ind119(x, y);
 input [46:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[136] ^ x[45];
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[2]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[7]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[17];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[12]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[17]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[18] & t[19];
  assign t[120] = (x[22]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[27]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[32]);
  assign t[129] = (x[37]);
  assign t[12] = t[20] ^ t[11];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[37]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[136] = (x[42]);
  assign t[13] = t[39] ^ t[18];
  assign t[14] = t[21] ^ t[22];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[40] ^ t[41];
  assign t[17] = t[18] & t[25];
  assign t[18] = ~(t[41]);
  assign t[19] = ~(t[39] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[39] & t[26];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[42] ^ t[29];
  assign t[25] = t[39] ^ t[32];
  assign t[26] = t[33] ^ t[17];
  assign t[27] = t[43] ^ t[44];
  assign t[28] = t[29] & t[34];
  assign t[29] = ~(t[44]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[42] ^ t[29]);
  assign t[31] = t[42] & t[35];
  assign t[32] = t[41] ^ t[45];
  assign t[33] = t[39] ^ t[16];
  assign t[34] = t[42] ^ t[36];
  assign t[35] = t[37] ^ t[28];
  assign t[36] = t[44] ^ t[46];
  assign t[37] = t[42] ^ t[27];
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = (t[55]);
  assign t[47] = t[56] ^ x[6];
  assign t[48] = t[57] ^ x[11];
  assign t[49] = t[58] ^ x[16];
  assign t[4] = ~(t[6] ^ t[38]);
  assign t[50] = t[59] ^ x[21];
  assign t[51] = t[60] ^ x[26];
  assign t[52] = t[61] ^ x[31];
  assign t[53] = t[62] ^ x[36];
  assign t[54] = t[63] ^ x[41];
  assign t[55] = t[64] ^ x[46];
  assign t[56] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[57] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[58] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[59] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[60] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[61] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[62] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[63] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[64] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[65] = t[101] ^ x[6];
  assign t[66] = t[102] ^ x[3];
  assign t[67] = t[103] ^ x[4];
  assign t[68] = t[104] ^ x[5];
  assign t[69] = t[105] ^ x[11];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[8];
  assign t[71] = t[107] ^ x[9];
  assign t[72] = t[108] ^ x[10];
  assign t[73] = t[109] ^ x[16];
  assign t[74] = t[110] ^ x[13];
  assign t[75] = t[111] ^ x[14];
  assign t[76] = t[112] ^ x[15];
  assign t[77] = t[113] ^ x[21];
  assign t[78] = t[114] ^ x[18];
  assign t[79] = t[115] ^ x[19];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[20];
  assign t[81] = t[117] ^ x[26];
  assign t[82] = t[118] ^ x[23];
  assign t[83] = t[119] ^ x[24];
  assign t[84] = t[120] ^ x[25];
  assign t[85] = t[121] ^ x[31];
  assign t[86] = t[122] ^ x[28];
  assign t[87] = t[123] ^ x[29];
  assign t[88] = t[124] ^ x[30];
  assign t[89] = t[125] ^ x[36];
  assign t[8] = t[12] ^ t[13];
  assign t[90] = t[126] ^ x[33];
  assign t[91] = t[127] ^ x[34];
  assign t[92] = t[128] ^ x[35];
  assign t[93] = t[129] ^ x[41];
  assign t[94] = t[130] ^ x[38];
  assign t[95] = t[131] ^ x[39];
  assign t[96] = t[132] ^ x[40];
  assign t[97] = t[133] ^ x[46];
  assign t[98] = t[134] ^ x[43];
  assign t[99] = t[135] ^ x[44];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = (t[0]);
endmodule

module R2ind120(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind121(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind122(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind123(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind124(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind125(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind126(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind127(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind128(x, y);
 input [51:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ^ x[40];
  assign t[101] = t[141] ^ x[46];
  assign t[102] = t[142] ^ x[43];
  assign t[103] = t[143] ^ x[44];
  assign t[104] = t[144] ^ x[45];
  assign t[105] = t[145] ^ x[51];
  assign t[106] = t[146] ^ x[48];
  assign t[107] = t[147] ^ x[49];
  assign t[108] = t[148] ^ x[50];
  assign t[109] = (x[2]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[2]);
  assign t[111] = (x[2]);
  assign t[112] = (x[2]);
  assign t[113] = (x[7]);
  assign t[114] = (x[7]);
  assign t[115] = (x[7]);
  assign t[116] = (x[7]);
  assign t[117] = (x[12]);
  assign t[118] = (x[12]);
  assign t[119] = (x[12]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[12]);
  assign t[121] = (x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[17]);
  assign t[124] = (x[17]);
  assign t[125] = (x[22]);
  assign t[126] = (x[22]);
  assign t[127] = (x[22]);
  assign t[128] = (x[22]);
  assign t[129] = (x[27]);
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[130] = (x[27]);
  assign t[131] = (x[27]);
  assign t[132] = (x[27]);
  assign t[133] = (x[32]);
  assign t[134] = (x[32]);
  assign t[135] = (x[32]);
  assign t[136] = (x[32]);
  assign t[137] = (x[37]);
  assign t[138] = (x[37]);
  assign t[139] = (x[37]);
  assign t[13] = t[19] ^ t[20];
  assign t[140] = (x[37]);
  assign t[141] = (x[42]);
  assign t[142] = (x[42]);
  assign t[143] = (x[42]);
  assign t[144] = (x[42]);
  assign t[145] = (x[47]);
  assign t[146] = (x[47]);
  assign t[147] = (x[47]);
  assign t[148] = (x[47]);
  assign t[14] = ~(t[42]);
  assign t[15] = ~(t[40] ^ t[14]);
  assign t[16] = t[43] ^ t[42];
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[18] = ~t[22];
  assign t[19] = t[40] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[40] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[42] ^ t[44];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[45] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[45] ^ t[31]);
  assign t[33] = t[47] ^ t[46];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[45] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[45] ^ t[38];
  assign t[38] = t[46] ^ t[48];
  assign t[39] = (t[49]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[6];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[11];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[21];
  assign t[53] = t[63] ^ x[26];
  assign t[54] = t[64] ^ x[31];
  assign t[55] = t[65] ^ x[36];
  assign t[56] = t[66] ^ x[41];
  assign t[57] = t[67] ^ x[46];
  assign t[58] = t[68] ^ x[51];
  assign t[59] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[61] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[62] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[63] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[64] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[65] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[66] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[67] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[68] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[69] = t[109] ^ x[6];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[110] ^ x[3];
  assign t[71] = t[111] ^ x[4];
  assign t[72] = t[112] ^ x[5];
  assign t[73] = t[113] ^ x[11];
  assign t[74] = t[114] ^ x[8];
  assign t[75] = t[115] ^ x[9];
  assign t[76] = t[116] ^ x[10];
  assign t[77] = t[117] ^ x[16];
  assign t[78] = t[118] ^ x[13];
  assign t[79] = t[119] ^ x[14];
  assign t[7] = ~t[12];
  assign t[80] = t[120] ^ x[15];
  assign t[81] = t[121] ^ x[21];
  assign t[82] = t[122] ^ x[18];
  assign t[83] = t[123] ^ x[19];
  assign t[84] = t[124] ^ x[20];
  assign t[85] = t[125] ^ x[26];
  assign t[86] = t[126] ^ x[23];
  assign t[87] = t[127] ^ x[24];
  assign t[88] = t[128] ^ x[25];
  assign t[89] = t[129] ^ x[31];
  assign t[8] = t[40] & t[13];
  assign t[90] = t[130] ^ x[28];
  assign t[91] = t[131] ^ x[29];
  assign t[92] = t[132] ^ x[30];
  assign t[93] = t[133] ^ x[36];
  assign t[94] = t[134] ^ x[33];
  assign t[95] = t[135] ^ x[34];
  assign t[96] = t[136] ^ x[35];
  assign t[97] = t[137] ^ x[41];
  assign t[98] = t[138] ^ x[38];
  assign t[99] = t[139] ^ x[39];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind129(x, y);
 input [51:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ^ x[40];
  assign t[101] = t[141] ^ x[46];
  assign t[102] = t[142] ^ x[43];
  assign t[103] = t[143] ^ x[44];
  assign t[104] = t[144] ^ x[45];
  assign t[105] = t[145] ^ x[51];
  assign t[106] = t[146] ^ x[48];
  assign t[107] = t[147] ^ x[49];
  assign t[108] = t[148] ^ x[50];
  assign t[109] = (x[2]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[2]);
  assign t[111] = (x[2]);
  assign t[112] = (x[2]);
  assign t[113] = (x[7]);
  assign t[114] = (x[7]);
  assign t[115] = (x[7]);
  assign t[116] = (x[7]);
  assign t[117] = (x[12]);
  assign t[118] = (x[12]);
  assign t[119] = (x[12]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[12]);
  assign t[121] = (x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[17]);
  assign t[124] = (x[17]);
  assign t[125] = (x[22]);
  assign t[126] = (x[22]);
  assign t[127] = (x[22]);
  assign t[128] = (x[22]);
  assign t[129] = (x[27]);
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[130] = (x[27]);
  assign t[131] = (x[27]);
  assign t[132] = (x[27]);
  assign t[133] = (x[32]);
  assign t[134] = (x[32]);
  assign t[135] = (x[32]);
  assign t[136] = (x[32]);
  assign t[137] = (x[37]);
  assign t[138] = (x[37]);
  assign t[139] = (x[37]);
  assign t[13] = t[19] ^ t[20];
  assign t[140] = (x[37]);
  assign t[141] = (x[42]);
  assign t[142] = (x[42]);
  assign t[143] = (x[42]);
  assign t[144] = (x[42]);
  assign t[145] = (x[47]);
  assign t[146] = (x[47]);
  assign t[147] = (x[47]);
  assign t[148] = (x[47]);
  assign t[14] = ~(t[42]);
  assign t[15] = ~(t[40] ^ t[14]);
  assign t[16] = t[43] ^ t[42];
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[18] = ~t[22];
  assign t[19] = t[40] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[40] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[42] ^ t[44];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[45] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[45] ^ t[31]);
  assign t[33] = t[47] ^ t[46];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[45] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[45] ^ t[38];
  assign t[38] = t[46] ^ t[48];
  assign t[39] = (t[49]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[6];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[11];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[21];
  assign t[53] = t[63] ^ x[26];
  assign t[54] = t[64] ^ x[31];
  assign t[55] = t[65] ^ x[36];
  assign t[56] = t[66] ^ x[41];
  assign t[57] = t[67] ^ x[46];
  assign t[58] = t[68] ^ x[51];
  assign t[59] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[61] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[62] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[63] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[64] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[65] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[66] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[67] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[68] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[69] = t[109] ^ x[6];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[110] ^ x[3];
  assign t[71] = t[111] ^ x[4];
  assign t[72] = t[112] ^ x[5];
  assign t[73] = t[113] ^ x[11];
  assign t[74] = t[114] ^ x[8];
  assign t[75] = t[115] ^ x[9];
  assign t[76] = t[116] ^ x[10];
  assign t[77] = t[117] ^ x[16];
  assign t[78] = t[118] ^ x[13];
  assign t[79] = t[119] ^ x[14];
  assign t[7] = ~t[12];
  assign t[80] = t[120] ^ x[15];
  assign t[81] = t[121] ^ x[21];
  assign t[82] = t[122] ^ x[18];
  assign t[83] = t[123] ^ x[19];
  assign t[84] = t[124] ^ x[20];
  assign t[85] = t[125] ^ x[26];
  assign t[86] = t[126] ^ x[23];
  assign t[87] = t[127] ^ x[24];
  assign t[88] = t[128] ^ x[25];
  assign t[89] = t[129] ^ x[31];
  assign t[8] = t[40] & t[13];
  assign t[90] = t[130] ^ x[28];
  assign t[91] = t[131] ^ x[29];
  assign t[92] = t[132] ^ x[30];
  assign t[93] = t[133] ^ x[36];
  assign t[94] = t[134] ^ x[33];
  assign t[95] = t[135] ^ x[34];
  assign t[96] = t[136] ^ x[35];
  assign t[97] = t[137] ^ x[41];
  assign t[98] = t[138] ^ x[38];
  assign t[99] = t[139] ^ x[39];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind130(x, y);
 input [51:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ^ x[40];
  assign t[101] = t[141] ^ x[46];
  assign t[102] = t[142] ^ x[43];
  assign t[103] = t[143] ^ x[44];
  assign t[104] = t[144] ^ x[45];
  assign t[105] = t[145] ^ x[51];
  assign t[106] = t[146] ^ x[48];
  assign t[107] = t[147] ^ x[49];
  assign t[108] = t[148] ^ x[50];
  assign t[109] = (x[2]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[2]);
  assign t[111] = (x[2]);
  assign t[112] = (x[2]);
  assign t[113] = (x[7]);
  assign t[114] = (x[7]);
  assign t[115] = (x[7]);
  assign t[116] = (x[7]);
  assign t[117] = (x[12]);
  assign t[118] = (x[12]);
  assign t[119] = (x[12]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[12]);
  assign t[121] = (x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[17]);
  assign t[124] = (x[17]);
  assign t[125] = (x[22]);
  assign t[126] = (x[22]);
  assign t[127] = (x[22]);
  assign t[128] = (x[22]);
  assign t[129] = (x[27]);
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[130] = (x[27]);
  assign t[131] = (x[27]);
  assign t[132] = (x[27]);
  assign t[133] = (x[32]);
  assign t[134] = (x[32]);
  assign t[135] = (x[32]);
  assign t[136] = (x[32]);
  assign t[137] = (x[37]);
  assign t[138] = (x[37]);
  assign t[139] = (x[37]);
  assign t[13] = t[19] ^ t[20];
  assign t[140] = (x[37]);
  assign t[141] = (x[42]);
  assign t[142] = (x[42]);
  assign t[143] = (x[42]);
  assign t[144] = (x[42]);
  assign t[145] = (x[47]);
  assign t[146] = (x[47]);
  assign t[147] = (x[47]);
  assign t[148] = (x[47]);
  assign t[14] = ~(t[42]);
  assign t[15] = ~(t[40] ^ t[14]);
  assign t[16] = t[43] ^ t[42];
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[18] = ~t[22];
  assign t[19] = t[40] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[40] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[42] ^ t[44];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[45] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[45] ^ t[31]);
  assign t[33] = t[47] ^ t[46];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[45] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[45] ^ t[38];
  assign t[38] = t[46] ^ t[48];
  assign t[39] = (t[49]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[6];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[11];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[21];
  assign t[53] = t[63] ^ x[26];
  assign t[54] = t[64] ^ x[31];
  assign t[55] = t[65] ^ x[36];
  assign t[56] = t[66] ^ x[41];
  assign t[57] = t[67] ^ x[46];
  assign t[58] = t[68] ^ x[51];
  assign t[59] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[61] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[62] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[63] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[64] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[65] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[66] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[67] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[68] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[69] = t[109] ^ x[6];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[110] ^ x[3];
  assign t[71] = t[111] ^ x[4];
  assign t[72] = t[112] ^ x[5];
  assign t[73] = t[113] ^ x[11];
  assign t[74] = t[114] ^ x[8];
  assign t[75] = t[115] ^ x[9];
  assign t[76] = t[116] ^ x[10];
  assign t[77] = t[117] ^ x[16];
  assign t[78] = t[118] ^ x[13];
  assign t[79] = t[119] ^ x[14];
  assign t[7] = ~t[12];
  assign t[80] = t[120] ^ x[15];
  assign t[81] = t[121] ^ x[21];
  assign t[82] = t[122] ^ x[18];
  assign t[83] = t[123] ^ x[19];
  assign t[84] = t[124] ^ x[20];
  assign t[85] = t[125] ^ x[26];
  assign t[86] = t[126] ^ x[23];
  assign t[87] = t[127] ^ x[24];
  assign t[88] = t[128] ^ x[25];
  assign t[89] = t[129] ^ x[31];
  assign t[8] = t[40] & t[13];
  assign t[90] = t[130] ^ x[28];
  assign t[91] = t[131] ^ x[29];
  assign t[92] = t[132] ^ x[30];
  assign t[93] = t[133] ^ x[36];
  assign t[94] = t[134] ^ x[33];
  assign t[95] = t[135] ^ x[34];
  assign t[96] = t[136] ^ x[35];
  assign t[97] = t[137] ^ x[41];
  assign t[98] = t[138] ^ x[38];
  assign t[99] = t[139] ^ x[39];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind131(x, y);
 input [51:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ^ x[40];
  assign t[101] = t[141] ^ x[46];
  assign t[102] = t[142] ^ x[43];
  assign t[103] = t[143] ^ x[44];
  assign t[104] = t[144] ^ x[45];
  assign t[105] = t[145] ^ x[51];
  assign t[106] = t[146] ^ x[48];
  assign t[107] = t[147] ^ x[49];
  assign t[108] = t[148] ^ x[50];
  assign t[109] = (x[2]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[2]);
  assign t[111] = (x[2]);
  assign t[112] = (x[2]);
  assign t[113] = (x[7]);
  assign t[114] = (x[7]);
  assign t[115] = (x[7]);
  assign t[116] = (x[7]);
  assign t[117] = (x[12]);
  assign t[118] = (x[12]);
  assign t[119] = (x[12]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[12]);
  assign t[121] = (x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[17]);
  assign t[124] = (x[17]);
  assign t[125] = (x[22]);
  assign t[126] = (x[22]);
  assign t[127] = (x[22]);
  assign t[128] = (x[22]);
  assign t[129] = (x[27]);
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[130] = (x[27]);
  assign t[131] = (x[27]);
  assign t[132] = (x[27]);
  assign t[133] = (x[32]);
  assign t[134] = (x[32]);
  assign t[135] = (x[32]);
  assign t[136] = (x[32]);
  assign t[137] = (x[37]);
  assign t[138] = (x[37]);
  assign t[139] = (x[37]);
  assign t[13] = t[19] ^ t[20];
  assign t[140] = (x[37]);
  assign t[141] = (x[42]);
  assign t[142] = (x[42]);
  assign t[143] = (x[42]);
  assign t[144] = (x[42]);
  assign t[145] = (x[47]);
  assign t[146] = (x[47]);
  assign t[147] = (x[47]);
  assign t[148] = (x[47]);
  assign t[14] = ~(t[42]);
  assign t[15] = ~(t[40] ^ t[14]);
  assign t[16] = t[43] ^ t[42];
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[18] = ~t[22];
  assign t[19] = t[40] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[40] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[42] ^ t[44];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[45] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[45] ^ t[31]);
  assign t[33] = t[47] ^ t[46];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[45] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[45] ^ t[38];
  assign t[38] = t[46] ^ t[48];
  assign t[39] = (t[49]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[6];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[11];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[21];
  assign t[53] = t[63] ^ x[26];
  assign t[54] = t[64] ^ x[31];
  assign t[55] = t[65] ^ x[36];
  assign t[56] = t[66] ^ x[41];
  assign t[57] = t[67] ^ x[46];
  assign t[58] = t[68] ^ x[51];
  assign t[59] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[61] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[62] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[63] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[64] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[65] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[66] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[67] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[68] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[69] = t[109] ^ x[6];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[110] ^ x[3];
  assign t[71] = t[111] ^ x[4];
  assign t[72] = t[112] ^ x[5];
  assign t[73] = t[113] ^ x[11];
  assign t[74] = t[114] ^ x[8];
  assign t[75] = t[115] ^ x[9];
  assign t[76] = t[116] ^ x[10];
  assign t[77] = t[117] ^ x[16];
  assign t[78] = t[118] ^ x[13];
  assign t[79] = t[119] ^ x[14];
  assign t[7] = ~t[12];
  assign t[80] = t[120] ^ x[15];
  assign t[81] = t[121] ^ x[21];
  assign t[82] = t[122] ^ x[18];
  assign t[83] = t[123] ^ x[19];
  assign t[84] = t[124] ^ x[20];
  assign t[85] = t[125] ^ x[26];
  assign t[86] = t[126] ^ x[23];
  assign t[87] = t[127] ^ x[24];
  assign t[88] = t[128] ^ x[25];
  assign t[89] = t[129] ^ x[31];
  assign t[8] = t[40] & t[13];
  assign t[90] = t[130] ^ x[28];
  assign t[91] = t[131] ^ x[29];
  assign t[92] = t[132] ^ x[30];
  assign t[93] = t[133] ^ x[36];
  assign t[94] = t[134] ^ x[33];
  assign t[95] = t[135] ^ x[34];
  assign t[96] = t[136] ^ x[35];
  assign t[97] = t[137] ^ x[41];
  assign t[98] = t[138] ^ x[38];
  assign t[99] = t[139] ^ x[39];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind132(x, y);
 input [51:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ^ x[40];
  assign t[101] = t[141] ^ x[46];
  assign t[102] = t[142] ^ x[43];
  assign t[103] = t[143] ^ x[44];
  assign t[104] = t[144] ^ x[45];
  assign t[105] = t[145] ^ x[51];
  assign t[106] = t[146] ^ x[48];
  assign t[107] = t[147] ^ x[49];
  assign t[108] = t[148] ^ x[50];
  assign t[109] = (x[2]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[2]);
  assign t[111] = (x[2]);
  assign t[112] = (x[2]);
  assign t[113] = (x[7]);
  assign t[114] = (x[7]);
  assign t[115] = (x[7]);
  assign t[116] = (x[7]);
  assign t[117] = (x[12]);
  assign t[118] = (x[12]);
  assign t[119] = (x[12]);
  assign t[11] = t[40] ^ t[15];
  assign t[120] = (x[12]);
  assign t[121] = (x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[17]);
  assign t[124] = (x[17]);
  assign t[125] = (x[22]);
  assign t[126] = (x[22]);
  assign t[127] = (x[22]);
  assign t[128] = (x[22]);
  assign t[129] = (x[27]);
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[130] = (x[27]);
  assign t[131] = (x[27]);
  assign t[132] = (x[27]);
  assign t[133] = (x[32]);
  assign t[134] = (x[32]);
  assign t[135] = (x[32]);
  assign t[136] = (x[32]);
  assign t[137] = (x[37]);
  assign t[138] = (x[37]);
  assign t[139] = (x[37]);
  assign t[13] = t[42] ^ t[43];
  assign t[140] = (x[37]);
  assign t[141] = (x[42]);
  assign t[142] = (x[42]);
  assign t[143] = (x[42]);
  assign t[144] = (x[42]);
  assign t[145] = (x[47]);
  assign t[146] = (x[47]);
  assign t[147] = (x[47]);
  assign t[148] = (x[47]);
  assign t[14] = t[15] & t[19];
  assign t[15] = ~(t[43]);
  assign t[16] = ~(t[40] ^ t[15]);
  assign t[17] = t[40] & t[20];
  assign t[18] = ~t[21];
  assign t[19] = t[40] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] ^ t[14];
  assign t[21] = ~(t[24] ^ t[25]);
  assign t[22] = t[43] ^ t[44];
  assign t[23] = t[40] ^ t[13];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[34] ^ t[27];
  assign t[29] = t[45] ^ t[32];
  assign t[2] = ~t[4];
  assign t[30] = t[46] ^ t[47];
  assign t[31] = t[32] & t[35];
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[45] ^ t[32]);
  assign t[34] = t[45] & t[36];
  assign t[35] = t[45] ^ t[37];
  assign t[36] = t[38] ^ t[31];
  assign t[37] = t[47] ^ t[48];
  assign t[38] = t[45] ^ t[30];
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[6];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[11];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[21];
  assign t[53] = t[63] ^ x[26];
  assign t[54] = t[64] ^ x[31];
  assign t[55] = t[65] ^ x[36];
  assign t[56] = t[66] ^ x[41];
  assign t[57] = t[67] ^ x[46];
  assign t[58] = t[68] ^ x[51];
  assign t[59] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[61] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[62] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[63] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[64] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[65] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[66] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[67] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[68] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[69] = t[109] ^ x[6];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[110] ^ x[3];
  assign t[71] = t[111] ^ x[4];
  assign t[72] = t[112] ^ x[5];
  assign t[73] = t[113] ^ x[11];
  assign t[74] = t[114] ^ x[8];
  assign t[75] = t[115] ^ x[9];
  assign t[76] = t[116] ^ x[10];
  assign t[77] = t[117] ^ x[16];
  assign t[78] = t[118] ^ x[13];
  assign t[79] = t[119] ^ x[14];
  assign t[7] = ~t[12];
  assign t[80] = t[120] ^ x[15];
  assign t[81] = t[121] ^ x[21];
  assign t[82] = t[122] ^ x[18];
  assign t[83] = t[123] ^ x[19];
  assign t[84] = t[124] ^ x[20];
  assign t[85] = t[125] ^ x[26];
  assign t[86] = t[126] ^ x[23];
  assign t[87] = t[127] ^ x[24];
  assign t[88] = t[128] ^ x[25];
  assign t[89] = t[129] ^ x[31];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[130] ^ x[28];
  assign t[91] = t[131] ^ x[29];
  assign t[92] = t[132] ^ x[30];
  assign t[93] = t[133] ^ x[36];
  assign t[94] = t[134] ^ x[33];
  assign t[95] = t[135] ^ x[34];
  assign t[96] = t[136] ^ x[35];
  assign t[97] = t[137] ^ x[41];
  assign t[98] = t[138] ^ x[38];
  assign t[99] = t[139] ^ x[39];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind133(x, y);
 input [51:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ^ x[40];
  assign t[101] = t[141] ^ x[46];
  assign t[102] = t[142] ^ x[43];
  assign t[103] = t[143] ^ x[44];
  assign t[104] = t[144] ^ x[45];
  assign t[105] = t[145] ^ x[51];
  assign t[106] = t[146] ^ x[48];
  assign t[107] = t[147] ^ x[49];
  assign t[108] = t[148] ^ x[50];
  assign t[109] = (x[2]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[2]);
  assign t[111] = (x[2]);
  assign t[112] = (x[2]);
  assign t[113] = (x[7]);
  assign t[114] = (x[7]);
  assign t[115] = (x[7]);
  assign t[116] = (x[7]);
  assign t[117] = (x[12]);
  assign t[118] = (x[12]);
  assign t[119] = (x[12]);
  assign t[11] = t[40] ^ t[15];
  assign t[120] = (x[12]);
  assign t[121] = (x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[17]);
  assign t[124] = (x[17]);
  assign t[125] = (x[22]);
  assign t[126] = (x[22]);
  assign t[127] = (x[22]);
  assign t[128] = (x[22]);
  assign t[129] = (x[27]);
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[130] = (x[27]);
  assign t[131] = (x[27]);
  assign t[132] = (x[27]);
  assign t[133] = (x[32]);
  assign t[134] = (x[32]);
  assign t[135] = (x[32]);
  assign t[136] = (x[32]);
  assign t[137] = (x[37]);
  assign t[138] = (x[37]);
  assign t[139] = (x[37]);
  assign t[13] = t[42] ^ t[43];
  assign t[140] = (x[37]);
  assign t[141] = (x[42]);
  assign t[142] = (x[42]);
  assign t[143] = (x[42]);
  assign t[144] = (x[42]);
  assign t[145] = (x[47]);
  assign t[146] = (x[47]);
  assign t[147] = (x[47]);
  assign t[148] = (x[47]);
  assign t[14] = t[15] & t[19];
  assign t[15] = ~(t[43]);
  assign t[16] = ~(t[40] ^ t[15]);
  assign t[17] = t[40] & t[20];
  assign t[18] = ~t[21];
  assign t[19] = t[40] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] ^ t[14];
  assign t[21] = ~(t[24] ^ t[25]);
  assign t[22] = t[43] ^ t[44];
  assign t[23] = t[40] ^ t[13];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[34] ^ t[27];
  assign t[29] = t[45] ^ t[32];
  assign t[2] = ~t[4];
  assign t[30] = t[46] ^ t[47];
  assign t[31] = t[32] & t[35];
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[45] ^ t[32]);
  assign t[34] = t[45] & t[36];
  assign t[35] = t[45] ^ t[37];
  assign t[36] = t[38] ^ t[31];
  assign t[37] = t[47] ^ t[48];
  assign t[38] = t[45] ^ t[30];
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[6];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[11];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[21];
  assign t[53] = t[63] ^ x[26];
  assign t[54] = t[64] ^ x[31];
  assign t[55] = t[65] ^ x[36];
  assign t[56] = t[66] ^ x[41];
  assign t[57] = t[67] ^ x[46];
  assign t[58] = t[68] ^ x[51];
  assign t[59] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[61] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[62] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[63] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[64] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[65] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[66] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[67] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[68] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[69] = t[109] ^ x[6];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[110] ^ x[3];
  assign t[71] = t[111] ^ x[4];
  assign t[72] = t[112] ^ x[5];
  assign t[73] = t[113] ^ x[11];
  assign t[74] = t[114] ^ x[8];
  assign t[75] = t[115] ^ x[9];
  assign t[76] = t[116] ^ x[10];
  assign t[77] = t[117] ^ x[16];
  assign t[78] = t[118] ^ x[13];
  assign t[79] = t[119] ^ x[14];
  assign t[7] = ~t[12];
  assign t[80] = t[120] ^ x[15];
  assign t[81] = t[121] ^ x[21];
  assign t[82] = t[122] ^ x[18];
  assign t[83] = t[123] ^ x[19];
  assign t[84] = t[124] ^ x[20];
  assign t[85] = t[125] ^ x[26];
  assign t[86] = t[126] ^ x[23];
  assign t[87] = t[127] ^ x[24];
  assign t[88] = t[128] ^ x[25];
  assign t[89] = t[129] ^ x[31];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[130] ^ x[28];
  assign t[91] = t[131] ^ x[29];
  assign t[92] = t[132] ^ x[30];
  assign t[93] = t[133] ^ x[36];
  assign t[94] = t[134] ^ x[33];
  assign t[95] = t[135] ^ x[34];
  assign t[96] = t[136] ^ x[35];
  assign t[97] = t[137] ^ x[41];
  assign t[98] = t[138] ^ x[38];
  assign t[99] = t[139] ^ x[39];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind134(x, y);
 input [51:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ^ x[40];
  assign t[101] = t[141] ^ x[46];
  assign t[102] = t[142] ^ x[43];
  assign t[103] = t[143] ^ x[44];
  assign t[104] = t[144] ^ x[45];
  assign t[105] = t[145] ^ x[51];
  assign t[106] = t[146] ^ x[48];
  assign t[107] = t[147] ^ x[49];
  assign t[108] = t[148] ^ x[50];
  assign t[109] = (x[2]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[2]);
  assign t[111] = (x[2]);
  assign t[112] = (x[2]);
  assign t[113] = (x[7]);
  assign t[114] = (x[7]);
  assign t[115] = (x[7]);
  assign t[116] = (x[7]);
  assign t[117] = (x[12]);
  assign t[118] = (x[12]);
  assign t[119] = (x[12]);
  assign t[11] = t[40] ^ t[15];
  assign t[120] = (x[12]);
  assign t[121] = (x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[17]);
  assign t[124] = (x[17]);
  assign t[125] = (x[22]);
  assign t[126] = (x[22]);
  assign t[127] = (x[22]);
  assign t[128] = (x[22]);
  assign t[129] = (x[27]);
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[130] = (x[27]);
  assign t[131] = (x[27]);
  assign t[132] = (x[27]);
  assign t[133] = (x[32]);
  assign t[134] = (x[32]);
  assign t[135] = (x[32]);
  assign t[136] = (x[32]);
  assign t[137] = (x[37]);
  assign t[138] = (x[37]);
  assign t[139] = (x[37]);
  assign t[13] = t[42] ^ t[43];
  assign t[140] = (x[37]);
  assign t[141] = (x[42]);
  assign t[142] = (x[42]);
  assign t[143] = (x[42]);
  assign t[144] = (x[42]);
  assign t[145] = (x[47]);
  assign t[146] = (x[47]);
  assign t[147] = (x[47]);
  assign t[148] = (x[47]);
  assign t[14] = t[15] & t[19];
  assign t[15] = ~(t[43]);
  assign t[16] = ~(t[40] ^ t[15]);
  assign t[17] = t[40] & t[20];
  assign t[18] = ~t[21];
  assign t[19] = t[40] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] ^ t[14];
  assign t[21] = ~(t[24] ^ t[25]);
  assign t[22] = t[43] ^ t[44];
  assign t[23] = t[40] ^ t[13];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[34] ^ t[27];
  assign t[29] = t[45] ^ t[32];
  assign t[2] = ~t[4];
  assign t[30] = t[46] ^ t[47];
  assign t[31] = t[32] & t[35];
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[45] ^ t[32]);
  assign t[34] = t[45] & t[36];
  assign t[35] = t[45] ^ t[37];
  assign t[36] = t[38] ^ t[31];
  assign t[37] = t[47] ^ t[48];
  assign t[38] = t[45] ^ t[30];
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[6];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[11];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[21];
  assign t[53] = t[63] ^ x[26];
  assign t[54] = t[64] ^ x[31];
  assign t[55] = t[65] ^ x[36];
  assign t[56] = t[66] ^ x[41];
  assign t[57] = t[67] ^ x[46];
  assign t[58] = t[68] ^ x[51];
  assign t[59] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[61] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[62] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[63] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[64] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[65] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[66] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[67] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[68] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[69] = t[109] ^ x[6];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[110] ^ x[3];
  assign t[71] = t[111] ^ x[4];
  assign t[72] = t[112] ^ x[5];
  assign t[73] = t[113] ^ x[11];
  assign t[74] = t[114] ^ x[8];
  assign t[75] = t[115] ^ x[9];
  assign t[76] = t[116] ^ x[10];
  assign t[77] = t[117] ^ x[16];
  assign t[78] = t[118] ^ x[13];
  assign t[79] = t[119] ^ x[14];
  assign t[7] = ~t[12];
  assign t[80] = t[120] ^ x[15];
  assign t[81] = t[121] ^ x[21];
  assign t[82] = t[122] ^ x[18];
  assign t[83] = t[123] ^ x[19];
  assign t[84] = t[124] ^ x[20];
  assign t[85] = t[125] ^ x[26];
  assign t[86] = t[126] ^ x[23];
  assign t[87] = t[127] ^ x[24];
  assign t[88] = t[128] ^ x[25];
  assign t[89] = t[129] ^ x[31];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[130] ^ x[28];
  assign t[91] = t[131] ^ x[29];
  assign t[92] = t[132] ^ x[30];
  assign t[93] = t[133] ^ x[36];
  assign t[94] = t[134] ^ x[33];
  assign t[95] = t[135] ^ x[34];
  assign t[96] = t[136] ^ x[35];
  assign t[97] = t[137] ^ x[41];
  assign t[98] = t[138] ^ x[38];
  assign t[99] = t[139] ^ x[39];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind135(x, y);
 input [51:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[140] ^ x[40];
  assign t[101] = t[141] ^ x[46];
  assign t[102] = t[142] ^ x[43];
  assign t[103] = t[143] ^ x[44];
  assign t[104] = t[144] ^ x[45];
  assign t[105] = t[145] ^ x[51];
  assign t[106] = t[146] ^ x[48];
  assign t[107] = t[147] ^ x[49];
  assign t[108] = t[148] ^ x[50];
  assign t[109] = (x[2]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[2]);
  assign t[111] = (x[2]);
  assign t[112] = (x[2]);
  assign t[113] = (x[7]);
  assign t[114] = (x[7]);
  assign t[115] = (x[7]);
  assign t[116] = (x[7]);
  assign t[117] = (x[12]);
  assign t[118] = (x[12]);
  assign t[119] = (x[12]);
  assign t[11] = t[40] ^ t[15];
  assign t[120] = (x[12]);
  assign t[121] = (x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[17]);
  assign t[124] = (x[17]);
  assign t[125] = (x[22]);
  assign t[126] = (x[22]);
  assign t[127] = (x[22]);
  assign t[128] = (x[22]);
  assign t[129] = (x[27]);
  assign t[12] = ~(t[18] ^ t[41]);
  assign t[130] = (x[27]);
  assign t[131] = (x[27]);
  assign t[132] = (x[27]);
  assign t[133] = (x[32]);
  assign t[134] = (x[32]);
  assign t[135] = (x[32]);
  assign t[136] = (x[32]);
  assign t[137] = (x[37]);
  assign t[138] = (x[37]);
  assign t[139] = (x[37]);
  assign t[13] = t[42] ^ t[43];
  assign t[140] = (x[37]);
  assign t[141] = (x[42]);
  assign t[142] = (x[42]);
  assign t[143] = (x[42]);
  assign t[144] = (x[42]);
  assign t[145] = (x[47]);
  assign t[146] = (x[47]);
  assign t[147] = (x[47]);
  assign t[148] = (x[47]);
  assign t[14] = t[15] & t[19];
  assign t[15] = ~(t[43]);
  assign t[16] = ~(t[40] ^ t[15]);
  assign t[17] = t[40] & t[20];
  assign t[18] = ~t[21];
  assign t[19] = t[40] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] ^ t[14];
  assign t[21] = ~(t[24] ^ t[25]);
  assign t[22] = t[43] ^ t[44];
  assign t[23] = t[40] ^ t[13];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[34] ^ t[27];
  assign t[29] = t[45] ^ t[32];
  assign t[2] = ~t[4];
  assign t[30] = t[46] ^ t[47];
  assign t[31] = t[32] & t[35];
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[45] ^ t[32]);
  assign t[34] = t[45] & t[36];
  assign t[35] = t[45] ^ t[37];
  assign t[36] = t[38] ^ t[31];
  assign t[37] = t[47] ^ t[48];
  assign t[38] = t[45] ^ t[30];
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = t[59] ^ x[6];
  assign t[4] = ~(t[7] ^ t[39]);
  assign t[50] = t[60] ^ x[11];
  assign t[51] = t[61] ^ x[16];
  assign t[52] = t[62] ^ x[21];
  assign t[53] = t[63] ^ x[26];
  assign t[54] = t[64] ^ x[31];
  assign t[55] = t[65] ^ x[36];
  assign t[56] = t[66] ^ x[41];
  assign t[57] = t[67] ^ x[46];
  assign t[58] = t[68] ^ x[51];
  assign t[59] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[61] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[62] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[63] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[64] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[65] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[66] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[67] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[68] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[69] = t[109] ^ x[6];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[110] ^ x[3];
  assign t[71] = t[111] ^ x[4];
  assign t[72] = t[112] ^ x[5];
  assign t[73] = t[113] ^ x[11];
  assign t[74] = t[114] ^ x[8];
  assign t[75] = t[115] ^ x[9];
  assign t[76] = t[116] ^ x[10];
  assign t[77] = t[117] ^ x[16];
  assign t[78] = t[118] ^ x[13];
  assign t[79] = t[119] ^ x[14];
  assign t[7] = ~t[12];
  assign t[80] = t[120] ^ x[15];
  assign t[81] = t[121] ^ x[21];
  assign t[82] = t[122] ^ x[18];
  assign t[83] = t[123] ^ x[19];
  assign t[84] = t[124] ^ x[20];
  assign t[85] = t[125] ^ x[26];
  assign t[86] = t[126] ^ x[23];
  assign t[87] = t[127] ^ x[24];
  assign t[88] = t[128] ^ x[25];
  assign t[89] = t[129] ^ x[31];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[130] ^ x[28];
  assign t[91] = t[131] ^ x[29];
  assign t[92] = t[132] ^ x[30];
  assign t[93] = t[133] ^ x[36];
  assign t[94] = t[134] ^ x[33];
  assign t[95] = t[135] ^ x[34];
  assign t[96] = t[136] ^ x[35];
  assign t[97] = t[137] ^ x[41];
  assign t[98] = t[138] ^ x[38];
  assign t[99] = t[139] ^ x[39];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind136(x, y);
 input [36:0] x;
 output y;

 wire [95:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[22] ^ t[10]);
  assign t[12] = ~t[13];
  assign t[13] = ~(t[14]);
  assign t[14] = t[15] ^ t[16];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[17] & t[18];
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[25] ^ t[17]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = (t[31]);
  assign t[25] = (t[32]);
  assign t[26] = t[33] ^ x[6];
  assign t[27] = t[34] ^ x[11];
  assign t[28] = t[35] ^ x[16];
  assign t[29] = t[36] ^ x[21];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[26];
  assign t[31] = t[38] ^ x[31];
  assign t[32] = t[39] ^ x[36];
  assign t[33] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[34] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[35] = (~t[48] & t[49] & t[50] & t[51]) | (t[48] & ~t[50] & ~t[51]) | (t[48] & ~t[49] & ~t[51]) | (t[48] & ~t[49] & ~t[50]);
  assign t[36] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[37] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[38] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[39] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[6];
  assign t[41] = t[69] ^ x[3];
  assign t[42] = t[70] ^ x[4];
  assign t[43] = t[71] ^ x[5];
  assign t[44] = t[72] ^ x[11];
  assign t[45] = t[73] ^ x[8];
  assign t[46] = t[74] ^ x[9];
  assign t[47] = t[75] ^ x[10];
  assign t[48] = t[76] ^ x[16];
  assign t[49] = t[77] ^ x[13];
  assign t[4] = ~(t[6] ^ t[19]);
  assign t[50] = t[78] ^ x[14];
  assign t[51] = t[79] ^ x[15];
  assign t[52] = t[80] ^ x[21];
  assign t[53] = t[81] ^ x[18];
  assign t[54] = t[82] ^ x[19];
  assign t[55] = t[83] ^ x[20];
  assign t[56] = t[84] ^ x[26];
  assign t[57] = t[85] ^ x[23];
  assign t[58] = t[86] ^ x[24];
  assign t[59] = t[87] ^ x[25];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[31];
  assign t[61] = t[89] ^ x[28];
  assign t[62] = t[90] ^ x[29];
  assign t[63] = t[91] ^ x[30];
  assign t[64] = t[92] ^ x[36];
  assign t[65] = t[93] ^ x[33];
  assign t[66] = t[94] ^ x[34];
  assign t[67] = t[95] ^ x[35];
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[2]);
  assign t[71] = (x[2]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[7]);
  assign t[75] = (x[7]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[12]);
  assign t[79] = (x[12]);
  assign t[7] = t[20] ^ t[21];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[17]);
  assign t[83] = (x[17]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[22]);
  assign t[87] = (x[22]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[27]);
  assign t[91] = (x[27]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[94] = (x[32]);
  assign t[95] = (x[32]);
  assign t[9] = ~t[12];
  assign y = (t[0]);
endmodule

module R2ind137(x, y);
 input [36:0] x;
 output y;

 wire [95:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[22] ^ t[10]);
  assign t[12] = ~t[13];
  assign t[13] = ~(t[14]);
  assign t[14] = t[15] ^ t[16];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[17] & t[18];
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[25] ^ t[17]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = (t[31]);
  assign t[25] = (t[32]);
  assign t[26] = t[33] ^ x[6];
  assign t[27] = t[34] ^ x[11];
  assign t[28] = t[35] ^ x[16];
  assign t[29] = t[36] ^ x[21];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[26];
  assign t[31] = t[38] ^ x[31];
  assign t[32] = t[39] ^ x[36];
  assign t[33] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[34] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[35] = (~t[48] & t[49] & t[50] & t[51]) | (t[48] & ~t[50] & ~t[51]) | (t[48] & ~t[49] & ~t[51]) | (t[48] & ~t[49] & ~t[50]);
  assign t[36] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[37] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[38] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[39] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[6];
  assign t[41] = t[69] ^ x[3];
  assign t[42] = t[70] ^ x[4];
  assign t[43] = t[71] ^ x[5];
  assign t[44] = t[72] ^ x[11];
  assign t[45] = t[73] ^ x[8];
  assign t[46] = t[74] ^ x[9];
  assign t[47] = t[75] ^ x[10];
  assign t[48] = t[76] ^ x[16];
  assign t[49] = t[77] ^ x[13];
  assign t[4] = ~(t[6] ^ t[19]);
  assign t[50] = t[78] ^ x[14];
  assign t[51] = t[79] ^ x[15];
  assign t[52] = t[80] ^ x[21];
  assign t[53] = t[81] ^ x[18];
  assign t[54] = t[82] ^ x[19];
  assign t[55] = t[83] ^ x[20];
  assign t[56] = t[84] ^ x[26];
  assign t[57] = t[85] ^ x[23];
  assign t[58] = t[86] ^ x[24];
  assign t[59] = t[87] ^ x[25];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[31];
  assign t[61] = t[89] ^ x[28];
  assign t[62] = t[90] ^ x[29];
  assign t[63] = t[91] ^ x[30];
  assign t[64] = t[92] ^ x[36];
  assign t[65] = t[93] ^ x[33];
  assign t[66] = t[94] ^ x[34];
  assign t[67] = t[95] ^ x[35];
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[2]);
  assign t[71] = (x[2]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[7]);
  assign t[75] = (x[7]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[12]);
  assign t[79] = (x[12]);
  assign t[7] = t[20] ^ t[21];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[17]);
  assign t[83] = (x[17]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[22]);
  assign t[87] = (x[22]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[27]);
  assign t[91] = (x[27]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[94] = (x[32]);
  assign t[95] = (x[32]);
  assign t[9] = ~t[12];
  assign y = (t[0]);
endmodule

module R2ind138(x, y);
 input [36:0] x;
 output y;

 wire [95:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[22] ^ t[10]);
  assign t[12] = ~t[13];
  assign t[13] = ~(t[14]);
  assign t[14] = t[15] ^ t[16];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[17] & t[18];
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[25] ^ t[17]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = (t[31]);
  assign t[25] = (t[32]);
  assign t[26] = t[33] ^ x[6];
  assign t[27] = t[34] ^ x[11];
  assign t[28] = t[35] ^ x[16];
  assign t[29] = t[36] ^ x[21];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[26];
  assign t[31] = t[38] ^ x[31];
  assign t[32] = t[39] ^ x[36];
  assign t[33] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[34] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[35] = (~t[48] & t[49] & t[50] & t[51]) | (t[48] & ~t[50] & ~t[51]) | (t[48] & ~t[49] & ~t[51]) | (t[48] & ~t[49] & ~t[50]);
  assign t[36] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[37] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[38] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[39] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[6];
  assign t[41] = t[69] ^ x[3];
  assign t[42] = t[70] ^ x[4];
  assign t[43] = t[71] ^ x[5];
  assign t[44] = t[72] ^ x[11];
  assign t[45] = t[73] ^ x[8];
  assign t[46] = t[74] ^ x[9];
  assign t[47] = t[75] ^ x[10];
  assign t[48] = t[76] ^ x[16];
  assign t[49] = t[77] ^ x[13];
  assign t[4] = ~(t[6] ^ t[19]);
  assign t[50] = t[78] ^ x[14];
  assign t[51] = t[79] ^ x[15];
  assign t[52] = t[80] ^ x[21];
  assign t[53] = t[81] ^ x[18];
  assign t[54] = t[82] ^ x[19];
  assign t[55] = t[83] ^ x[20];
  assign t[56] = t[84] ^ x[26];
  assign t[57] = t[85] ^ x[23];
  assign t[58] = t[86] ^ x[24];
  assign t[59] = t[87] ^ x[25];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[31];
  assign t[61] = t[89] ^ x[28];
  assign t[62] = t[90] ^ x[29];
  assign t[63] = t[91] ^ x[30];
  assign t[64] = t[92] ^ x[36];
  assign t[65] = t[93] ^ x[33];
  assign t[66] = t[94] ^ x[34];
  assign t[67] = t[95] ^ x[35];
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[2]);
  assign t[71] = (x[2]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[7]);
  assign t[75] = (x[7]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[12]);
  assign t[79] = (x[12]);
  assign t[7] = t[20] ^ t[21];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[17]);
  assign t[83] = (x[17]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[22]);
  assign t[87] = (x[22]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[27]);
  assign t[91] = (x[27]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[94] = (x[32]);
  assign t[95] = (x[32]);
  assign t[9] = ~t[12];
  assign y = (t[0]);
endmodule

module R2ind139(x, y);
 input [36:0] x;
 output y;

 wire [95:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[22] ^ t[10]);
  assign t[12] = ~t[13];
  assign t[13] = ~(t[14]);
  assign t[14] = t[15] ^ t[16];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[17] & t[18];
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[25] ^ t[17]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = (t[31]);
  assign t[25] = (t[32]);
  assign t[26] = t[33] ^ x[6];
  assign t[27] = t[34] ^ x[11];
  assign t[28] = t[35] ^ x[16];
  assign t[29] = t[36] ^ x[21];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[26];
  assign t[31] = t[38] ^ x[31];
  assign t[32] = t[39] ^ x[36];
  assign t[33] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[34] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[35] = (~t[48] & t[49] & t[50] & t[51]) | (t[48] & ~t[50] & ~t[51]) | (t[48] & ~t[49] & ~t[51]) | (t[48] & ~t[49] & ~t[50]);
  assign t[36] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[37] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[38] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[39] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[6];
  assign t[41] = t[69] ^ x[3];
  assign t[42] = t[70] ^ x[4];
  assign t[43] = t[71] ^ x[5];
  assign t[44] = t[72] ^ x[11];
  assign t[45] = t[73] ^ x[8];
  assign t[46] = t[74] ^ x[9];
  assign t[47] = t[75] ^ x[10];
  assign t[48] = t[76] ^ x[16];
  assign t[49] = t[77] ^ x[13];
  assign t[4] = ~(t[6] ^ t[19]);
  assign t[50] = t[78] ^ x[14];
  assign t[51] = t[79] ^ x[15];
  assign t[52] = t[80] ^ x[21];
  assign t[53] = t[81] ^ x[18];
  assign t[54] = t[82] ^ x[19];
  assign t[55] = t[83] ^ x[20];
  assign t[56] = t[84] ^ x[26];
  assign t[57] = t[85] ^ x[23];
  assign t[58] = t[86] ^ x[24];
  assign t[59] = t[87] ^ x[25];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[31];
  assign t[61] = t[89] ^ x[28];
  assign t[62] = t[90] ^ x[29];
  assign t[63] = t[91] ^ x[30];
  assign t[64] = t[92] ^ x[36];
  assign t[65] = t[93] ^ x[33];
  assign t[66] = t[94] ^ x[34];
  assign t[67] = t[95] ^ x[35];
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[2]);
  assign t[71] = (x[2]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[7]);
  assign t[75] = (x[7]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[12]);
  assign t[79] = (x[12]);
  assign t[7] = t[20] ^ t[21];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[17]);
  assign t[83] = (x[17]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[22]);
  assign t[87] = (x[22]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[27]);
  assign t[91] = (x[27]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[94] = (x[32]);
  assign t[95] = (x[32]);
  assign t[9] = ~t[12];
  assign y = (t[0]);
endmodule

module R2ind140(x, y);
 input [46:0] x;
 output y;

 wire [125:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[12]);
  assign t[101] = (x[12]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[17]);
  assign t[105] = (x[17]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[22]);
  assign t[10] = t[28] ^ t[29];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[27]);
  assign t[113] = (x[27]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[32]);
  assign t[117] = (x[32]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[37]);
  assign t[121] = (x[37]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[124] = (x[42]);
  assign t[125] = (x[42]);
  assign t[12] = ~(t[29]);
  assign t[13] = ~(t[30] ^ t[12]);
  assign t[14] = ~t[16];
  assign t[15] = t[30] ^ t[17];
  assign t[16] = ~(t[18]);
  assign t[17] = t[29] ^ t[31];
  assign t[18] = t[19] ^ t[20];
  assign t[19] = t[21] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] & t[24];
  assign t[21] = t[32] ^ t[33];
  assign t[22] = t[23] & t[25];
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[34] ^ t[23]);
  assign t[25] = t[34] ^ t[26];
  assign t[26] = t[33] ^ t[35];
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = (t[43]);
  assign t[35] = (t[44]);
  assign t[36] = t[45] ^ x[6];
  assign t[37] = t[46] ^ x[11];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[26];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = t[51] ^ x[36];
  assign t[43] = t[52] ^ x[41];
  assign t[44] = t[53] ^ x[46];
  assign t[45] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[46] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[47] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[48] = (~t[66] & t[67] & t[68] & t[69]) | (t[66] & ~t[68] & ~t[69]) | (t[66] & ~t[67] & ~t[69]) | (t[66] & ~t[67] & ~t[68]);
  assign t[49] = (~t[70] & t[71] & t[72] & t[73]) | (t[70] & ~t[72] & ~t[73]) | (t[70] & ~t[71] & ~t[73]) | (t[70] & ~t[71] & ~t[72]);
  assign t[4] = ~(t[6] ^ t[27]);
  assign t[50] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[51] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[52] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[53] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[54] = t[90] ^ x[6];
  assign t[55] = t[91] ^ x[3];
  assign t[56] = t[92] ^ x[4];
  assign t[57] = t[93] ^ x[5];
  assign t[58] = t[94] ^ x[11];
  assign t[59] = t[95] ^ x[8];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[9];
  assign t[61] = t[97] ^ x[10];
  assign t[62] = t[98] ^ x[16];
  assign t[63] = t[99] ^ x[13];
  assign t[64] = t[100] ^ x[14];
  assign t[65] = t[101] ^ x[15];
  assign t[66] = t[102] ^ x[21];
  assign t[67] = t[103] ^ x[18];
  assign t[68] = t[104] ^ x[19];
  assign t[69] = t[105] ^ x[20];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[26];
  assign t[71] = t[107] ^ x[23];
  assign t[72] = t[108] ^ x[24];
  assign t[73] = t[109] ^ x[25];
  assign t[74] = t[110] ^ x[31];
  assign t[75] = t[111] ^ x[28];
  assign t[76] = t[112] ^ x[29];
  assign t[77] = t[113] ^ x[30];
  assign t[78] = t[114] ^ x[36];
  assign t[79] = t[115] ^ x[33];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[34];
  assign t[81] = t[117] ^ x[35];
  assign t[82] = t[118] ^ x[41];
  assign t[83] = t[119] ^ x[38];
  assign t[84] = t[120] ^ x[39];
  assign t[85] = t[121] ^ x[40];
  assign t[86] = t[122] ^ x[46];
  assign t[87] = t[123] ^ x[43];
  assign t[88] = t[124] ^ x[44];
  assign t[89] = t[125] ^ x[45];
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[2]);
  assign t[93] = (x[2]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[7]);
  assign t[97] = (x[7]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~t[14];
  assign y = (t[0]);
endmodule

module R2ind141(x, y);
 input [46:0] x;
 output y;

 wire [125:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[12]);
  assign t[101] = (x[12]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[17]);
  assign t[105] = (x[17]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[22]);
  assign t[10] = t[28] ^ t[29];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[27]);
  assign t[113] = (x[27]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[32]);
  assign t[117] = (x[32]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[37]);
  assign t[121] = (x[37]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[124] = (x[42]);
  assign t[125] = (x[42]);
  assign t[12] = ~(t[29]);
  assign t[13] = ~(t[30] ^ t[12]);
  assign t[14] = ~t[16];
  assign t[15] = t[30] ^ t[17];
  assign t[16] = ~(t[18]);
  assign t[17] = t[29] ^ t[31];
  assign t[18] = t[19] ^ t[20];
  assign t[19] = t[21] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] & t[24];
  assign t[21] = t[32] ^ t[33];
  assign t[22] = t[23] & t[25];
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[34] ^ t[23]);
  assign t[25] = t[34] ^ t[26];
  assign t[26] = t[33] ^ t[35];
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = (t[43]);
  assign t[35] = (t[44]);
  assign t[36] = t[45] ^ x[6];
  assign t[37] = t[46] ^ x[11];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[26];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = t[51] ^ x[36];
  assign t[43] = t[52] ^ x[41];
  assign t[44] = t[53] ^ x[46];
  assign t[45] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[46] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[47] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[48] = (~t[66] & t[67] & t[68] & t[69]) | (t[66] & ~t[68] & ~t[69]) | (t[66] & ~t[67] & ~t[69]) | (t[66] & ~t[67] & ~t[68]);
  assign t[49] = (~t[70] & t[71] & t[72] & t[73]) | (t[70] & ~t[72] & ~t[73]) | (t[70] & ~t[71] & ~t[73]) | (t[70] & ~t[71] & ~t[72]);
  assign t[4] = ~(t[6] ^ t[27]);
  assign t[50] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[51] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[52] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[53] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[54] = t[90] ^ x[6];
  assign t[55] = t[91] ^ x[3];
  assign t[56] = t[92] ^ x[4];
  assign t[57] = t[93] ^ x[5];
  assign t[58] = t[94] ^ x[11];
  assign t[59] = t[95] ^ x[8];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[9];
  assign t[61] = t[97] ^ x[10];
  assign t[62] = t[98] ^ x[16];
  assign t[63] = t[99] ^ x[13];
  assign t[64] = t[100] ^ x[14];
  assign t[65] = t[101] ^ x[15];
  assign t[66] = t[102] ^ x[21];
  assign t[67] = t[103] ^ x[18];
  assign t[68] = t[104] ^ x[19];
  assign t[69] = t[105] ^ x[20];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[26];
  assign t[71] = t[107] ^ x[23];
  assign t[72] = t[108] ^ x[24];
  assign t[73] = t[109] ^ x[25];
  assign t[74] = t[110] ^ x[31];
  assign t[75] = t[111] ^ x[28];
  assign t[76] = t[112] ^ x[29];
  assign t[77] = t[113] ^ x[30];
  assign t[78] = t[114] ^ x[36];
  assign t[79] = t[115] ^ x[33];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[34];
  assign t[81] = t[117] ^ x[35];
  assign t[82] = t[118] ^ x[41];
  assign t[83] = t[119] ^ x[38];
  assign t[84] = t[120] ^ x[39];
  assign t[85] = t[121] ^ x[40];
  assign t[86] = t[122] ^ x[46];
  assign t[87] = t[123] ^ x[43];
  assign t[88] = t[124] ^ x[44];
  assign t[89] = t[125] ^ x[45];
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[2]);
  assign t[93] = (x[2]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[7]);
  assign t[97] = (x[7]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~t[14];
  assign y = (t[0]);
endmodule

module R2ind142(x, y);
 input [46:0] x;
 output y;

 wire [125:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[12]);
  assign t[101] = (x[12]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[17]);
  assign t[105] = (x[17]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[22]);
  assign t[10] = t[28] ^ t[29];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[27]);
  assign t[113] = (x[27]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[32]);
  assign t[117] = (x[32]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[37]);
  assign t[121] = (x[37]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[124] = (x[42]);
  assign t[125] = (x[42]);
  assign t[12] = ~(t[29]);
  assign t[13] = ~(t[30] ^ t[12]);
  assign t[14] = ~t[16];
  assign t[15] = t[30] ^ t[17];
  assign t[16] = ~(t[18]);
  assign t[17] = t[29] ^ t[31];
  assign t[18] = t[19] ^ t[20];
  assign t[19] = t[21] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] & t[24];
  assign t[21] = t[32] ^ t[33];
  assign t[22] = t[23] & t[25];
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[34] ^ t[23]);
  assign t[25] = t[34] ^ t[26];
  assign t[26] = t[33] ^ t[35];
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = (t[43]);
  assign t[35] = (t[44]);
  assign t[36] = t[45] ^ x[6];
  assign t[37] = t[46] ^ x[11];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[26];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = t[51] ^ x[36];
  assign t[43] = t[52] ^ x[41];
  assign t[44] = t[53] ^ x[46];
  assign t[45] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[46] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[47] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[48] = (~t[66] & t[67] & t[68] & t[69]) | (t[66] & ~t[68] & ~t[69]) | (t[66] & ~t[67] & ~t[69]) | (t[66] & ~t[67] & ~t[68]);
  assign t[49] = (~t[70] & t[71] & t[72] & t[73]) | (t[70] & ~t[72] & ~t[73]) | (t[70] & ~t[71] & ~t[73]) | (t[70] & ~t[71] & ~t[72]);
  assign t[4] = ~(t[6] ^ t[27]);
  assign t[50] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[51] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[52] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[53] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[54] = t[90] ^ x[6];
  assign t[55] = t[91] ^ x[3];
  assign t[56] = t[92] ^ x[4];
  assign t[57] = t[93] ^ x[5];
  assign t[58] = t[94] ^ x[11];
  assign t[59] = t[95] ^ x[8];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[9];
  assign t[61] = t[97] ^ x[10];
  assign t[62] = t[98] ^ x[16];
  assign t[63] = t[99] ^ x[13];
  assign t[64] = t[100] ^ x[14];
  assign t[65] = t[101] ^ x[15];
  assign t[66] = t[102] ^ x[21];
  assign t[67] = t[103] ^ x[18];
  assign t[68] = t[104] ^ x[19];
  assign t[69] = t[105] ^ x[20];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[26];
  assign t[71] = t[107] ^ x[23];
  assign t[72] = t[108] ^ x[24];
  assign t[73] = t[109] ^ x[25];
  assign t[74] = t[110] ^ x[31];
  assign t[75] = t[111] ^ x[28];
  assign t[76] = t[112] ^ x[29];
  assign t[77] = t[113] ^ x[30];
  assign t[78] = t[114] ^ x[36];
  assign t[79] = t[115] ^ x[33];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[34];
  assign t[81] = t[117] ^ x[35];
  assign t[82] = t[118] ^ x[41];
  assign t[83] = t[119] ^ x[38];
  assign t[84] = t[120] ^ x[39];
  assign t[85] = t[121] ^ x[40];
  assign t[86] = t[122] ^ x[46];
  assign t[87] = t[123] ^ x[43];
  assign t[88] = t[124] ^ x[44];
  assign t[89] = t[125] ^ x[45];
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[2]);
  assign t[93] = (x[2]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[7]);
  assign t[97] = (x[7]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~t[14];
  assign y = (t[0]);
endmodule

module R2ind143(x, y);
 input [46:0] x;
 output y;

 wire [125:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[12]);
  assign t[101] = (x[12]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[17]);
  assign t[105] = (x[17]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[22]);
  assign t[10] = t[28] ^ t[29];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[27]);
  assign t[113] = (x[27]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[32]);
  assign t[117] = (x[32]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[37]);
  assign t[121] = (x[37]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[124] = (x[42]);
  assign t[125] = (x[42]);
  assign t[12] = ~(t[29]);
  assign t[13] = ~(t[30] ^ t[12]);
  assign t[14] = ~t[16];
  assign t[15] = t[30] ^ t[17];
  assign t[16] = ~(t[18]);
  assign t[17] = t[29] ^ t[31];
  assign t[18] = t[19] ^ t[20];
  assign t[19] = t[21] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] & t[24];
  assign t[21] = t[32] ^ t[33];
  assign t[22] = t[23] & t[25];
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[34] ^ t[23]);
  assign t[25] = t[34] ^ t[26];
  assign t[26] = t[33] ^ t[35];
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = (t[43]);
  assign t[35] = (t[44]);
  assign t[36] = t[45] ^ x[6];
  assign t[37] = t[46] ^ x[11];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[26];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = t[51] ^ x[36];
  assign t[43] = t[52] ^ x[41];
  assign t[44] = t[53] ^ x[46];
  assign t[45] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[46] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[47] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[48] = (~t[66] & t[67] & t[68] & t[69]) | (t[66] & ~t[68] & ~t[69]) | (t[66] & ~t[67] & ~t[69]) | (t[66] & ~t[67] & ~t[68]);
  assign t[49] = (~t[70] & t[71] & t[72] & t[73]) | (t[70] & ~t[72] & ~t[73]) | (t[70] & ~t[71] & ~t[73]) | (t[70] & ~t[71] & ~t[72]);
  assign t[4] = ~(t[6] ^ t[27]);
  assign t[50] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[51] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[52] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[53] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[54] = t[90] ^ x[6];
  assign t[55] = t[91] ^ x[3];
  assign t[56] = t[92] ^ x[4];
  assign t[57] = t[93] ^ x[5];
  assign t[58] = t[94] ^ x[11];
  assign t[59] = t[95] ^ x[8];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[9];
  assign t[61] = t[97] ^ x[10];
  assign t[62] = t[98] ^ x[16];
  assign t[63] = t[99] ^ x[13];
  assign t[64] = t[100] ^ x[14];
  assign t[65] = t[101] ^ x[15];
  assign t[66] = t[102] ^ x[21];
  assign t[67] = t[103] ^ x[18];
  assign t[68] = t[104] ^ x[19];
  assign t[69] = t[105] ^ x[20];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[26];
  assign t[71] = t[107] ^ x[23];
  assign t[72] = t[108] ^ x[24];
  assign t[73] = t[109] ^ x[25];
  assign t[74] = t[110] ^ x[31];
  assign t[75] = t[111] ^ x[28];
  assign t[76] = t[112] ^ x[29];
  assign t[77] = t[113] ^ x[30];
  assign t[78] = t[114] ^ x[36];
  assign t[79] = t[115] ^ x[33];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[34];
  assign t[81] = t[117] ^ x[35];
  assign t[82] = t[118] ^ x[41];
  assign t[83] = t[119] ^ x[38];
  assign t[84] = t[120] ^ x[39];
  assign t[85] = t[121] ^ x[40];
  assign t[86] = t[122] ^ x[46];
  assign t[87] = t[123] ^ x[43];
  assign t[88] = t[124] ^ x[44];
  assign t[89] = t[125] ^ x[45];
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[2]);
  assign t[93] = (x[2]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[7]);
  assign t[97] = (x[7]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~t[14];
  assign y = (t[0]);
endmodule

module R2ind144(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind145(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind146(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind147(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[38] ^ t[14]);
  assign t[16] = t[40] ^ t[39];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[38] ^ t[27];
  assign t[23] = t[41] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[39] ^ t[42];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[43]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[41] ^ t[29]);
  assign t[31] = t[44] ^ t[43];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[41] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[41] ^ t[36];
  assign t[36] = t[43] ^ t[45];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[38] & t[13];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind148(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[38] ^ t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind149(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[38] ^ t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind150(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[38] ^ t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind151(x, y);
 input [46:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2]);
  assign t[101] = (x[2]);
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[12]);
  assign t[109] = (x[12]);
  assign t[10] = t[17] ^ t[9];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[17]);
  assign t[113] = (x[17]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[22]);
  assign t[117] = (x[22]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[38] ^ t[15];
  assign t[120] = (x[27]);
  assign t[121] = (x[27]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[32]);
  assign t[125] = (x[32]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[37]);
  assign t[129] = (x[37]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[42]);
  assign t[133] = (x[42]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[13] = t[39] ^ t[40];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[40]);
  assign t[16] = ~(t[38] ^ t[15]);
  assign t[17] = t[38] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[41] ^ t[30];
  assign t[26] = t[40] ^ t[42];
  assign t[27] = t[38] ^ t[13];
  assign t[28] = t[43] ^ t[44];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[41] ^ t[30]);
  assign t[32] = t[41] & t[34];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[44] ^ t[45];
  assign t[36] = t[41] ^ t[28];
  assign t[37] = (t[46]);
  assign t[38] = (t[47]);
  assign t[39] = (t[48]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49]);
  assign t[41] = (t[50]);
  assign t[42] = (t[51]);
  assign t[43] = (t[52]);
  assign t[44] = (t[53]);
  assign t[45] = (t[54]);
  assign t[46] = t[55] ^ x[6];
  assign t[47] = t[56] ^ x[11];
  assign t[48] = t[57] ^ x[16];
  assign t[49] = t[58] ^ x[21];
  assign t[4] = ~(t[7] ^ t[37]);
  assign t[50] = t[59] ^ x[26];
  assign t[51] = t[60] ^ x[31];
  assign t[52] = t[61] ^ x[36];
  assign t[53] = t[62] ^ x[41];
  assign t[54] = t[63] ^ x[46];
  assign t[55] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[56] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[57] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[58] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[59] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[61] = (~t[88] & t[89] & t[90] & t[91]) | (t[88] & ~t[90] & ~t[91]) | (t[88] & ~t[89] & ~t[91]) | (t[88] & ~t[89] & ~t[90]);
  assign t[62] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[63] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[64] = t[100] ^ x[6];
  assign t[65] = t[101] ^ x[3];
  assign t[66] = t[102] ^ x[4];
  assign t[67] = t[103] ^ x[5];
  assign t[68] = t[104] ^ x[11];
  assign t[69] = t[105] ^ x[8];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[106] ^ x[9];
  assign t[71] = t[107] ^ x[10];
  assign t[72] = t[108] ^ x[16];
  assign t[73] = t[109] ^ x[13];
  assign t[74] = t[110] ^ x[14];
  assign t[75] = t[111] ^ x[15];
  assign t[76] = t[112] ^ x[21];
  assign t[77] = t[113] ^ x[18];
  assign t[78] = t[114] ^ x[19];
  assign t[79] = t[115] ^ x[20];
  assign t[7] = ~t[12];
  assign t[80] = t[116] ^ x[26];
  assign t[81] = t[117] ^ x[23];
  assign t[82] = t[118] ^ x[24];
  assign t[83] = t[119] ^ x[25];
  assign t[84] = t[120] ^ x[31];
  assign t[85] = t[121] ^ x[28];
  assign t[86] = t[122] ^ x[29];
  assign t[87] = t[123] ^ x[30];
  assign t[88] = t[124] ^ x[36];
  assign t[89] = t[125] ^ x[33];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[126] ^ x[34];
  assign t[91] = t[127] ^ x[35];
  assign t[92] = t[128] ^ x[41];
  assign t[93] = t[129] ^ x[38];
  assign t[94] = t[130] ^ x[39];
  assign t[95] = t[131] ^ x[40];
  assign t[96] = t[132] ^ x[46];
  assign t[97] = t[133] ^ x[43];
  assign t[98] = t[134] ^ x[44];
  assign t[99] = t[135] ^ x[45];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind152(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind153(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind154(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind155(x, y);
 input [36:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[18]);
  assign t[11] = ~(t[20] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[21] ^ t[22];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[21]);
  assign t[16] = ~(t[23] ^ t[15]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = t[31] ^ x[6];
  assign t[25] = t[32] ^ x[11];
  assign t[26] = t[33] ^ x[16];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = t[35] ^ x[26];
  assign t[29] = t[36] ^ x[31];
  assign t[2] = ~t[4];
  assign t[30] = t[37] ^ x[36];
  assign t[31] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[32] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[33] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[34] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[35] = (~t[54] & t[55] & t[56] & t[57]) | (t[54] & ~t[56] & ~t[57]) | (t[54] & ~t[55] & ~t[57]) | (t[54] & ~t[55] & ~t[56]);
  assign t[36] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[37] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[38] = t[66] ^ x[6];
  assign t[39] = t[67] ^ x[3];
  assign t[3] = ~(t[5]);
  assign t[40] = t[68] ^ x[4];
  assign t[41] = t[69] ^ x[5];
  assign t[42] = t[70] ^ x[11];
  assign t[43] = t[71] ^ x[8];
  assign t[44] = t[72] ^ x[9];
  assign t[45] = t[73] ^ x[10];
  assign t[46] = t[74] ^ x[16];
  assign t[47] = t[75] ^ x[13];
  assign t[48] = t[76] ^ x[14];
  assign t[49] = t[77] ^ x[15];
  assign t[4] = ~(t[6] ^ t[17]);
  assign t[50] = t[78] ^ x[21];
  assign t[51] = t[79] ^ x[18];
  assign t[52] = t[80] ^ x[19];
  assign t[53] = t[81] ^ x[20];
  assign t[54] = t[82] ^ x[26];
  assign t[55] = t[83] ^ x[23];
  assign t[56] = t[84] ^ x[24];
  assign t[57] = t[85] ^ x[25];
  assign t[58] = t[86] ^ x[31];
  assign t[59] = t[87] ^ x[28];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[88] ^ x[29];
  assign t[61] = t[89] ^ x[30];
  assign t[62] = t[90] ^ x[36];
  assign t[63] = t[91] ^ x[33];
  assign t[64] = t[92] ^ x[34];
  assign t[65] = t[93] ^ x[35];
  assign t[66] = (x[2]);
  assign t[67] = (x[2]);
  assign t[68] = (x[2]);
  assign t[69] = (x[2]);
  assign t[6] = ~t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[7]);
  assign t[72] = (x[7]);
  assign t[73] = (x[7]);
  assign t[74] = (x[12]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[12]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = t[18] ^ t[19];
  assign t[80] = (x[17]);
  assign t[81] = (x[17]);
  assign t[82] = (x[22]);
  assign t[83] = (x[22]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[27]);
  assign t[87] = (x[27]);
  assign t[88] = (x[27]);
  assign t[89] = (x[27]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (x[32]);
  assign t[91] = (x[32]);
  assign t[92] = (x[32]);
  assign t[93] = (x[32]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind156(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind157(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind158(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind159(x, y);
 input [46:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[17]);
  assign t[101] = (x[17]);
  assign t[102] = (x[17]);
  assign t[103] = (x[17]);
  assign t[104] = (x[22]);
  assign t[105] = (x[22]);
  assign t[106] = (x[22]);
  assign t[107] = (x[22]);
  assign t[108] = (x[27]);
  assign t[109] = (x[27]);
  assign t[10] = t[26] ^ t[27];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[32]);
  assign t[113] = (x[32]);
  assign t[114] = (x[32]);
  assign t[115] = (x[32]);
  assign t[116] = (x[37]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[37]);
  assign t[11] = t[12] & t[15];
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[28] ^ t[12]);
  assign t[14] = t[16] ^ t[17];
  assign t[15] = t[28] ^ t[18];
  assign t[16] = t[19] ^ t[20];
  assign t[17] = t[21] & t[22];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = t[30] ^ t[31];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] & t[23];
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = t[32] ^ t[24];
  assign t[24] = t[31] ^ t[33];
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[6];
  assign t[35] = t[44] ^ x[11];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[26];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5]);
  assign t[40] = t[49] ^ x[36];
  assign t[41] = t[50] ^ x[41];
  assign t[42] = t[51] ^ x[46];
  assign t[43] = (~t[52] & t[53] & t[54] & t[55]) | (t[52] & ~t[54] & ~t[55]) | (t[52] & ~t[53] & ~t[55]) | (t[52] & ~t[53] & ~t[54]);
  assign t[44] = (~t[56] & t[57] & t[58] & t[59]) | (t[56] & ~t[58] & ~t[59]) | (t[56] & ~t[57] & ~t[59]) | (t[56] & ~t[57] & ~t[58]);
  assign t[45] = (~t[60] & t[61] & t[62] & t[63]) | (t[60] & ~t[62] & ~t[63]) | (t[60] & ~t[61] & ~t[63]) | (t[60] & ~t[61] & ~t[62]);
  assign t[46] = (~t[64] & t[65] & t[66] & t[67]) | (t[64] & ~t[66] & ~t[67]) | (t[64] & ~t[65] & ~t[67]) | (t[64] & ~t[65] & ~t[66]);
  assign t[47] = (~t[68] & t[69] & t[70] & t[71]) | (t[68] & ~t[70] & ~t[71]) | (t[68] & ~t[69] & ~t[71]) | (t[68] & ~t[69] & ~t[70]);
  assign t[48] = (~t[72] & t[73] & t[74] & t[75]) | (t[72] & ~t[74] & ~t[75]) | (t[72] & ~t[73] & ~t[75]) | (t[72] & ~t[73] & ~t[74]);
  assign t[49] = (~t[76] & t[77] & t[78] & t[79]) | (t[76] & ~t[78] & ~t[79]) | (t[76] & ~t[77] & ~t[79]) | (t[76] & ~t[77] & ~t[78]);
  assign t[4] = ~(t[6] ^ t[25]);
  assign t[50] = (~t[80] & t[81] & t[82] & t[83]) | (t[80] & ~t[82] & ~t[83]) | (t[80] & ~t[81] & ~t[83]) | (t[80] & ~t[81] & ~t[82]);
  assign t[51] = (~t[84] & t[85] & t[86] & t[87]) | (t[84] & ~t[86] & ~t[87]) | (t[84] & ~t[85] & ~t[87]) | (t[84] & ~t[85] & ~t[86]);
  assign t[52] = t[88] ^ x[6];
  assign t[53] = t[89] ^ x[3];
  assign t[54] = t[90] ^ x[4];
  assign t[55] = t[91] ^ x[5];
  assign t[56] = t[92] ^ x[11];
  assign t[57] = t[93] ^ x[8];
  assign t[58] = t[94] ^ x[9];
  assign t[59] = t[95] ^ x[10];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[96] ^ x[16];
  assign t[61] = t[97] ^ x[13];
  assign t[62] = t[98] ^ x[14];
  assign t[63] = t[99] ^ x[15];
  assign t[64] = t[100] ^ x[21];
  assign t[65] = t[101] ^ x[18];
  assign t[66] = t[102] ^ x[19];
  assign t[67] = t[103] ^ x[20];
  assign t[68] = t[104] ^ x[26];
  assign t[69] = t[105] ^ x[23];
  assign t[6] = ~t[9];
  assign t[70] = t[106] ^ x[24];
  assign t[71] = t[107] ^ x[25];
  assign t[72] = t[108] ^ x[31];
  assign t[73] = t[109] ^ x[28];
  assign t[74] = t[110] ^ x[29];
  assign t[75] = t[111] ^ x[30];
  assign t[76] = t[112] ^ x[36];
  assign t[77] = t[113] ^ x[33];
  assign t[78] = t[114] ^ x[34];
  assign t[79] = t[115] ^ x[35];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[116] ^ x[41];
  assign t[81] = t[117] ^ x[38];
  assign t[82] = t[118] ^ x[39];
  assign t[83] = t[119] ^ x[40];
  assign t[84] = t[120] ^ x[46];
  assign t[85] = t[121] ^ x[43];
  assign t[86] = t[122] ^ x[44];
  assign t[87] = t[123] ^ x[45];
  assign t[88] = (x[2]);
  assign t[89] = (x[2]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[2]);
  assign t[91] = (x[2]);
  assign t[92] = (x[7]);
  assign t[93] = (x[7]);
  assign t[94] = (x[7]);
  assign t[95] = (x[7]);
  assign t[96] = (x[12]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[12]);
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind160(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[20] ^ t[11]);
  assign t[13] = t[22] ^ t[21];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[20] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[20] ^ t[18];
  assign t[18] = t[21] ^ t[23];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[20] & t[10];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0]);
endmodule

module R2ind161(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[20] ^ t[11]);
  assign t[13] = t[22] ^ t[21];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[20] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[20] ^ t[18];
  assign t[18] = t[21] ^ t[23];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[20] & t[10];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0]);
endmodule

module R2ind162(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[20] ^ t[11]);
  assign t[13] = t[22] ^ t[21];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[20] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[20] ^ t[18];
  assign t[18] = t[21] ^ t[23];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[20] & t[10];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0]);
endmodule

module R2ind163(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[20] ^ t[11]);
  assign t[13] = t[22] ^ t[21];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[20] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[20] ^ t[18];
  assign t[18] = t[21] ^ t[23];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[20] & t[10];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0]);
endmodule

module R2ind164(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[21] ^ t[22];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[20] ^ t[12]);
  assign t[14] = t[20] & t[16];
  assign t[15] = t[20] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[20] ^ t[10];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[20] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind165(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[21] ^ t[22];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[20] ^ t[12]);
  assign t[14] = t[20] & t[16];
  assign t[15] = t[20] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[20] ^ t[10];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[20] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind166(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[21] ^ t[22];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[20] ^ t[12]);
  assign t[14] = t[20] & t[16];
  assign t[15] = t[20] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[20] ^ t[10];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[20] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind167(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[21] ^ t[22];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[20] ^ t[12]);
  assign t[14] = t[20] & t[16];
  assign t[15] = t[20] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[20] ^ t[10];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[20] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind168(x, y);
 input [21:0] x;
 output y;

 wire [52:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[16];
  assign t[16] = t[20] ^ x[21];
  assign t[17] = (~t[21] & t[22] & t[23] & t[24]) | (t[21] & ~t[23] & ~t[24]) | (t[21] & ~t[22] & ~t[24]) | (t[21] & ~t[22] & ~t[23]);
  assign t[18] = (~t[25] & t[26] & t[27] & t[28]) | (t[25] & ~t[27] & ~t[28]) | (t[25] & ~t[26] & ~t[28]) | (t[25] & ~t[26] & ~t[27]);
  assign t[19] = (~t[29] & t[30] & t[31] & t[32]) | (t[29] & ~t[31] & ~t[32]) | (t[29] & ~t[30] & ~t[32]) | (t[29] & ~t[30] & ~t[31]);
  assign t[1] = ~(t[2] ^ t[9]);
  assign t[20] = (~t[33] & t[34] & t[35] & t[36]) | (t[33] & ~t[35] & ~t[36]) | (t[33] & ~t[34] & ~t[36]) | (t[33] & ~t[34] & ~t[35]);
  assign t[21] = t[37] ^ x[6];
  assign t[22] = t[38] ^ x[3];
  assign t[23] = t[39] ^ x[4];
  assign t[24] = t[40] ^ x[5];
  assign t[25] = t[41] ^ x[11];
  assign t[26] = t[42] ^ x[8];
  assign t[27] = t[43] ^ x[9];
  assign t[28] = t[44] ^ x[10];
  assign t[29] = t[45] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[46] ^ x[13];
  assign t[31] = t[47] ^ x[14];
  assign t[32] = t[48] ^ x[15];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[18];
  assign t[35] = t[51] ^ x[19];
  assign t[36] = t[52] ^ x[20];
  assign t[37] = (x[2]);
  assign t[38] = (x[2]);
  assign t[39] = (x[2]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[2]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[7]);
  assign t[45] = (x[12]);
  assign t[46] = (x[12]);
  assign t[47] = (x[12]);
  assign t[48] = (x[12]);
  assign t[49] = (x[17]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[52] = (x[17]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[12] ^ t[7]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind169(x, y);
 input [21:0] x;
 output y;

 wire [52:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[16];
  assign t[16] = t[20] ^ x[21];
  assign t[17] = (~t[21] & t[22] & t[23] & t[24]) | (t[21] & ~t[23] & ~t[24]) | (t[21] & ~t[22] & ~t[24]) | (t[21] & ~t[22] & ~t[23]);
  assign t[18] = (~t[25] & t[26] & t[27] & t[28]) | (t[25] & ~t[27] & ~t[28]) | (t[25] & ~t[26] & ~t[28]) | (t[25] & ~t[26] & ~t[27]);
  assign t[19] = (~t[29] & t[30] & t[31] & t[32]) | (t[29] & ~t[31] & ~t[32]) | (t[29] & ~t[30] & ~t[32]) | (t[29] & ~t[30] & ~t[31]);
  assign t[1] = ~(t[2] ^ t[9]);
  assign t[20] = (~t[33] & t[34] & t[35] & t[36]) | (t[33] & ~t[35] & ~t[36]) | (t[33] & ~t[34] & ~t[36]) | (t[33] & ~t[34] & ~t[35]);
  assign t[21] = t[37] ^ x[6];
  assign t[22] = t[38] ^ x[3];
  assign t[23] = t[39] ^ x[4];
  assign t[24] = t[40] ^ x[5];
  assign t[25] = t[41] ^ x[11];
  assign t[26] = t[42] ^ x[8];
  assign t[27] = t[43] ^ x[9];
  assign t[28] = t[44] ^ x[10];
  assign t[29] = t[45] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[46] ^ x[13];
  assign t[31] = t[47] ^ x[14];
  assign t[32] = t[48] ^ x[15];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[18];
  assign t[35] = t[51] ^ x[19];
  assign t[36] = t[52] ^ x[20];
  assign t[37] = (x[2]);
  assign t[38] = (x[2]);
  assign t[39] = (x[2]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[2]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[7]);
  assign t[45] = (x[12]);
  assign t[46] = (x[12]);
  assign t[47] = (x[12]);
  assign t[48] = (x[12]);
  assign t[49] = (x[17]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[52] = (x[17]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[12] ^ t[7]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind170(x, y);
 input [21:0] x;
 output y;

 wire [52:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[16];
  assign t[16] = t[20] ^ x[21];
  assign t[17] = (~t[21] & t[22] & t[23] & t[24]) | (t[21] & ~t[23] & ~t[24]) | (t[21] & ~t[22] & ~t[24]) | (t[21] & ~t[22] & ~t[23]);
  assign t[18] = (~t[25] & t[26] & t[27] & t[28]) | (t[25] & ~t[27] & ~t[28]) | (t[25] & ~t[26] & ~t[28]) | (t[25] & ~t[26] & ~t[27]);
  assign t[19] = (~t[29] & t[30] & t[31] & t[32]) | (t[29] & ~t[31] & ~t[32]) | (t[29] & ~t[30] & ~t[32]) | (t[29] & ~t[30] & ~t[31]);
  assign t[1] = ~(t[2] ^ t[9]);
  assign t[20] = (~t[33] & t[34] & t[35] & t[36]) | (t[33] & ~t[35] & ~t[36]) | (t[33] & ~t[34] & ~t[36]) | (t[33] & ~t[34] & ~t[35]);
  assign t[21] = t[37] ^ x[6];
  assign t[22] = t[38] ^ x[3];
  assign t[23] = t[39] ^ x[4];
  assign t[24] = t[40] ^ x[5];
  assign t[25] = t[41] ^ x[11];
  assign t[26] = t[42] ^ x[8];
  assign t[27] = t[43] ^ x[9];
  assign t[28] = t[44] ^ x[10];
  assign t[29] = t[45] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[46] ^ x[13];
  assign t[31] = t[47] ^ x[14];
  assign t[32] = t[48] ^ x[15];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[18];
  assign t[35] = t[51] ^ x[19];
  assign t[36] = t[52] ^ x[20];
  assign t[37] = (x[2]);
  assign t[38] = (x[2]);
  assign t[39] = (x[2]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[2]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[7]);
  assign t[45] = (x[12]);
  assign t[46] = (x[12]);
  assign t[47] = (x[12]);
  assign t[48] = (x[12]);
  assign t[49] = (x[17]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[52] = (x[17]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[12] ^ t[7]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind171(x, y);
 input [21:0] x;
 output y;

 wire [52:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[16];
  assign t[16] = t[20] ^ x[21];
  assign t[17] = (~t[21] & t[22] & t[23] & t[24]) | (t[21] & ~t[23] & ~t[24]) | (t[21] & ~t[22] & ~t[24]) | (t[21] & ~t[22] & ~t[23]);
  assign t[18] = (~t[25] & t[26] & t[27] & t[28]) | (t[25] & ~t[27] & ~t[28]) | (t[25] & ~t[26] & ~t[28]) | (t[25] & ~t[26] & ~t[27]);
  assign t[19] = (~t[29] & t[30] & t[31] & t[32]) | (t[29] & ~t[31] & ~t[32]) | (t[29] & ~t[30] & ~t[32]) | (t[29] & ~t[30] & ~t[31]);
  assign t[1] = ~(t[2] ^ t[9]);
  assign t[20] = (~t[33] & t[34] & t[35] & t[36]) | (t[33] & ~t[35] & ~t[36]) | (t[33] & ~t[34] & ~t[36]) | (t[33] & ~t[34] & ~t[35]);
  assign t[21] = t[37] ^ x[6];
  assign t[22] = t[38] ^ x[3];
  assign t[23] = t[39] ^ x[4];
  assign t[24] = t[40] ^ x[5];
  assign t[25] = t[41] ^ x[11];
  assign t[26] = t[42] ^ x[8];
  assign t[27] = t[43] ^ x[9];
  assign t[28] = t[44] ^ x[10];
  assign t[29] = t[45] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[46] ^ x[13];
  assign t[31] = t[47] ^ x[14];
  assign t[32] = t[48] ^ x[15];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[18];
  assign t[35] = t[51] ^ x[19];
  assign t[36] = t[52] ^ x[20];
  assign t[37] = (x[2]);
  assign t[38] = (x[2]);
  assign t[39] = (x[2]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[2]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[7]);
  assign t[45] = (x[12]);
  assign t[46] = (x[12]);
  assign t[47] = (x[12]);
  assign t[48] = (x[12]);
  assign t[49] = (x[17]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[52] = (x[17]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[12] ^ t[7]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind172(x, y);
 input [26:0] x;
 output y;

 wire [67:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] ^ t[12];
  assign t[12] = t[15] ^ t[17];
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~(t[2] ^ t[13]);
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[24] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[25] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[26] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[27] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[28] = t[48] ^ x[6];
  assign t[29] = t[49] ^ x[3];
  assign t[2] = ~t[3];
  assign t[30] = t[50] ^ x[4];
  assign t[31] = t[51] ^ x[5];
  assign t[32] = t[52] ^ x[11];
  assign t[33] = t[53] ^ x[8];
  assign t[34] = t[54] ^ x[9];
  assign t[35] = t[55] ^ x[10];
  assign t[36] = t[56] ^ x[16];
  assign t[37] = t[57] ^ x[13];
  assign t[38] = t[58] ^ x[14];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[4]);
  assign t[40] = t[60] ^ x[21];
  assign t[41] = t[61] ^ x[18];
  assign t[42] = t[62] ^ x[19];
  assign t[43] = t[63] ^ x[20];
  assign t[44] = t[64] ^ x[26];
  assign t[45] = t[65] ^ x[23];
  assign t[46] = t[66] ^ x[24];
  assign t[47] = t[67] ^ x[25];
  assign t[48] = (x[2]);
  assign t[49] = (x[2]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[2]);
  assign t[51] = (x[2]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[7]);
  assign t[55] = (x[7]);
  assign t[56] = (x[12]);
  assign t[57] = (x[12]);
  assign t[58] = (x[12]);
  assign t[59] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[60] = (x[17]);
  assign t[61] = (x[17]);
  assign t[62] = (x[17]);
  assign t[63] = (x[17]);
  assign t[64] = (x[22]);
  assign t[65] = (x[22]);
  assign t[66] = (x[22]);
  assign t[67] = (x[22]);
  assign t[6] = t[9] & t[10];
  assign t[7] = t[14] ^ t[15];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind173(x, y);
 input [26:0] x;
 output y;

 wire [67:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] ^ t[12];
  assign t[12] = t[15] ^ t[17];
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~(t[2] ^ t[13]);
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[24] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[25] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[26] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[27] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[28] = t[48] ^ x[6];
  assign t[29] = t[49] ^ x[3];
  assign t[2] = ~t[3];
  assign t[30] = t[50] ^ x[4];
  assign t[31] = t[51] ^ x[5];
  assign t[32] = t[52] ^ x[11];
  assign t[33] = t[53] ^ x[8];
  assign t[34] = t[54] ^ x[9];
  assign t[35] = t[55] ^ x[10];
  assign t[36] = t[56] ^ x[16];
  assign t[37] = t[57] ^ x[13];
  assign t[38] = t[58] ^ x[14];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[4]);
  assign t[40] = t[60] ^ x[21];
  assign t[41] = t[61] ^ x[18];
  assign t[42] = t[62] ^ x[19];
  assign t[43] = t[63] ^ x[20];
  assign t[44] = t[64] ^ x[26];
  assign t[45] = t[65] ^ x[23];
  assign t[46] = t[66] ^ x[24];
  assign t[47] = t[67] ^ x[25];
  assign t[48] = (x[2]);
  assign t[49] = (x[2]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[2]);
  assign t[51] = (x[2]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[7]);
  assign t[55] = (x[7]);
  assign t[56] = (x[12]);
  assign t[57] = (x[12]);
  assign t[58] = (x[12]);
  assign t[59] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[60] = (x[17]);
  assign t[61] = (x[17]);
  assign t[62] = (x[17]);
  assign t[63] = (x[17]);
  assign t[64] = (x[22]);
  assign t[65] = (x[22]);
  assign t[66] = (x[22]);
  assign t[67] = (x[22]);
  assign t[6] = t[9] & t[10];
  assign t[7] = t[14] ^ t[15];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind174(x, y);
 input [26:0] x;
 output y;

 wire [67:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] ^ t[12];
  assign t[12] = t[15] ^ t[17];
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~(t[2] ^ t[13]);
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[24] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[25] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[26] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[27] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[28] = t[48] ^ x[6];
  assign t[29] = t[49] ^ x[3];
  assign t[2] = ~t[3];
  assign t[30] = t[50] ^ x[4];
  assign t[31] = t[51] ^ x[5];
  assign t[32] = t[52] ^ x[11];
  assign t[33] = t[53] ^ x[8];
  assign t[34] = t[54] ^ x[9];
  assign t[35] = t[55] ^ x[10];
  assign t[36] = t[56] ^ x[16];
  assign t[37] = t[57] ^ x[13];
  assign t[38] = t[58] ^ x[14];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[4]);
  assign t[40] = t[60] ^ x[21];
  assign t[41] = t[61] ^ x[18];
  assign t[42] = t[62] ^ x[19];
  assign t[43] = t[63] ^ x[20];
  assign t[44] = t[64] ^ x[26];
  assign t[45] = t[65] ^ x[23];
  assign t[46] = t[66] ^ x[24];
  assign t[47] = t[67] ^ x[25];
  assign t[48] = (x[2]);
  assign t[49] = (x[2]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[2]);
  assign t[51] = (x[2]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[7]);
  assign t[55] = (x[7]);
  assign t[56] = (x[12]);
  assign t[57] = (x[12]);
  assign t[58] = (x[12]);
  assign t[59] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[60] = (x[17]);
  assign t[61] = (x[17]);
  assign t[62] = (x[17]);
  assign t[63] = (x[17]);
  assign t[64] = (x[22]);
  assign t[65] = (x[22]);
  assign t[66] = (x[22]);
  assign t[67] = (x[22]);
  assign t[6] = t[9] & t[10];
  assign t[7] = t[14] ^ t[15];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind175(x, y);
 input [26:0] x;
 output y;

 wire [67:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] ^ t[12];
  assign t[12] = t[15] ^ t[17];
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~(t[2] ^ t[13]);
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[24] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[25] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[26] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[27] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[28] = t[48] ^ x[6];
  assign t[29] = t[49] ^ x[3];
  assign t[2] = ~t[3];
  assign t[30] = t[50] ^ x[4];
  assign t[31] = t[51] ^ x[5];
  assign t[32] = t[52] ^ x[11];
  assign t[33] = t[53] ^ x[8];
  assign t[34] = t[54] ^ x[9];
  assign t[35] = t[55] ^ x[10];
  assign t[36] = t[56] ^ x[16];
  assign t[37] = t[57] ^ x[13];
  assign t[38] = t[58] ^ x[14];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[4]);
  assign t[40] = t[60] ^ x[21];
  assign t[41] = t[61] ^ x[18];
  assign t[42] = t[62] ^ x[19];
  assign t[43] = t[63] ^ x[20];
  assign t[44] = t[64] ^ x[26];
  assign t[45] = t[65] ^ x[23];
  assign t[46] = t[66] ^ x[24];
  assign t[47] = t[67] ^ x[25];
  assign t[48] = (x[2]);
  assign t[49] = (x[2]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[2]);
  assign t[51] = (x[2]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[7]);
  assign t[55] = (x[7]);
  assign t[56] = (x[12]);
  assign t[57] = (x[12]);
  assign t[58] = (x[12]);
  assign t[59] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[60] = (x[17]);
  assign t[61] = (x[17]);
  assign t[62] = (x[17]);
  assign t[63] = (x[17]);
  assign t[64] = (x[22]);
  assign t[65] = (x[22]);
  assign t[66] = (x[22]);
  assign t[67] = (x[22]);
  assign t[6] = t[9] & t[10];
  assign t[7] = t[14] ^ t[15];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind176(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[20] ^ t[11]);
  assign t[13] = t[22] ^ t[21];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[20] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[20] ^ t[18];
  assign t[18] = t[21] ^ t[23];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[20] & t[10];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0]);
endmodule

module R2ind177(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[20] ^ t[11]);
  assign t[13] = t[22] ^ t[21];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[20] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[20] ^ t[18];
  assign t[18] = t[21] ^ t[23];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[20] & t[10];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0]);
endmodule

module R2ind178(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[20] ^ t[11]);
  assign t[13] = t[22] ^ t[21];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[20] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[20] ^ t[18];
  assign t[18] = t[21] ^ t[23];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[20] & t[10];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0]);
endmodule

module R2ind179(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[20] ^ t[11]);
  assign t[13] = t[22] ^ t[21];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[20] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[20] ^ t[18];
  assign t[18] = t[21] ^ t[23];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[20] & t[10];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0]);
endmodule

module R2ind180(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[21] ^ t[22];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[20] ^ t[12]);
  assign t[14] = t[20] & t[16];
  assign t[15] = t[20] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[20] ^ t[10];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[20] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind181(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[21] ^ t[22];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[20] ^ t[12]);
  assign t[14] = t[20] & t[16];
  assign t[15] = t[20] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[20] ^ t[10];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[20] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind182(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[21] ^ t[22];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[20] ^ t[12]);
  assign t[14] = t[20] & t[16];
  assign t[15] = t[20] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[20] ^ t[10];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[20] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind183(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[21] ^ t[22];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[20] ^ t[12]);
  assign t[14] = t[20] & t[16];
  assign t[15] = t[20] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[20] ^ t[10];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[20] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind184(x, y);
 input [21:0] x;
 output y;

 wire [52:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[16];
  assign t[16] = t[20] ^ x[21];
  assign t[17] = (~t[21] & t[22] & t[23] & t[24]) | (t[21] & ~t[23] & ~t[24]) | (t[21] & ~t[22] & ~t[24]) | (t[21] & ~t[22] & ~t[23]);
  assign t[18] = (~t[25] & t[26] & t[27] & t[28]) | (t[25] & ~t[27] & ~t[28]) | (t[25] & ~t[26] & ~t[28]) | (t[25] & ~t[26] & ~t[27]);
  assign t[19] = (~t[29] & t[30] & t[31] & t[32]) | (t[29] & ~t[31] & ~t[32]) | (t[29] & ~t[30] & ~t[32]) | (t[29] & ~t[30] & ~t[31]);
  assign t[1] = ~(t[2] ^ t[9]);
  assign t[20] = (~t[33] & t[34] & t[35] & t[36]) | (t[33] & ~t[35] & ~t[36]) | (t[33] & ~t[34] & ~t[36]) | (t[33] & ~t[34] & ~t[35]);
  assign t[21] = t[37] ^ x[6];
  assign t[22] = t[38] ^ x[3];
  assign t[23] = t[39] ^ x[4];
  assign t[24] = t[40] ^ x[5];
  assign t[25] = t[41] ^ x[11];
  assign t[26] = t[42] ^ x[8];
  assign t[27] = t[43] ^ x[9];
  assign t[28] = t[44] ^ x[10];
  assign t[29] = t[45] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[46] ^ x[13];
  assign t[31] = t[47] ^ x[14];
  assign t[32] = t[48] ^ x[15];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[18];
  assign t[35] = t[51] ^ x[19];
  assign t[36] = t[52] ^ x[20];
  assign t[37] = (x[2]);
  assign t[38] = (x[2]);
  assign t[39] = (x[2]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[2]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[7]);
  assign t[45] = (x[12]);
  assign t[46] = (x[12]);
  assign t[47] = (x[12]);
  assign t[48] = (x[12]);
  assign t[49] = (x[17]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[52] = (x[17]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[12] ^ t[7]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind185(x, y);
 input [21:0] x;
 output y;

 wire [52:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[16];
  assign t[16] = t[20] ^ x[21];
  assign t[17] = (~t[21] & t[22] & t[23] & t[24]) | (t[21] & ~t[23] & ~t[24]) | (t[21] & ~t[22] & ~t[24]) | (t[21] & ~t[22] & ~t[23]);
  assign t[18] = (~t[25] & t[26] & t[27] & t[28]) | (t[25] & ~t[27] & ~t[28]) | (t[25] & ~t[26] & ~t[28]) | (t[25] & ~t[26] & ~t[27]);
  assign t[19] = (~t[29] & t[30] & t[31] & t[32]) | (t[29] & ~t[31] & ~t[32]) | (t[29] & ~t[30] & ~t[32]) | (t[29] & ~t[30] & ~t[31]);
  assign t[1] = ~(t[2] ^ t[9]);
  assign t[20] = (~t[33] & t[34] & t[35] & t[36]) | (t[33] & ~t[35] & ~t[36]) | (t[33] & ~t[34] & ~t[36]) | (t[33] & ~t[34] & ~t[35]);
  assign t[21] = t[37] ^ x[6];
  assign t[22] = t[38] ^ x[3];
  assign t[23] = t[39] ^ x[4];
  assign t[24] = t[40] ^ x[5];
  assign t[25] = t[41] ^ x[11];
  assign t[26] = t[42] ^ x[8];
  assign t[27] = t[43] ^ x[9];
  assign t[28] = t[44] ^ x[10];
  assign t[29] = t[45] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[46] ^ x[13];
  assign t[31] = t[47] ^ x[14];
  assign t[32] = t[48] ^ x[15];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[18];
  assign t[35] = t[51] ^ x[19];
  assign t[36] = t[52] ^ x[20];
  assign t[37] = (x[2]);
  assign t[38] = (x[2]);
  assign t[39] = (x[2]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[2]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[7]);
  assign t[45] = (x[12]);
  assign t[46] = (x[12]);
  assign t[47] = (x[12]);
  assign t[48] = (x[12]);
  assign t[49] = (x[17]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[52] = (x[17]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[12] ^ t[7]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind186(x, y);
 input [21:0] x;
 output y;

 wire [52:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[16];
  assign t[16] = t[20] ^ x[21];
  assign t[17] = (~t[21] & t[22] & t[23] & t[24]) | (t[21] & ~t[23] & ~t[24]) | (t[21] & ~t[22] & ~t[24]) | (t[21] & ~t[22] & ~t[23]);
  assign t[18] = (~t[25] & t[26] & t[27] & t[28]) | (t[25] & ~t[27] & ~t[28]) | (t[25] & ~t[26] & ~t[28]) | (t[25] & ~t[26] & ~t[27]);
  assign t[19] = (~t[29] & t[30] & t[31] & t[32]) | (t[29] & ~t[31] & ~t[32]) | (t[29] & ~t[30] & ~t[32]) | (t[29] & ~t[30] & ~t[31]);
  assign t[1] = ~(t[2] ^ t[9]);
  assign t[20] = (~t[33] & t[34] & t[35] & t[36]) | (t[33] & ~t[35] & ~t[36]) | (t[33] & ~t[34] & ~t[36]) | (t[33] & ~t[34] & ~t[35]);
  assign t[21] = t[37] ^ x[6];
  assign t[22] = t[38] ^ x[3];
  assign t[23] = t[39] ^ x[4];
  assign t[24] = t[40] ^ x[5];
  assign t[25] = t[41] ^ x[11];
  assign t[26] = t[42] ^ x[8];
  assign t[27] = t[43] ^ x[9];
  assign t[28] = t[44] ^ x[10];
  assign t[29] = t[45] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[46] ^ x[13];
  assign t[31] = t[47] ^ x[14];
  assign t[32] = t[48] ^ x[15];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[18];
  assign t[35] = t[51] ^ x[19];
  assign t[36] = t[52] ^ x[20];
  assign t[37] = (x[2]);
  assign t[38] = (x[2]);
  assign t[39] = (x[2]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[2]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[7]);
  assign t[45] = (x[12]);
  assign t[46] = (x[12]);
  assign t[47] = (x[12]);
  assign t[48] = (x[12]);
  assign t[49] = (x[17]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[52] = (x[17]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[12] ^ t[7]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind187(x, y);
 input [21:0] x;
 output y;

 wire [52:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[16];
  assign t[16] = t[20] ^ x[21];
  assign t[17] = (~t[21] & t[22] & t[23] & t[24]) | (t[21] & ~t[23] & ~t[24]) | (t[21] & ~t[22] & ~t[24]) | (t[21] & ~t[22] & ~t[23]);
  assign t[18] = (~t[25] & t[26] & t[27] & t[28]) | (t[25] & ~t[27] & ~t[28]) | (t[25] & ~t[26] & ~t[28]) | (t[25] & ~t[26] & ~t[27]);
  assign t[19] = (~t[29] & t[30] & t[31] & t[32]) | (t[29] & ~t[31] & ~t[32]) | (t[29] & ~t[30] & ~t[32]) | (t[29] & ~t[30] & ~t[31]);
  assign t[1] = ~(t[2] ^ t[9]);
  assign t[20] = (~t[33] & t[34] & t[35] & t[36]) | (t[33] & ~t[35] & ~t[36]) | (t[33] & ~t[34] & ~t[36]) | (t[33] & ~t[34] & ~t[35]);
  assign t[21] = t[37] ^ x[6];
  assign t[22] = t[38] ^ x[3];
  assign t[23] = t[39] ^ x[4];
  assign t[24] = t[40] ^ x[5];
  assign t[25] = t[41] ^ x[11];
  assign t[26] = t[42] ^ x[8];
  assign t[27] = t[43] ^ x[9];
  assign t[28] = t[44] ^ x[10];
  assign t[29] = t[45] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[46] ^ x[13];
  assign t[31] = t[47] ^ x[14];
  assign t[32] = t[48] ^ x[15];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[18];
  assign t[35] = t[51] ^ x[19];
  assign t[36] = t[52] ^ x[20];
  assign t[37] = (x[2]);
  assign t[38] = (x[2]);
  assign t[39] = (x[2]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[2]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[7]);
  assign t[45] = (x[12]);
  assign t[46] = (x[12]);
  assign t[47] = (x[12]);
  assign t[48] = (x[12]);
  assign t[49] = (x[17]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[52] = (x[17]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[12] ^ t[7]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind188(x, y);
 input [26:0] x;
 output y;

 wire [67:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] ^ t[12];
  assign t[12] = t[15] ^ t[17];
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~(t[2] ^ t[13]);
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[24] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[25] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[26] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[27] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[28] = t[48] ^ x[6];
  assign t[29] = t[49] ^ x[3];
  assign t[2] = ~t[3];
  assign t[30] = t[50] ^ x[4];
  assign t[31] = t[51] ^ x[5];
  assign t[32] = t[52] ^ x[11];
  assign t[33] = t[53] ^ x[8];
  assign t[34] = t[54] ^ x[9];
  assign t[35] = t[55] ^ x[10];
  assign t[36] = t[56] ^ x[16];
  assign t[37] = t[57] ^ x[13];
  assign t[38] = t[58] ^ x[14];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[4]);
  assign t[40] = t[60] ^ x[21];
  assign t[41] = t[61] ^ x[18];
  assign t[42] = t[62] ^ x[19];
  assign t[43] = t[63] ^ x[20];
  assign t[44] = t[64] ^ x[26];
  assign t[45] = t[65] ^ x[23];
  assign t[46] = t[66] ^ x[24];
  assign t[47] = t[67] ^ x[25];
  assign t[48] = (x[2]);
  assign t[49] = (x[2]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[2]);
  assign t[51] = (x[2]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[7]);
  assign t[55] = (x[7]);
  assign t[56] = (x[12]);
  assign t[57] = (x[12]);
  assign t[58] = (x[12]);
  assign t[59] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[60] = (x[17]);
  assign t[61] = (x[17]);
  assign t[62] = (x[17]);
  assign t[63] = (x[17]);
  assign t[64] = (x[22]);
  assign t[65] = (x[22]);
  assign t[66] = (x[22]);
  assign t[67] = (x[22]);
  assign t[6] = t[9] & t[10];
  assign t[7] = t[14] ^ t[15];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind189(x, y);
 input [26:0] x;
 output y;

 wire [67:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] ^ t[12];
  assign t[12] = t[15] ^ t[17];
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~(t[2] ^ t[13]);
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[24] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[25] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[26] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[27] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[28] = t[48] ^ x[6];
  assign t[29] = t[49] ^ x[3];
  assign t[2] = ~t[3];
  assign t[30] = t[50] ^ x[4];
  assign t[31] = t[51] ^ x[5];
  assign t[32] = t[52] ^ x[11];
  assign t[33] = t[53] ^ x[8];
  assign t[34] = t[54] ^ x[9];
  assign t[35] = t[55] ^ x[10];
  assign t[36] = t[56] ^ x[16];
  assign t[37] = t[57] ^ x[13];
  assign t[38] = t[58] ^ x[14];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[4]);
  assign t[40] = t[60] ^ x[21];
  assign t[41] = t[61] ^ x[18];
  assign t[42] = t[62] ^ x[19];
  assign t[43] = t[63] ^ x[20];
  assign t[44] = t[64] ^ x[26];
  assign t[45] = t[65] ^ x[23];
  assign t[46] = t[66] ^ x[24];
  assign t[47] = t[67] ^ x[25];
  assign t[48] = (x[2]);
  assign t[49] = (x[2]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[2]);
  assign t[51] = (x[2]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[7]);
  assign t[55] = (x[7]);
  assign t[56] = (x[12]);
  assign t[57] = (x[12]);
  assign t[58] = (x[12]);
  assign t[59] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[60] = (x[17]);
  assign t[61] = (x[17]);
  assign t[62] = (x[17]);
  assign t[63] = (x[17]);
  assign t[64] = (x[22]);
  assign t[65] = (x[22]);
  assign t[66] = (x[22]);
  assign t[67] = (x[22]);
  assign t[6] = t[9] & t[10];
  assign t[7] = t[14] ^ t[15];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind190(x, y);
 input [26:0] x;
 output y;

 wire [67:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] ^ t[12];
  assign t[12] = t[15] ^ t[17];
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~(t[2] ^ t[13]);
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[24] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[25] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[26] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[27] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[28] = t[48] ^ x[6];
  assign t[29] = t[49] ^ x[3];
  assign t[2] = ~t[3];
  assign t[30] = t[50] ^ x[4];
  assign t[31] = t[51] ^ x[5];
  assign t[32] = t[52] ^ x[11];
  assign t[33] = t[53] ^ x[8];
  assign t[34] = t[54] ^ x[9];
  assign t[35] = t[55] ^ x[10];
  assign t[36] = t[56] ^ x[16];
  assign t[37] = t[57] ^ x[13];
  assign t[38] = t[58] ^ x[14];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[4]);
  assign t[40] = t[60] ^ x[21];
  assign t[41] = t[61] ^ x[18];
  assign t[42] = t[62] ^ x[19];
  assign t[43] = t[63] ^ x[20];
  assign t[44] = t[64] ^ x[26];
  assign t[45] = t[65] ^ x[23];
  assign t[46] = t[66] ^ x[24];
  assign t[47] = t[67] ^ x[25];
  assign t[48] = (x[2]);
  assign t[49] = (x[2]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[2]);
  assign t[51] = (x[2]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[7]);
  assign t[55] = (x[7]);
  assign t[56] = (x[12]);
  assign t[57] = (x[12]);
  assign t[58] = (x[12]);
  assign t[59] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[60] = (x[17]);
  assign t[61] = (x[17]);
  assign t[62] = (x[17]);
  assign t[63] = (x[17]);
  assign t[64] = (x[22]);
  assign t[65] = (x[22]);
  assign t[66] = (x[22]);
  assign t[67] = (x[22]);
  assign t[6] = t[9] & t[10];
  assign t[7] = t[14] ^ t[15];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind191(x, y);
 input [26:0] x;
 output y;

 wire [67:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] ^ t[12];
  assign t[12] = t[15] ^ t[17];
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~(t[2] ^ t[13]);
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[24] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[25] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[26] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[27] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[28] = t[48] ^ x[6];
  assign t[29] = t[49] ^ x[3];
  assign t[2] = ~t[3];
  assign t[30] = t[50] ^ x[4];
  assign t[31] = t[51] ^ x[5];
  assign t[32] = t[52] ^ x[11];
  assign t[33] = t[53] ^ x[8];
  assign t[34] = t[54] ^ x[9];
  assign t[35] = t[55] ^ x[10];
  assign t[36] = t[56] ^ x[16];
  assign t[37] = t[57] ^ x[13];
  assign t[38] = t[58] ^ x[14];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[4]);
  assign t[40] = t[60] ^ x[21];
  assign t[41] = t[61] ^ x[18];
  assign t[42] = t[62] ^ x[19];
  assign t[43] = t[63] ^ x[20];
  assign t[44] = t[64] ^ x[26];
  assign t[45] = t[65] ^ x[23];
  assign t[46] = t[66] ^ x[24];
  assign t[47] = t[67] ^ x[25];
  assign t[48] = (x[2]);
  assign t[49] = (x[2]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[2]);
  assign t[51] = (x[2]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[7]);
  assign t[55] = (x[7]);
  assign t[56] = (x[12]);
  assign t[57] = (x[12]);
  assign t[58] = (x[12]);
  assign t[59] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[60] = (x[17]);
  assign t[61] = (x[17]);
  assign t[62] = (x[17]);
  assign t[63] = (x[17]);
  assign t[64] = (x[22]);
  assign t[65] = (x[22]);
  assign t[66] = (x[22]);
  assign t[67] = (x[22]);
  assign t[6] = t[9] & t[10];
  assign t[7] = t[14] ^ t[15];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind192(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[20] ^ t[11]);
  assign t[13] = t[22] ^ t[21];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[20] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[20] ^ t[18];
  assign t[18] = t[21] ^ t[23];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[20] & t[10];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0]);
endmodule

module R2ind193(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[20] ^ t[11]);
  assign t[13] = t[22] ^ t[21];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[20] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[20] ^ t[18];
  assign t[18] = t[21] ^ t[23];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[20] & t[10];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0]);
endmodule

module R2ind194(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[20] ^ t[11]);
  assign t[13] = t[22] ^ t[21];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[20] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[20] ^ t[18];
  assign t[18] = t[21] ^ t[23];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[20] & t[10];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0]);
endmodule

module R2ind195(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[20] ^ t[11]);
  assign t[13] = t[22] ^ t[21];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[20] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[20] ^ t[18];
  assign t[18] = t[21] ^ t[23];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[20] & t[10];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0]);
endmodule

module R2ind196(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[21] ^ t[22];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[20] ^ t[12]);
  assign t[14] = t[20] & t[16];
  assign t[15] = t[20] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[20] ^ t[10];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[20] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind197(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[21] ^ t[22];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[20] ^ t[12]);
  assign t[14] = t[20] & t[16];
  assign t[15] = t[20] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[20] ^ t[10];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[20] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind198(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[21] ^ t[22];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[20] ^ t[12]);
  assign t[14] = t[20] & t[16];
  assign t[15] = t[20] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[20] ^ t[10];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[20] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind199(x, y);
 input [26:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[21] ^ t[22];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[20] ^ t[12]);
  assign t[14] = t[20] & t[16];
  assign t[15] = t[20] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[20] ^ t[10];
  assign t[19] = (t[24]);
  assign t[1] = ~(t[2] ^ t[19]);
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = (t[28]);
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[11];
  assign t[26] = t[31] ^ x[16];
  assign t[27] = t[32] ^ x[21];
  assign t[28] = t[33] ^ x[26];
  assign t[29] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[31] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[32] = (~t[46] & t[47] & t[48] & t[49]) | (t[46] & ~t[48] & ~t[49]) | (t[46] & ~t[47] & ~t[49]) | (t[46] & ~t[47] & ~t[48]);
  assign t[33] = (~t[50] & t[51] & t[52] & t[53]) | (t[50] & ~t[52] & ~t[53]) | (t[50] & ~t[51] & ~t[53]) | (t[50] & ~t[51] & ~t[52]);
  assign t[34] = t[54] ^ x[6];
  assign t[35] = t[55] ^ x[3];
  assign t[36] = t[56] ^ x[4];
  assign t[37] = t[57] ^ x[5];
  assign t[38] = t[58] ^ x[11];
  assign t[39] = t[59] ^ x[8];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[60] ^ x[9];
  assign t[41] = t[61] ^ x[10];
  assign t[42] = t[62] ^ x[16];
  assign t[43] = t[63] ^ x[13];
  assign t[44] = t[64] ^ x[14];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[21];
  assign t[47] = t[67] ^ x[18];
  assign t[48] = t[68] ^ x[19];
  assign t[49] = t[69] ^ x[20];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[70] ^ x[26];
  assign t[51] = t[71] ^ x[23];
  assign t[52] = t[72] ^ x[24];
  assign t[53] = t[73] ^ x[25];
  assign t[54] = (x[2]);
  assign t[55] = (x[2]);
  assign t[56] = (x[2]);
  assign t[57] = (x[2]);
  assign t[58] = (x[7]);
  assign t[59] = (x[7]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[12]);
  assign t[66] = (x[17]);
  assign t[67] = (x[17]);
  assign t[68] = (x[17]);
  assign t[69] = (x[17]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[20] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind200(x, y);
 input [21:0] x;
 output y;

 wire [52:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[16];
  assign t[16] = t[20] ^ x[21];
  assign t[17] = (~t[21] & t[22] & t[23] & t[24]) | (t[21] & ~t[23] & ~t[24]) | (t[21] & ~t[22] & ~t[24]) | (t[21] & ~t[22] & ~t[23]);
  assign t[18] = (~t[25] & t[26] & t[27] & t[28]) | (t[25] & ~t[27] & ~t[28]) | (t[25] & ~t[26] & ~t[28]) | (t[25] & ~t[26] & ~t[27]);
  assign t[19] = (~t[29] & t[30] & t[31] & t[32]) | (t[29] & ~t[31] & ~t[32]) | (t[29] & ~t[30] & ~t[32]) | (t[29] & ~t[30] & ~t[31]);
  assign t[1] = ~(t[2] ^ t[9]);
  assign t[20] = (~t[33] & t[34] & t[35] & t[36]) | (t[33] & ~t[35] & ~t[36]) | (t[33] & ~t[34] & ~t[36]) | (t[33] & ~t[34] & ~t[35]);
  assign t[21] = t[37] ^ x[6];
  assign t[22] = t[38] ^ x[3];
  assign t[23] = t[39] ^ x[4];
  assign t[24] = t[40] ^ x[5];
  assign t[25] = t[41] ^ x[11];
  assign t[26] = t[42] ^ x[8];
  assign t[27] = t[43] ^ x[9];
  assign t[28] = t[44] ^ x[10];
  assign t[29] = t[45] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[46] ^ x[13];
  assign t[31] = t[47] ^ x[14];
  assign t[32] = t[48] ^ x[15];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[18];
  assign t[35] = t[51] ^ x[19];
  assign t[36] = t[52] ^ x[20];
  assign t[37] = (x[2]);
  assign t[38] = (x[2]);
  assign t[39] = (x[2]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[2]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[7]);
  assign t[45] = (x[12]);
  assign t[46] = (x[12]);
  assign t[47] = (x[12]);
  assign t[48] = (x[12]);
  assign t[49] = (x[17]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[52] = (x[17]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[12] ^ t[7]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind201(x, y);
 input [21:0] x;
 output y;

 wire [52:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[16];
  assign t[16] = t[20] ^ x[21];
  assign t[17] = (~t[21] & t[22] & t[23] & t[24]) | (t[21] & ~t[23] & ~t[24]) | (t[21] & ~t[22] & ~t[24]) | (t[21] & ~t[22] & ~t[23]);
  assign t[18] = (~t[25] & t[26] & t[27] & t[28]) | (t[25] & ~t[27] & ~t[28]) | (t[25] & ~t[26] & ~t[28]) | (t[25] & ~t[26] & ~t[27]);
  assign t[19] = (~t[29] & t[30] & t[31] & t[32]) | (t[29] & ~t[31] & ~t[32]) | (t[29] & ~t[30] & ~t[32]) | (t[29] & ~t[30] & ~t[31]);
  assign t[1] = ~(t[2] ^ t[9]);
  assign t[20] = (~t[33] & t[34] & t[35] & t[36]) | (t[33] & ~t[35] & ~t[36]) | (t[33] & ~t[34] & ~t[36]) | (t[33] & ~t[34] & ~t[35]);
  assign t[21] = t[37] ^ x[6];
  assign t[22] = t[38] ^ x[3];
  assign t[23] = t[39] ^ x[4];
  assign t[24] = t[40] ^ x[5];
  assign t[25] = t[41] ^ x[11];
  assign t[26] = t[42] ^ x[8];
  assign t[27] = t[43] ^ x[9];
  assign t[28] = t[44] ^ x[10];
  assign t[29] = t[45] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[46] ^ x[13];
  assign t[31] = t[47] ^ x[14];
  assign t[32] = t[48] ^ x[15];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[18];
  assign t[35] = t[51] ^ x[19];
  assign t[36] = t[52] ^ x[20];
  assign t[37] = (x[2]);
  assign t[38] = (x[2]);
  assign t[39] = (x[2]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[2]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[7]);
  assign t[45] = (x[12]);
  assign t[46] = (x[12]);
  assign t[47] = (x[12]);
  assign t[48] = (x[12]);
  assign t[49] = (x[17]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[52] = (x[17]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[12] ^ t[7]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind202(x, y);
 input [21:0] x;
 output y;

 wire [52:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[16];
  assign t[16] = t[20] ^ x[21];
  assign t[17] = (~t[21] & t[22] & t[23] & t[24]) | (t[21] & ~t[23] & ~t[24]) | (t[21] & ~t[22] & ~t[24]) | (t[21] & ~t[22] & ~t[23]);
  assign t[18] = (~t[25] & t[26] & t[27] & t[28]) | (t[25] & ~t[27] & ~t[28]) | (t[25] & ~t[26] & ~t[28]) | (t[25] & ~t[26] & ~t[27]);
  assign t[19] = (~t[29] & t[30] & t[31] & t[32]) | (t[29] & ~t[31] & ~t[32]) | (t[29] & ~t[30] & ~t[32]) | (t[29] & ~t[30] & ~t[31]);
  assign t[1] = ~(t[2] ^ t[9]);
  assign t[20] = (~t[33] & t[34] & t[35] & t[36]) | (t[33] & ~t[35] & ~t[36]) | (t[33] & ~t[34] & ~t[36]) | (t[33] & ~t[34] & ~t[35]);
  assign t[21] = t[37] ^ x[6];
  assign t[22] = t[38] ^ x[3];
  assign t[23] = t[39] ^ x[4];
  assign t[24] = t[40] ^ x[5];
  assign t[25] = t[41] ^ x[11];
  assign t[26] = t[42] ^ x[8];
  assign t[27] = t[43] ^ x[9];
  assign t[28] = t[44] ^ x[10];
  assign t[29] = t[45] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[46] ^ x[13];
  assign t[31] = t[47] ^ x[14];
  assign t[32] = t[48] ^ x[15];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[18];
  assign t[35] = t[51] ^ x[19];
  assign t[36] = t[52] ^ x[20];
  assign t[37] = (x[2]);
  assign t[38] = (x[2]);
  assign t[39] = (x[2]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[2]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[7]);
  assign t[45] = (x[12]);
  assign t[46] = (x[12]);
  assign t[47] = (x[12]);
  assign t[48] = (x[12]);
  assign t[49] = (x[17]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[52] = (x[17]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[12] ^ t[7]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind203(x, y);
 input [21:0] x;
 output y;

 wire [52:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[16];
  assign t[16] = t[20] ^ x[21];
  assign t[17] = (~t[21] & t[22] & t[23] & t[24]) | (t[21] & ~t[23] & ~t[24]) | (t[21] & ~t[22] & ~t[24]) | (t[21] & ~t[22] & ~t[23]);
  assign t[18] = (~t[25] & t[26] & t[27] & t[28]) | (t[25] & ~t[27] & ~t[28]) | (t[25] & ~t[26] & ~t[28]) | (t[25] & ~t[26] & ~t[27]);
  assign t[19] = (~t[29] & t[30] & t[31] & t[32]) | (t[29] & ~t[31] & ~t[32]) | (t[29] & ~t[30] & ~t[32]) | (t[29] & ~t[30] & ~t[31]);
  assign t[1] = ~(t[2] ^ t[9]);
  assign t[20] = (~t[33] & t[34] & t[35] & t[36]) | (t[33] & ~t[35] & ~t[36]) | (t[33] & ~t[34] & ~t[36]) | (t[33] & ~t[34] & ~t[35]);
  assign t[21] = t[37] ^ x[6];
  assign t[22] = t[38] ^ x[3];
  assign t[23] = t[39] ^ x[4];
  assign t[24] = t[40] ^ x[5];
  assign t[25] = t[41] ^ x[11];
  assign t[26] = t[42] ^ x[8];
  assign t[27] = t[43] ^ x[9];
  assign t[28] = t[44] ^ x[10];
  assign t[29] = t[45] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[46] ^ x[13];
  assign t[31] = t[47] ^ x[14];
  assign t[32] = t[48] ^ x[15];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[18];
  assign t[35] = t[51] ^ x[19];
  assign t[36] = t[52] ^ x[20];
  assign t[37] = (x[2]);
  assign t[38] = (x[2]);
  assign t[39] = (x[2]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[2]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[7]);
  assign t[45] = (x[12]);
  assign t[46] = (x[12]);
  assign t[47] = (x[12]);
  assign t[48] = (x[12]);
  assign t[49] = (x[17]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[52] = (x[17]);
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[12] ^ t[7]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind204(x, y);
 input [26:0] x;
 output y;

 wire [67:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] ^ t[12];
  assign t[12] = t[15] ^ t[17];
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~(t[2] ^ t[13]);
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[24] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[25] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[26] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[27] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[28] = t[48] ^ x[6];
  assign t[29] = t[49] ^ x[3];
  assign t[2] = ~t[3];
  assign t[30] = t[50] ^ x[4];
  assign t[31] = t[51] ^ x[5];
  assign t[32] = t[52] ^ x[11];
  assign t[33] = t[53] ^ x[8];
  assign t[34] = t[54] ^ x[9];
  assign t[35] = t[55] ^ x[10];
  assign t[36] = t[56] ^ x[16];
  assign t[37] = t[57] ^ x[13];
  assign t[38] = t[58] ^ x[14];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[4]);
  assign t[40] = t[60] ^ x[21];
  assign t[41] = t[61] ^ x[18];
  assign t[42] = t[62] ^ x[19];
  assign t[43] = t[63] ^ x[20];
  assign t[44] = t[64] ^ x[26];
  assign t[45] = t[65] ^ x[23];
  assign t[46] = t[66] ^ x[24];
  assign t[47] = t[67] ^ x[25];
  assign t[48] = (x[2]);
  assign t[49] = (x[2]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[2]);
  assign t[51] = (x[2]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[7]);
  assign t[55] = (x[7]);
  assign t[56] = (x[12]);
  assign t[57] = (x[12]);
  assign t[58] = (x[12]);
  assign t[59] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[60] = (x[17]);
  assign t[61] = (x[17]);
  assign t[62] = (x[17]);
  assign t[63] = (x[17]);
  assign t[64] = (x[22]);
  assign t[65] = (x[22]);
  assign t[66] = (x[22]);
  assign t[67] = (x[22]);
  assign t[6] = t[9] & t[10];
  assign t[7] = t[14] ^ t[15];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind205(x, y);
 input [26:0] x;
 output y;

 wire [67:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] ^ t[12];
  assign t[12] = t[15] ^ t[17];
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~(t[2] ^ t[13]);
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[24] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[25] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[26] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[27] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[28] = t[48] ^ x[6];
  assign t[29] = t[49] ^ x[3];
  assign t[2] = ~t[3];
  assign t[30] = t[50] ^ x[4];
  assign t[31] = t[51] ^ x[5];
  assign t[32] = t[52] ^ x[11];
  assign t[33] = t[53] ^ x[8];
  assign t[34] = t[54] ^ x[9];
  assign t[35] = t[55] ^ x[10];
  assign t[36] = t[56] ^ x[16];
  assign t[37] = t[57] ^ x[13];
  assign t[38] = t[58] ^ x[14];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[4]);
  assign t[40] = t[60] ^ x[21];
  assign t[41] = t[61] ^ x[18];
  assign t[42] = t[62] ^ x[19];
  assign t[43] = t[63] ^ x[20];
  assign t[44] = t[64] ^ x[26];
  assign t[45] = t[65] ^ x[23];
  assign t[46] = t[66] ^ x[24];
  assign t[47] = t[67] ^ x[25];
  assign t[48] = (x[2]);
  assign t[49] = (x[2]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[2]);
  assign t[51] = (x[2]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[7]);
  assign t[55] = (x[7]);
  assign t[56] = (x[12]);
  assign t[57] = (x[12]);
  assign t[58] = (x[12]);
  assign t[59] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[60] = (x[17]);
  assign t[61] = (x[17]);
  assign t[62] = (x[17]);
  assign t[63] = (x[17]);
  assign t[64] = (x[22]);
  assign t[65] = (x[22]);
  assign t[66] = (x[22]);
  assign t[67] = (x[22]);
  assign t[6] = t[9] & t[10];
  assign t[7] = t[14] ^ t[15];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind206(x, y);
 input [26:0] x;
 output y;

 wire [67:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] ^ t[12];
  assign t[12] = t[15] ^ t[17];
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~(t[2] ^ t[13]);
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[24] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[25] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[26] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[27] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[28] = t[48] ^ x[6];
  assign t[29] = t[49] ^ x[3];
  assign t[2] = ~t[3];
  assign t[30] = t[50] ^ x[4];
  assign t[31] = t[51] ^ x[5];
  assign t[32] = t[52] ^ x[11];
  assign t[33] = t[53] ^ x[8];
  assign t[34] = t[54] ^ x[9];
  assign t[35] = t[55] ^ x[10];
  assign t[36] = t[56] ^ x[16];
  assign t[37] = t[57] ^ x[13];
  assign t[38] = t[58] ^ x[14];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[4]);
  assign t[40] = t[60] ^ x[21];
  assign t[41] = t[61] ^ x[18];
  assign t[42] = t[62] ^ x[19];
  assign t[43] = t[63] ^ x[20];
  assign t[44] = t[64] ^ x[26];
  assign t[45] = t[65] ^ x[23];
  assign t[46] = t[66] ^ x[24];
  assign t[47] = t[67] ^ x[25];
  assign t[48] = (x[2]);
  assign t[49] = (x[2]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[2]);
  assign t[51] = (x[2]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[7]);
  assign t[55] = (x[7]);
  assign t[56] = (x[12]);
  assign t[57] = (x[12]);
  assign t[58] = (x[12]);
  assign t[59] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[60] = (x[17]);
  assign t[61] = (x[17]);
  assign t[62] = (x[17]);
  assign t[63] = (x[17]);
  assign t[64] = (x[22]);
  assign t[65] = (x[22]);
  assign t[66] = (x[22]);
  assign t[67] = (x[22]);
  assign t[6] = t[9] & t[10];
  assign t[7] = t[14] ^ t[15];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind207(x, y);
 input [26:0] x;
 output y;

 wire [67:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] ^ t[12];
  assign t[12] = t[15] ^ t[17];
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = ~(t[2] ^ t[13]);
  assign t[20] = t[25] ^ x[16];
  assign t[21] = t[26] ^ x[21];
  assign t[22] = t[27] ^ x[26];
  assign t[23] = (~t[28] & t[29] & t[30] & t[31]) | (t[28] & ~t[30] & ~t[31]) | (t[28] & ~t[29] & ~t[31]) | (t[28] & ~t[29] & ~t[30]);
  assign t[24] = (~t[32] & t[33] & t[34] & t[35]) | (t[32] & ~t[34] & ~t[35]) | (t[32] & ~t[33] & ~t[35]) | (t[32] & ~t[33] & ~t[34]);
  assign t[25] = (~t[36] & t[37] & t[38] & t[39]) | (t[36] & ~t[38] & ~t[39]) | (t[36] & ~t[37] & ~t[39]) | (t[36] & ~t[37] & ~t[38]);
  assign t[26] = (~t[40] & t[41] & t[42] & t[43]) | (t[40] & ~t[42] & ~t[43]) | (t[40] & ~t[41] & ~t[43]) | (t[40] & ~t[41] & ~t[42]);
  assign t[27] = (~t[44] & t[45] & t[46] & t[47]) | (t[44] & ~t[46] & ~t[47]) | (t[44] & ~t[45] & ~t[47]) | (t[44] & ~t[45] & ~t[46]);
  assign t[28] = t[48] ^ x[6];
  assign t[29] = t[49] ^ x[3];
  assign t[2] = ~t[3];
  assign t[30] = t[50] ^ x[4];
  assign t[31] = t[51] ^ x[5];
  assign t[32] = t[52] ^ x[11];
  assign t[33] = t[53] ^ x[8];
  assign t[34] = t[54] ^ x[9];
  assign t[35] = t[55] ^ x[10];
  assign t[36] = t[56] ^ x[16];
  assign t[37] = t[57] ^ x[13];
  assign t[38] = t[58] ^ x[14];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[4]);
  assign t[40] = t[60] ^ x[21];
  assign t[41] = t[61] ^ x[18];
  assign t[42] = t[62] ^ x[19];
  assign t[43] = t[63] ^ x[20];
  assign t[44] = t[64] ^ x[26];
  assign t[45] = t[65] ^ x[23];
  assign t[46] = t[66] ^ x[24];
  assign t[47] = t[67] ^ x[25];
  assign t[48] = (x[2]);
  assign t[49] = (x[2]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[2]);
  assign t[51] = (x[2]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[7]);
  assign t[55] = (x[7]);
  assign t[56] = (x[12]);
  assign t[57] = (x[12]);
  assign t[58] = (x[12]);
  assign t[59] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[60] = (x[17]);
  assign t[61] = (x[17]);
  assign t[62] = (x[17]);
  assign t[63] = (x[17]);
  assign t[64] = (x[22]);
  assign t[65] = (x[22]);
  assign t[66] = (x[22]);
  assign t[67] = (x[22]);
  assign t[6] = t[9] & t[10];
  assign t[7] = t[14] ^ t[15];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind208(x, y);
 input [31:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[13];
  assign t[11] = t[16] ^ t[9];
  assign t[12] = t[17] ^ t[18];
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[23] ^ t[13]);
  assign t[15] = t[25] ^ t[24];
  assign t[16] = ~(t[19] ^ t[10]);
  assign t[17] = t[23] ^ t[15];
  assign t[18] = t[13] & t[19];
  assign t[19] = t[23] ^ t[20];
  assign t[1] = ~(t[2] ^ t[21]);
  assign t[20] = t[24] ^ t[26];
  assign t[21] = (t[27]);
  assign t[22] = (t[28]);
  assign t[23] = (t[29]);
  assign t[24] = (t[30]);
  assign t[25] = (t[31]);
  assign t[26] = (t[32]);
  assign t[27] = t[33] ^ x[6];
  assign t[28] = t[34] ^ x[11];
  assign t[29] = t[35] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[36] ^ x[21];
  assign t[31] = t[37] ^ x[26];
  assign t[32] = t[38] ^ x[31];
  assign t[33] = (~t[39] & t[40] & t[41] & t[42]) | (t[39] & ~t[41] & ~t[42]) | (t[39] & ~t[40] & ~t[42]) | (t[39] & ~t[40] & ~t[41]);
  assign t[34] = (~t[43] & t[44] & t[45] & t[46]) | (t[43] & ~t[45] & ~t[46]) | (t[43] & ~t[44] & ~t[46]) | (t[43] & ~t[44] & ~t[45]);
  assign t[35] = (~t[47] & t[48] & t[49] & t[50]) | (t[47] & ~t[49] & ~t[50]) | (t[47] & ~t[48] & ~t[50]) | (t[47] & ~t[48] & ~t[49]);
  assign t[36] = (~t[51] & t[52] & t[53] & t[54]) | (t[51] & ~t[53] & ~t[54]) | (t[51] & ~t[52] & ~t[54]) | (t[51] & ~t[52] & ~t[53]);
  assign t[37] = (~t[55] & t[56] & t[57] & t[58]) | (t[55] & ~t[57] & ~t[58]) | (t[55] & ~t[56] & ~t[58]) | (t[55] & ~t[56] & ~t[57]);
  assign t[38] = (~t[59] & t[60] & t[61] & t[62]) | (t[59] & ~t[61] & ~t[62]) | (t[59] & ~t[60] & ~t[62]) | (t[59] & ~t[60] & ~t[61]);
  assign t[39] = t[63] ^ x[6];
  assign t[3] = ~(t[4] ^ t[22]);
  assign t[40] = t[64] ^ x[3];
  assign t[41] = t[65] ^ x[4];
  assign t[42] = t[66] ^ x[5];
  assign t[43] = t[67] ^ x[11];
  assign t[44] = t[68] ^ x[8];
  assign t[45] = t[69] ^ x[9];
  assign t[46] = t[70] ^ x[10];
  assign t[47] = t[71] ^ x[16];
  assign t[48] = t[72] ^ x[13];
  assign t[49] = t[73] ^ x[14];
  assign t[4] = ~t[5];
  assign t[50] = t[74] ^ x[15];
  assign t[51] = t[75] ^ x[21];
  assign t[52] = t[76] ^ x[18];
  assign t[53] = t[77] ^ x[19];
  assign t[54] = t[78] ^ x[20];
  assign t[55] = t[79] ^ x[26];
  assign t[56] = t[80] ^ x[23];
  assign t[57] = t[81] ^ x[24];
  assign t[58] = t[82] ^ x[25];
  assign t[59] = t[83] ^ x[31];
  assign t[5] = t[6] ^ t[7];
  assign t[60] = t[84] ^ x[28];
  assign t[61] = t[85] ^ x[29];
  assign t[62] = t[86] ^ x[30];
  assign t[63] = (x[2]);
  assign t[64] = (x[2]);
  assign t[65] = (x[2]);
  assign t[66] = (x[2]);
  assign t[67] = (x[7]);
  assign t[68] = (x[7]);
  assign t[69] = (x[7]);
  assign t[6] = t[8] ^ t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[12]);
  assign t[72] = (x[12]);
  assign t[73] = (x[12]);
  assign t[74] = (x[12]);
  assign t[75] = (x[17]);
  assign t[76] = (x[17]);
  assign t[77] = (x[17]);
  assign t[78] = (x[17]);
  assign t[79] = (x[22]);
  assign t[7] = t[10] & t[11];
  assign t[80] = (x[22]);
  assign t[81] = (x[22]);
  assign t[82] = (x[22]);
  assign t[83] = (x[27]);
  assign t[84] = (x[27]);
  assign t[85] = (x[27]);
  assign t[86] = (x[27]);
  assign t[8] = t[23] & t[12];
  assign t[9] = t[13] & t[14];
  assign y = (t[0]);
endmodule

module R2ind209(x, y);
 input [31:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[13];
  assign t[11] = t[16] ^ t[9];
  assign t[12] = t[17] ^ t[18];
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[23] ^ t[13]);
  assign t[15] = t[25] ^ t[24];
  assign t[16] = ~(t[19] ^ t[10]);
  assign t[17] = t[23] ^ t[15];
  assign t[18] = t[13] & t[19];
  assign t[19] = t[23] ^ t[20];
  assign t[1] = ~(t[2] ^ t[21]);
  assign t[20] = t[24] ^ t[26];
  assign t[21] = (t[27]);
  assign t[22] = (t[28]);
  assign t[23] = (t[29]);
  assign t[24] = (t[30]);
  assign t[25] = (t[31]);
  assign t[26] = (t[32]);
  assign t[27] = t[33] ^ x[6];
  assign t[28] = t[34] ^ x[11];
  assign t[29] = t[35] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[36] ^ x[21];
  assign t[31] = t[37] ^ x[26];
  assign t[32] = t[38] ^ x[31];
  assign t[33] = (~t[39] & t[40] & t[41] & t[42]) | (t[39] & ~t[41] & ~t[42]) | (t[39] & ~t[40] & ~t[42]) | (t[39] & ~t[40] & ~t[41]);
  assign t[34] = (~t[43] & t[44] & t[45] & t[46]) | (t[43] & ~t[45] & ~t[46]) | (t[43] & ~t[44] & ~t[46]) | (t[43] & ~t[44] & ~t[45]);
  assign t[35] = (~t[47] & t[48] & t[49] & t[50]) | (t[47] & ~t[49] & ~t[50]) | (t[47] & ~t[48] & ~t[50]) | (t[47] & ~t[48] & ~t[49]);
  assign t[36] = (~t[51] & t[52] & t[53] & t[54]) | (t[51] & ~t[53] & ~t[54]) | (t[51] & ~t[52] & ~t[54]) | (t[51] & ~t[52] & ~t[53]);
  assign t[37] = (~t[55] & t[56] & t[57] & t[58]) | (t[55] & ~t[57] & ~t[58]) | (t[55] & ~t[56] & ~t[58]) | (t[55] & ~t[56] & ~t[57]);
  assign t[38] = (~t[59] & t[60] & t[61] & t[62]) | (t[59] & ~t[61] & ~t[62]) | (t[59] & ~t[60] & ~t[62]) | (t[59] & ~t[60] & ~t[61]);
  assign t[39] = t[63] ^ x[6];
  assign t[3] = ~(t[4] ^ t[22]);
  assign t[40] = t[64] ^ x[3];
  assign t[41] = t[65] ^ x[4];
  assign t[42] = t[66] ^ x[5];
  assign t[43] = t[67] ^ x[11];
  assign t[44] = t[68] ^ x[8];
  assign t[45] = t[69] ^ x[9];
  assign t[46] = t[70] ^ x[10];
  assign t[47] = t[71] ^ x[16];
  assign t[48] = t[72] ^ x[13];
  assign t[49] = t[73] ^ x[14];
  assign t[4] = ~t[5];
  assign t[50] = t[74] ^ x[15];
  assign t[51] = t[75] ^ x[21];
  assign t[52] = t[76] ^ x[18];
  assign t[53] = t[77] ^ x[19];
  assign t[54] = t[78] ^ x[20];
  assign t[55] = t[79] ^ x[26];
  assign t[56] = t[80] ^ x[23];
  assign t[57] = t[81] ^ x[24];
  assign t[58] = t[82] ^ x[25];
  assign t[59] = t[83] ^ x[31];
  assign t[5] = t[6] ^ t[7];
  assign t[60] = t[84] ^ x[28];
  assign t[61] = t[85] ^ x[29];
  assign t[62] = t[86] ^ x[30];
  assign t[63] = (x[2]);
  assign t[64] = (x[2]);
  assign t[65] = (x[2]);
  assign t[66] = (x[2]);
  assign t[67] = (x[7]);
  assign t[68] = (x[7]);
  assign t[69] = (x[7]);
  assign t[6] = t[8] ^ t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[12]);
  assign t[72] = (x[12]);
  assign t[73] = (x[12]);
  assign t[74] = (x[12]);
  assign t[75] = (x[17]);
  assign t[76] = (x[17]);
  assign t[77] = (x[17]);
  assign t[78] = (x[17]);
  assign t[79] = (x[22]);
  assign t[7] = t[10] & t[11];
  assign t[80] = (x[22]);
  assign t[81] = (x[22]);
  assign t[82] = (x[22]);
  assign t[83] = (x[27]);
  assign t[84] = (x[27]);
  assign t[85] = (x[27]);
  assign t[86] = (x[27]);
  assign t[8] = t[23] & t[12];
  assign t[9] = t[13] & t[14];
  assign y = (t[0]);
endmodule

module R2ind210(x, y);
 input [31:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[13];
  assign t[11] = t[16] ^ t[9];
  assign t[12] = t[17] ^ t[18];
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[23] ^ t[13]);
  assign t[15] = t[25] ^ t[24];
  assign t[16] = ~(t[19] ^ t[10]);
  assign t[17] = t[23] ^ t[15];
  assign t[18] = t[13] & t[19];
  assign t[19] = t[23] ^ t[20];
  assign t[1] = ~(t[2] ^ t[21]);
  assign t[20] = t[24] ^ t[26];
  assign t[21] = (t[27]);
  assign t[22] = (t[28]);
  assign t[23] = (t[29]);
  assign t[24] = (t[30]);
  assign t[25] = (t[31]);
  assign t[26] = (t[32]);
  assign t[27] = t[33] ^ x[6];
  assign t[28] = t[34] ^ x[11];
  assign t[29] = t[35] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[36] ^ x[21];
  assign t[31] = t[37] ^ x[26];
  assign t[32] = t[38] ^ x[31];
  assign t[33] = (~t[39] & t[40] & t[41] & t[42]) | (t[39] & ~t[41] & ~t[42]) | (t[39] & ~t[40] & ~t[42]) | (t[39] & ~t[40] & ~t[41]);
  assign t[34] = (~t[43] & t[44] & t[45] & t[46]) | (t[43] & ~t[45] & ~t[46]) | (t[43] & ~t[44] & ~t[46]) | (t[43] & ~t[44] & ~t[45]);
  assign t[35] = (~t[47] & t[48] & t[49] & t[50]) | (t[47] & ~t[49] & ~t[50]) | (t[47] & ~t[48] & ~t[50]) | (t[47] & ~t[48] & ~t[49]);
  assign t[36] = (~t[51] & t[52] & t[53] & t[54]) | (t[51] & ~t[53] & ~t[54]) | (t[51] & ~t[52] & ~t[54]) | (t[51] & ~t[52] & ~t[53]);
  assign t[37] = (~t[55] & t[56] & t[57] & t[58]) | (t[55] & ~t[57] & ~t[58]) | (t[55] & ~t[56] & ~t[58]) | (t[55] & ~t[56] & ~t[57]);
  assign t[38] = (~t[59] & t[60] & t[61] & t[62]) | (t[59] & ~t[61] & ~t[62]) | (t[59] & ~t[60] & ~t[62]) | (t[59] & ~t[60] & ~t[61]);
  assign t[39] = t[63] ^ x[6];
  assign t[3] = ~(t[4] ^ t[22]);
  assign t[40] = t[64] ^ x[3];
  assign t[41] = t[65] ^ x[4];
  assign t[42] = t[66] ^ x[5];
  assign t[43] = t[67] ^ x[11];
  assign t[44] = t[68] ^ x[8];
  assign t[45] = t[69] ^ x[9];
  assign t[46] = t[70] ^ x[10];
  assign t[47] = t[71] ^ x[16];
  assign t[48] = t[72] ^ x[13];
  assign t[49] = t[73] ^ x[14];
  assign t[4] = ~t[5];
  assign t[50] = t[74] ^ x[15];
  assign t[51] = t[75] ^ x[21];
  assign t[52] = t[76] ^ x[18];
  assign t[53] = t[77] ^ x[19];
  assign t[54] = t[78] ^ x[20];
  assign t[55] = t[79] ^ x[26];
  assign t[56] = t[80] ^ x[23];
  assign t[57] = t[81] ^ x[24];
  assign t[58] = t[82] ^ x[25];
  assign t[59] = t[83] ^ x[31];
  assign t[5] = t[6] ^ t[7];
  assign t[60] = t[84] ^ x[28];
  assign t[61] = t[85] ^ x[29];
  assign t[62] = t[86] ^ x[30];
  assign t[63] = (x[2]);
  assign t[64] = (x[2]);
  assign t[65] = (x[2]);
  assign t[66] = (x[2]);
  assign t[67] = (x[7]);
  assign t[68] = (x[7]);
  assign t[69] = (x[7]);
  assign t[6] = t[8] ^ t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[12]);
  assign t[72] = (x[12]);
  assign t[73] = (x[12]);
  assign t[74] = (x[12]);
  assign t[75] = (x[17]);
  assign t[76] = (x[17]);
  assign t[77] = (x[17]);
  assign t[78] = (x[17]);
  assign t[79] = (x[22]);
  assign t[7] = t[10] & t[11];
  assign t[80] = (x[22]);
  assign t[81] = (x[22]);
  assign t[82] = (x[22]);
  assign t[83] = (x[27]);
  assign t[84] = (x[27]);
  assign t[85] = (x[27]);
  assign t[86] = (x[27]);
  assign t[8] = t[23] & t[12];
  assign t[9] = t[13] & t[14];
  assign y = (t[0]);
endmodule

module R2ind211(x, y);
 input [31:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[13];
  assign t[11] = t[16] ^ t[9];
  assign t[12] = t[17] ^ t[18];
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[23] ^ t[13]);
  assign t[15] = t[25] ^ t[24];
  assign t[16] = ~(t[19] ^ t[10]);
  assign t[17] = t[23] ^ t[15];
  assign t[18] = t[13] & t[19];
  assign t[19] = t[23] ^ t[20];
  assign t[1] = ~(t[2] ^ t[21]);
  assign t[20] = t[24] ^ t[26];
  assign t[21] = (t[27]);
  assign t[22] = (t[28]);
  assign t[23] = (t[29]);
  assign t[24] = (t[30]);
  assign t[25] = (t[31]);
  assign t[26] = (t[32]);
  assign t[27] = t[33] ^ x[6];
  assign t[28] = t[34] ^ x[11];
  assign t[29] = t[35] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[36] ^ x[21];
  assign t[31] = t[37] ^ x[26];
  assign t[32] = t[38] ^ x[31];
  assign t[33] = (~t[39] & t[40] & t[41] & t[42]) | (t[39] & ~t[41] & ~t[42]) | (t[39] & ~t[40] & ~t[42]) | (t[39] & ~t[40] & ~t[41]);
  assign t[34] = (~t[43] & t[44] & t[45] & t[46]) | (t[43] & ~t[45] & ~t[46]) | (t[43] & ~t[44] & ~t[46]) | (t[43] & ~t[44] & ~t[45]);
  assign t[35] = (~t[47] & t[48] & t[49] & t[50]) | (t[47] & ~t[49] & ~t[50]) | (t[47] & ~t[48] & ~t[50]) | (t[47] & ~t[48] & ~t[49]);
  assign t[36] = (~t[51] & t[52] & t[53] & t[54]) | (t[51] & ~t[53] & ~t[54]) | (t[51] & ~t[52] & ~t[54]) | (t[51] & ~t[52] & ~t[53]);
  assign t[37] = (~t[55] & t[56] & t[57] & t[58]) | (t[55] & ~t[57] & ~t[58]) | (t[55] & ~t[56] & ~t[58]) | (t[55] & ~t[56] & ~t[57]);
  assign t[38] = (~t[59] & t[60] & t[61] & t[62]) | (t[59] & ~t[61] & ~t[62]) | (t[59] & ~t[60] & ~t[62]) | (t[59] & ~t[60] & ~t[61]);
  assign t[39] = t[63] ^ x[6];
  assign t[3] = ~(t[4] ^ t[22]);
  assign t[40] = t[64] ^ x[3];
  assign t[41] = t[65] ^ x[4];
  assign t[42] = t[66] ^ x[5];
  assign t[43] = t[67] ^ x[11];
  assign t[44] = t[68] ^ x[8];
  assign t[45] = t[69] ^ x[9];
  assign t[46] = t[70] ^ x[10];
  assign t[47] = t[71] ^ x[16];
  assign t[48] = t[72] ^ x[13];
  assign t[49] = t[73] ^ x[14];
  assign t[4] = ~t[5];
  assign t[50] = t[74] ^ x[15];
  assign t[51] = t[75] ^ x[21];
  assign t[52] = t[76] ^ x[18];
  assign t[53] = t[77] ^ x[19];
  assign t[54] = t[78] ^ x[20];
  assign t[55] = t[79] ^ x[26];
  assign t[56] = t[80] ^ x[23];
  assign t[57] = t[81] ^ x[24];
  assign t[58] = t[82] ^ x[25];
  assign t[59] = t[83] ^ x[31];
  assign t[5] = t[6] ^ t[7];
  assign t[60] = t[84] ^ x[28];
  assign t[61] = t[85] ^ x[29];
  assign t[62] = t[86] ^ x[30];
  assign t[63] = (x[2]);
  assign t[64] = (x[2]);
  assign t[65] = (x[2]);
  assign t[66] = (x[2]);
  assign t[67] = (x[7]);
  assign t[68] = (x[7]);
  assign t[69] = (x[7]);
  assign t[6] = t[8] ^ t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[12]);
  assign t[72] = (x[12]);
  assign t[73] = (x[12]);
  assign t[74] = (x[12]);
  assign t[75] = (x[17]);
  assign t[76] = (x[17]);
  assign t[77] = (x[17]);
  assign t[78] = (x[17]);
  assign t[79] = (x[22]);
  assign t[7] = t[10] & t[11];
  assign t[80] = (x[22]);
  assign t[81] = (x[22]);
  assign t[82] = (x[22]);
  assign t[83] = (x[27]);
  assign t[84] = (x[27]);
  assign t[85] = (x[27]);
  assign t[86] = (x[27]);
  assign t[8] = t[23] & t[12];
  assign t[9] = t[13] & t[14];
  assign y = (t[0]);
endmodule

module R2ind212(x, y);
 input [31:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[16] ^ t[9];
  assign t[11] = t[23] ^ t[14];
  assign t[12] = t[24] ^ t[25];
  assign t[13] = t[14] & t[17];
  assign t[14] = ~(t[25]);
  assign t[15] = ~(t[23] ^ t[14]);
  assign t[16] = t[23] & t[18];
  assign t[17] = t[23] ^ t[19];
  assign t[18] = t[20] ^ t[13];
  assign t[19] = t[25] ^ t[26];
  assign t[1] = ~(t[2] ^ t[21]);
  assign t[20] = t[23] ^ t[12];
  assign t[21] = (t[27]);
  assign t[22] = (t[28]);
  assign t[23] = (t[29]);
  assign t[24] = (t[30]);
  assign t[25] = (t[31]);
  assign t[26] = (t[32]);
  assign t[27] = t[33] ^ x[6];
  assign t[28] = t[34] ^ x[11];
  assign t[29] = t[35] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[36] ^ x[21];
  assign t[31] = t[37] ^ x[26];
  assign t[32] = t[38] ^ x[31];
  assign t[33] = (~t[39] & t[40] & t[41] & t[42]) | (t[39] & ~t[41] & ~t[42]) | (t[39] & ~t[40] & ~t[42]) | (t[39] & ~t[40] & ~t[41]);
  assign t[34] = (~t[43] & t[44] & t[45] & t[46]) | (t[43] & ~t[45] & ~t[46]) | (t[43] & ~t[44] & ~t[46]) | (t[43] & ~t[44] & ~t[45]);
  assign t[35] = (~t[47] & t[48] & t[49] & t[50]) | (t[47] & ~t[49] & ~t[50]) | (t[47] & ~t[48] & ~t[50]) | (t[47] & ~t[48] & ~t[49]);
  assign t[36] = (~t[51] & t[52] & t[53] & t[54]) | (t[51] & ~t[53] & ~t[54]) | (t[51] & ~t[52] & ~t[54]) | (t[51] & ~t[52] & ~t[53]);
  assign t[37] = (~t[55] & t[56] & t[57] & t[58]) | (t[55] & ~t[57] & ~t[58]) | (t[55] & ~t[56] & ~t[58]) | (t[55] & ~t[56] & ~t[57]);
  assign t[38] = (~t[59] & t[60] & t[61] & t[62]) | (t[59] & ~t[61] & ~t[62]) | (t[59] & ~t[60] & ~t[62]) | (t[59] & ~t[60] & ~t[61]);
  assign t[39] = t[63] ^ x[6];
  assign t[3] = ~(t[4] ^ t[22]);
  assign t[40] = t[64] ^ x[3];
  assign t[41] = t[65] ^ x[4];
  assign t[42] = t[66] ^ x[5];
  assign t[43] = t[67] ^ x[11];
  assign t[44] = t[68] ^ x[8];
  assign t[45] = t[69] ^ x[9];
  assign t[46] = t[70] ^ x[10];
  assign t[47] = t[71] ^ x[16];
  assign t[48] = t[72] ^ x[13];
  assign t[49] = t[73] ^ x[14];
  assign t[4] = ~t[5];
  assign t[50] = t[74] ^ x[15];
  assign t[51] = t[75] ^ x[21];
  assign t[52] = t[76] ^ x[18];
  assign t[53] = t[77] ^ x[19];
  assign t[54] = t[78] ^ x[20];
  assign t[55] = t[79] ^ x[26];
  assign t[56] = t[80] ^ x[23];
  assign t[57] = t[81] ^ x[24];
  assign t[58] = t[82] ^ x[25];
  assign t[59] = t[83] ^ x[31];
  assign t[5] = ~(t[6] ^ t[7]);
  assign t[60] = t[84] ^ x[28];
  assign t[61] = t[85] ^ x[29];
  assign t[62] = t[86] ^ x[30];
  assign t[63] = (x[2]);
  assign t[64] = (x[2]);
  assign t[65] = (x[2]);
  assign t[66] = (x[2]);
  assign t[67] = (x[7]);
  assign t[68] = (x[7]);
  assign t[69] = (x[7]);
  assign t[6] = t[8] ^ t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[12]);
  assign t[72] = (x[12]);
  assign t[73] = (x[12]);
  assign t[74] = (x[12]);
  assign t[75] = (x[17]);
  assign t[76] = (x[17]);
  assign t[77] = (x[17]);
  assign t[78] = (x[17]);
  assign t[79] = (x[22]);
  assign t[7] = t[10] ^ t[11];
  assign t[80] = (x[22]);
  assign t[81] = (x[22]);
  assign t[82] = (x[22]);
  assign t[83] = (x[27]);
  assign t[84] = (x[27]);
  assign t[85] = (x[27]);
  assign t[86] = (x[27]);
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind213(x, y);
 input [31:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[16] ^ t[9];
  assign t[11] = t[23] ^ t[14];
  assign t[12] = t[24] ^ t[25];
  assign t[13] = t[14] & t[17];
  assign t[14] = ~(t[25]);
  assign t[15] = ~(t[23] ^ t[14]);
  assign t[16] = t[23] & t[18];
  assign t[17] = t[23] ^ t[19];
  assign t[18] = t[20] ^ t[13];
  assign t[19] = t[25] ^ t[26];
  assign t[1] = ~(t[2] ^ t[21]);
  assign t[20] = t[23] ^ t[12];
  assign t[21] = (t[27]);
  assign t[22] = (t[28]);
  assign t[23] = (t[29]);
  assign t[24] = (t[30]);
  assign t[25] = (t[31]);
  assign t[26] = (t[32]);
  assign t[27] = t[33] ^ x[6];
  assign t[28] = t[34] ^ x[11];
  assign t[29] = t[35] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[36] ^ x[21];
  assign t[31] = t[37] ^ x[26];
  assign t[32] = t[38] ^ x[31];
  assign t[33] = (~t[39] & t[40] & t[41] & t[42]) | (t[39] & ~t[41] & ~t[42]) | (t[39] & ~t[40] & ~t[42]) | (t[39] & ~t[40] & ~t[41]);
  assign t[34] = (~t[43] & t[44] & t[45] & t[46]) | (t[43] & ~t[45] & ~t[46]) | (t[43] & ~t[44] & ~t[46]) | (t[43] & ~t[44] & ~t[45]);
  assign t[35] = (~t[47] & t[48] & t[49] & t[50]) | (t[47] & ~t[49] & ~t[50]) | (t[47] & ~t[48] & ~t[50]) | (t[47] & ~t[48] & ~t[49]);
  assign t[36] = (~t[51] & t[52] & t[53] & t[54]) | (t[51] & ~t[53] & ~t[54]) | (t[51] & ~t[52] & ~t[54]) | (t[51] & ~t[52] & ~t[53]);
  assign t[37] = (~t[55] & t[56] & t[57] & t[58]) | (t[55] & ~t[57] & ~t[58]) | (t[55] & ~t[56] & ~t[58]) | (t[55] & ~t[56] & ~t[57]);
  assign t[38] = (~t[59] & t[60] & t[61] & t[62]) | (t[59] & ~t[61] & ~t[62]) | (t[59] & ~t[60] & ~t[62]) | (t[59] & ~t[60] & ~t[61]);
  assign t[39] = t[63] ^ x[6];
  assign t[3] = ~(t[4] ^ t[22]);
  assign t[40] = t[64] ^ x[3];
  assign t[41] = t[65] ^ x[4];
  assign t[42] = t[66] ^ x[5];
  assign t[43] = t[67] ^ x[11];
  assign t[44] = t[68] ^ x[8];
  assign t[45] = t[69] ^ x[9];
  assign t[46] = t[70] ^ x[10];
  assign t[47] = t[71] ^ x[16];
  assign t[48] = t[72] ^ x[13];
  assign t[49] = t[73] ^ x[14];
  assign t[4] = ~t[5];
  assign t[50] = t[74] ^ x[15];
  assign t[51] = t[75] ^ x[21];
  assign t[52] = t[76] ^ x[18];
  assign t[53] = t[77] ^ x[19];
  assign t[54] = t[78] ^ x[20];
  assign t[55] = t[79] ^ x[26];
  assign t[56] = t[80] ^ x[23];
  assign t[57] = t[81] ^ x[24];
  assign t[58] = t[82] ^ x[25];
  assign t[59] = t[83] ^ x[31];
  assign t[5] = ~(t[6] ^ t[7]);
  assign t[60] = t[84] ^ x[28];
  assign t[61] = t[85] ^ x[29];
  assign t[62] = t[86] ^ x[30];
  assign t[63] = (x[2]);
  assign t[64] = (x[2]);
  assign t[65] = (x[2]);
  assign t[66] = (x[2]);
  assign t[67] = (x[7]);
  assign t[68] = (x[7]);
  assign t[69] = (x[7]);
  assign t[6] = t[8] ^ t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[12]);
  assign t[72] = (x[12]);
  assign t[73] = (x[12]);
  assign t[74] = (x[12]);
  assign t[75] = (x[17]);
  assign t[76] = (x[17]);
  assign t[77] = (x[17]);
  assign t[78] = (x[17]);
  assign t[79] = (x[22]);
  assign t[7] = t[10] ^ t[11];
  assign t[80] = (x[22]);
  assign t[81] = (x[22]);
  assign t[82] = (x[22]);
  assign t[83] = (x[27]);
  assign t[84] = (x[27]);
  assign t[85] = (x[27]);
  assign t[86] = (x[27]);
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind214(x, y);
 input [31:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[16] ^ t[9];
  assign t[11] = t[23] ^ t[14];
  assign t[12] = t[24] ^ t[25];
  assign t[13] = t[14] & t[17];
  assign t[14] = ~(t[25]);
  assign t[15] = ~(t[23] ^ t[14]);
  assign t[16] = t[23] & t[18];
  assign t[17] = t[23] ^ t[19];
  assign t[18] = t[20] ^ t[13];
  assign t[19] = t[25] ^ t[26];
  assign t[1] = ~(t[2] ^ t[21]);
  assign t[20] = t[23] ^ t[12];
  assign t[21] = (t[27]);
  assign t[22] = (t[28]);
  assign t[23] = (t[29]);
  assign t[24] = (t[30]);
  assign t[25] = (t[31]);
  assign t[26] = (t[32]);
  assign t[27] = t[33] ^ x[6];
  assign t[28] = t[34] ^ x[11];
  assign t[29] = t[35] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[36] ^ x[21];
  assign t[31] = t[37] ^ x[26];
  assign t[32] = t[38] ^ x[31];
  assign t[33] = (~t[39] & t[40] & t[41] & t[42]) | (t[39] & ~t[41] & ~t[42]) | (t[39] & ~t[40] & ~t[42]) | (t[39] & ~t[40] & ~t[41]);
  assign t[34] = (~t[43] & t[44] & t[45] & t[46]) | (t[43] & ~t[45] & ~t[46]) | (t[43] & ~t[44] & ~t[46]) | (t[43] & ~t[44] & ~t[45]);
  assign t[35] = (~t[47] & t[48] & t[49] & t[50]) | (t[47] & ~t[49] & ~t[50]) | (t[47] & ~t[48] & ~t[50]) | (t[47] & ~t[48] & ~t[49]);
  assign t[36] = (~t[51] & t[52] & t[53] & t[54]) | (t[51] & ~t[53] & ~t[54]) | (t[51] & ~t[52] & ~t[54]) | (t[51] & ~t[52] & ~t[53]);
  assign t[37] = (~t[55] & t[56] & t[57] & t[58]) | (t[55] & ~t[57] & ~t[58]) | (t[55] & ~t[56] & ~t[58]) | (t[55] & ~t[56] & ~t[57]);
  assign t[38] = (~t[59] & t[60] & t[61] & t[62]) | (t[59] & ~t[61] & ~t[62]) | (t[59] & ~t[60] & ~t[62]) | (t[59] & ~t[60] & ~t[61]);
  assign t[39] = t[63] ^ x[6];
  assign t[3] = ~(t[4] ^ t[22]);
  assign t[40] = t[64] ^ x[3];
  assign t[41] = t[65] ^ x[4];
  assign t[42] = t[66] ^ x[5];
  assign t[43] = t[67] ^ x[11];
  assign t[44] = t[68] ^ x[8];
  assign t[45] = t[69] ^ x[9];
  assign t[46] = t[70] ^ x[10];
  assign t[47] = t[71] ^ x[16];
  assign t[48] = t[72] ^ x[13];
  assign t[49] = t[73] ^ x[14];
  assign t[4] = ~t[5];
  assign t[50] = t[74] ^ x[15];
  assign t[51] = t[75] ^ x[21];
  assign t[52] = t[76] ^ x[18];
  assign t[53] = t[77] ^ x[19];
  assign t[54] = t[78] ^ x[20];
  assign t[55] = t[79] ^ x[26];
  assign t[56] = t[80] ^ x[23];
  assign t[57] = t[81] ^ x[24];
  assign t[58] = t[82] ^ x[25];
  assign t[59] = t[83] ^ x[31];
  assign t[5] = ~(t[6] ^ t[7]);
  assign t[60] = t[84] ^ x[28];
  assign t[61] = t[85] ^ x[29];
  assign t[62] = t[86] ^ x[30];
  assign t[63] = (x[2]);
  assign t[64] = (x[2]);
  assign t[65] = (x[2]);
  assign t[66] = (x[2]);
  assign t[67] = (x[7]);
  assign t[68] = (x[7]);
  assign t[69] = (x[7]);
  assign t[6] = t[8] ^ t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[12]);
  assign t[72] = (x[12]);
  assign t[73] = (x[12]);
  assign t[74] = (x[12]);
  assign t[75] = (x[17]);
  assign t[76] = (x[17]);
  assign t[77] = (x[17]);
  assign t[78] = (x[17]);
  assign t[79] = (x[22]);
  assign t[7] = t[10] ^ t[11];
  assign t[80] = (x[22]);
  assign t[81] = (x[22]);
  assign t[82] = (x[22]);
  assign t[83] = (x[27]);
  assign t[84] = (x[27]);
  assign t[85] = (x[27]);
  assign t[86] = (x[27]);
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind215(x, y);
 input [31:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[16] ^ t[9];
  assign t[11] = t[23] ^ t[14];
  assign t[12] = t[24] ^ t[25];
  assign t[13] = t[14] & t[17];
  assign t[14] = ~(t[25]);
  assign t[15] = ~(t[23] ^ t[14]);
  assign t[16] = t[23] & t[18];
  assign t[17] = t[23] ^ t[19];
  assign t[18] = t[20] ^ t[13];
  assign t[19] = t[25] ^ t[26];
  assign t[1] = ~(t[2] ^ t[21]);
  assign t[20] = t[23] ^ t[12];
  assign t[21] = (t[27]);
  assign t[22] = (t[28]);
  assign t[23] = (t[29]);
  assign t[24] = (t[30]);
  assign t[25] = (t[31]);
  assign t[26] = (t[32]);
  assign t[27] = t[33] ^ x[6];
  assign t[28] = t[34] ^ x[11];
  assign t[29] = t[35] ^ x[16];
  assign t[2] = ~t[3];
  assign t[30] = t[36] ^ x[21];
  assign t[31] = t[37] ^ x[26];
  assign t[32] = t[38] ^ x[31];
  assign t[33] = (~t[39] & t[40] & t[41] & t[42]) | (t[39] & ~t[41] & ~t[42]) | (t[39] & ~t[40] & ~t[42]) | (t[39] & ~t[40] & ~t[41]);
  assign t[34] = (~t[43] & t[44] & t[45] & t[46]) | (t[43] & ~t[45] & ~t[46]) | (t[43] & ~t[44] & ~t[46]) | (t[43] & ~t[44] & ~t[45]);
  assign t[35] = (~t[47] & t[48] & t[49] & t[50]) | (t[47] & ~t[49] & ~t[50]) | (t[47] & ~t[48] & ~t[50]) | (t[47] & ~t[48] & ~t[49]);
  assign t[36] = (~t[51] & t[52] & t[53] & t[54]) | (t[51] & ~t[53] & ~t[54]) | (t[51] & ~t[52] & ~t[54]) | (t[51] & ~t[52] & ~t[53]);
  assign t[37] = (~t[55] & t[56] & t[57] & t[58]) | (t[55] & ~t[57] & ~t[58]) | (t[55] & ~t[56] & ~t[58]) | (t[55] & ~t[56] & ~t[57]);
  assign t[38] = (~t[59] & t[60] & t[61] & t[62]) | (t[59] & ~t[61] & ~t[62]) | (t[59] & ~t[60] & ~t[62]) | (t[59] & ~t[60] & ~t[61]);
  assign t[39] = t[63] ^ x[6];
  assign t[3] = ~(t[4] ^ t[22]);
  assign t[40] = t[64] ^ x[3];
  assign t[41] = t[65] ^ x[4];
  assign t[42] = t[66] ^ x[5];
  assign t[43] = t[67] ^ x[11];
  assign t[44] = t[68] ^ x[8];
  assign t[45] = t[69] ^ x[9];
  assign t[46] = t[70] ^ x[10];
  assign t[47] = t[71] ^ x[16];
  assign t[48] = t[72] ^ x[13];
  assign t[49] = t[73] ^ x[14];
  assign t[4] = ~t[5];
  assign t[50] = t[74] ^ x[15];
  assign t[51] = t[75] ^ x[21];
  assign t[52] = t[76] ^ x[18];
  assign t[53] = t[77] ^ x[19];
  assign t[54] = t[78] ^ x[20];
  assign t[55] = t[79] ^ x[26];
  assign t[56] = t[80] ^ x[23];
  assign t[57] = t[81] ^ x[24];
  assign t[58] = t[82] ^ x[25];
  assign t[59] = t[83] ^ x[31];
  assign t[5] = ~(t[6] ^ t[7]);
  assign t[60] = t[84] ^ x[28];
  assign t[61] = t[85] ^ x[29];
  assign t[62] = t[86] ^ x[30];
  assign t[63] = (x[2]);
  assign t[64] = (x[2]);
  assign t[65] = (x[2]);
  assign t[66] = (x[2]);
  assign t[67] = (x[7]);
  assign t[68] = (x[7]);
  assign t[69] = (x[7]);
  assign t[6] = t[8] ^ t[9];
  assign t[70] = (x[7]);
  assign t[71] = (x[12]);
  assign t[72] = (x[12]);
  assign t[73] = (x[12]);
  assign t[74] = (x[12]);
  assign t[75] = (x[17]);
  assign t[76] = (x[17]);
  assign t[77] = (x[17]);
  assign t[78] = (x[17]);
  assign t[79] = (x[22]);
  assign t[7] = t[10] ^ t[11];
  assign t[80] = (x[22]);
  assign t[81] = (x[22]);
  assign t[82] = (x[22]);
  assign t[83] = (x[27]);
  assign t[84] = (x[27]);
  assign t[85] = (x[27]);
  assign t[86] = (x[27]);
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] & t[15];
  assign y = (t[0]);
endmodule

module R2ind216(x, y);
 input [26:0] x;
 output y;

 wire [65:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[15] ^ t[9]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[6];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[16];
  assign t[19] = t[24] ^ x[21];
  assign t[1] = ~(t[2] ^ t[11]);
  assign t[20] = t[25] ^ x[26];
  assign t[21] = (~t[26] & t[27] & t[28] & t[29]) | (t[26] & ~t[28] & ~t[29]) | (t[26] & ~t[27] & ~t[29]) | (t[26] & ~t[27] & ~t[28]);
  assign t[22] = (~t[30] & t[31] & t[32] & t[33]) | (t[30] & ~t[32] & ~t[33]) | (t[30] & ~t[31] & ~t[33]) | (t[30] & ~t[31] & ~t[32]);
  assign t[23] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[24] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[25] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[26] = t[46] ^ x[6];
  assign t[27] = t[47] ^ x[3];
  assign t[28] = t[48] ^ x[4];
  assign t[29] = t[49] ^ x[5];
  assign t[2] = ~t[3];
  assign t[30] = t[50] ^ x[11];
  assign t[31] = t[51] ^ x[8];
  assign t[32] = t[52] ^ x[9];
  assign t[33] = t[53] ^ x[10];
  assign t[34] = t[54] ^ x[16];
  assign t[35] = t[55] ^ x[13];
  assign t[36] = t[56] ^ x[14];
  assign t[37] = t[57] ^ x[15];
  assign t[38] = t[58] ^ x[21];
  assign t[39] = t[59] ^ x[18];
  assign t[3] = ~(t[4] ^ t[12]);
  assign t[40] = t[60] ^ x[19];
  assign t[41] = t[61] ^ x[20];
  assign t[42] = t[62] ^ x[26];
  assign t[43] = t[63] ^ x[23];
  assign t[44] = t[64] ^ x[24];
  assign t[45] = t[65] ^ x[25];
  assign t[46] = (x[2]);
  assign t[47] = (x[2]);
  assign t[48] = (x[2]);
  assign t[49] = (x[2]);
  assign t[4] = ~t[5];
  assign t[50] = (x[7]);
  assign t[51] = (x[7]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[12]);
  assign t[55] = (x[12]);
  assign t[56] = (x[12]);
  assign t[57] = (x[12]);
  assign t[58] = (x[17]);
  assign t[59] = (x[17]);
  assign t[5] = ~(t[6]);
  assign t[60] = (x[17]);
  assign t[61] = (x[17]);
  assign t[62] = (x[22]);
  assign t[63] = (x[22]);
  assign t[64] = (x[22]);
  assign t[65] = (x[22]);
  assign t[6] = t[7] ^ t[8];
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[9] & t[10];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind217(x, y);
 input [26:0] x;
 output y;

 wire [65:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[15] ^ t[9]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[6];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[16];
  assign t[19] = t[24] ^ x[21];
  assign t[1] = ~(t[2] ^ t[11]);
  assign t[20] = t[25] ^ x[26];
  assign t[21] = (~t[26] & t[27] & t[28] & t[29]) | (t[26] & ~t[28] & ~t[29]) | (t[26] & ~t[27] & ~t[29]) | (t[26] & ~t[27] & ~t[28]);
  assign t[22] = (~t[30] & t[31] & t[32] & t[33]) | (t[30] & ~t[32] & ~t[33]) | (t[30] & ~t[31] & ~t[33]) | (t[30] & ~t[31] & ~t[32]);
  assign t[23] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[24] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[25] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[26] = t[46] ^ x[6];
  assign t[27] = t[47] ^ x[3];
  assign t[28] = t[48] ^ x[4];
  assign t[29] = t[49] ^ x[5];
  assign t[2] = ~t[3];
  assign t[30] = t[50] ^ x[11];
  assign t[31] = t[51] ^ x[8];
  assign t[32] = t[52] ^ x[9];
  assign t[33] = t[53] ^ x[10];
  assign t[34] = t[54] ^ x[16];
  assign t[35] = t[55] ^ x[13];
  assign t[36] = t[56] ^ x[14];
  assign t[37] = t[57] ^ x[15];
  assign t[38] = t[58] ^ x[21];
  assign t[39] = t[59] ^ x[18];
  assign t[3] = ~(t[4] ^ t[12]);
  assign t[40] = t[60] ^ x[19];
  assign t[41] = t[61] ^ x[20];
  assign t[42] = t[62] ^ x[26];
  assign t[43] = t[63] ^ x[23];
  assign t[44] = t[64] ^ x[24];
  assign t[45] = t[65] ^ x[25];
  assign t[46] = (x[2]);
  assign t[47] = (x[2]);
  assign t[48] = (x[2]);
  assign t[49] = (x[2]);
  assign t[4] = ~t[5];
  assign t[50] = (x[7]);
  assign t[51] = (x[7]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[12]);
  assign t[55] = (x[12]);
  assign t[56] = (x[12]);
  assign t[57] = (x[12]);
  assign t[58] = (x[17]);
  assign t[59] = (x[17]);
  assign t[5] = ~(t[6]);
  assign t[60] = (x[17]);
  assign t[61] = (x[17]);
  assign t[62] = (x[22]);
  assign t[63] = (x[22]);
  assign t[64] = (x[22]);
  assign t[65] = (x[22]);
  assign t[6] = t[7] ^ t[8];
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[9] & t[10];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind218(x, y);
 input [26:0] x;
 output y;

 wire [65:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[15] ^ t[9]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[6];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[16];
  assign t[19] = t[24] ^ x[21];
  assign t[1] = ~(t[2] ^ t[11]);
  assign t[20] = t[25] ^ x[26];
  assign t[21] = (~t[26] & t[27] & t[28] & t[29]) | (t[26] & ~t[28] & ~t[29]) | (t[26] & ~t[27] & ~t[29]) | (t[26] & ~t[27] & ~t[28]);
  assign t[22] = (~t[30] & t[31] & t[32] & t[33]) | (t[30] & ~t[32] & ~t[33]) | (t[30] & ~t[31] & ~t[33]) | (t[30] & ~t[31] & ~t[32]);
  assign t[23] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[24] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[25] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[26] = t[46] ^ x[6];
  assign t[27] = t[47] ^ x[3];
  assign t[28] = t[48] ^ x[4];
  assign t[29] = t[49] ^ x[5];
  assign t[2] = ~t[3];
  assign t[30] = t[50] ^ x[11];
  assign t[31] = t[51] ^ x[8];
  assign t[32] = t[52] ^ x[9];
  assign t[33] = t[53] ^ x[10];
  assign t[34] = t[54] ^ x[16];
  assign t[35] = t[55] ^ x[13];
  assign t[36] = t[56] ^ x[14];
  assign t[37] = t[57] ^ x[15];
  assign t[38] = t[58] ^ x[21];
  assign t[39] = t[59] ^ x[18];
  assign t[3] = ~(t[4] ^ t[12]);
  assign t[40] = t[60] ^ x[19];
  assign t[41] = t[61] ^ x[20];
  assign t[42] = t[62] ^ x[26];
  assign t[43] = t[63] ^ x[23];
  assign t[44] = t[64] ^ x[24];
  assign t[45] = t[65] ^ x[25];
  assign t[46] = (x[2]);
  assign t[47] = (x[2]);
  assign t[48] = (x[2]);
  assign t[49] = (x[2]);
  assign t[4] = ~t[5];
  assign t[50] = (x[7]);
  assign t[51] = (x[7]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[12]);
  assign t[55] = (x[12]);
  assign t[56] = (x[12]);
  assign t[57] = (x[12]);
  assign t[58] = (x[17]);
  assign t[59] = (x[17]);
  assign t[5] = ~(t[6]);
  assign t[60] = (x[17]);
  assign t[61] = (x[17]);
  assign t[62] = (x[22]);
  assign t[63] = (x[22]);
  assign t[64] = (x[22]);
  assign t[65] = (x[22]);
  assign t[6] = t[7] ^ t[8];
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[9] & t[10];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind219(x, y);
 input [26:0] x;
 output y;

 wire [65:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[15] ^ t[9]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[6];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[16];
  assign t[19] = t[24] ^ x[21];
  assign t[1] = ~(t[2] ^ t[11]);
  assign t[20] = t[25] ^ x[26];
  assign t[21] = (~t[26] & t[27] & t[28] & t[29]) | (t[26] & ~t[28] & ~t[29]) | (t[26] & ~t[27] & ~t[29]) | (t[26] & ~t[27] & ~t[28]);
  assign t[22] = (~t[30] & t[31] & t[32] & t[33]) | (t[30] & ~t[32] & ~t[33]) | (t[30] & ~t[31] & ~t[33]) | (t[30] & ~t[31] & ~t[32]);
  assign t[23] = (~t[34] & t[35] & t[36] & t[37]) | (t[34] & ~t[36] & ~t[37]) | (t[34] & ~t[35] & ~t[37]) | (t[34] & ~t[35] & ~t[36]);
  assign t[24] = (~t[38] & t[39] & t[40] & t[41]) | (t[38] & ~t[40] & ~t[41]) | (t[38] & ~t[39] & ~t[41]) | (t[38] & ~t[39] & ~t[40]);
  assign t[25] = (~t[42] & t[43] & t[44] & t[45]) | (t[42] & ~t[44] & ~t[45]) | (t[42] & ~t[43] & ~t[45]) | (t[42] & ~t[43] & ~t[44]);
  assign t[26] = t[46] ^ x[6];
  assign t[27] = t[47] ^ x[3];
  assign t[28] = t[48] ^ x[4];
  assign t[29] = t[49] ^ x[5];
  assign t[2] = ~t[3];
  assign t[30] = t[50] ^ x[11];
  assign t[31] = t[51] ^ x[8];
  assign t[32] = t[52] ^ x[9];
  assign t[33] = t[53] ^ x[10];
  assign t[34] = t[54] ^ x[16];
  assign t[35] = t[55] ^ x[13];
  assign t[36] = t[56] ^ x[14];
  assign t[37] = t[57] ^ x[15];
  assign t[38] = t[58] ^ x[21];
  assign t[39] = t[59] ^ x[18];
  assign t[3] = ~(t[4] ^ t[12]);
  assign t[40] = t[60] ^ x[19];
  assign t[41] = t[61] ^ x[20];
  assign t[42] = t[62] ^ x[26];
  assign t[43] = t[63] ^ x[23];
  assign t[44] = t[64] ^ x[24];
  assign t[45] = t[65] ^ x[25];
  assign t[46] = (x[2]);
  assign t[47] = (x[2]);
  assign t[48] = (x[2]);
  assign t[49] = (x[2]);
  assign t[4] = ~t[5];
  assign t[50] = (x[7]);
  assign t[51] = (x[7]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[12]);
  assign t[55] = (x[12]);
  assign t[56] = (x[12]);
  assign t[57] = (x[12]);
  assign t[58] = (x[17]);
  assign t[59] = (x[17]);
  assign t[5] = ~(t[6]);
  assign t[60] = (x[17]);
  assign t[61] = (x[17]);
  assign t[62] = (x[22]);
  assign t[63] = (x[22]);
  assign t[64] = (x[22]);
  assign t[65] = (x[22]);
  assign t[6] = t[7] ^ t[8];
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[9] & t[10];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind220(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[11] & t[13];
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] ^ t[14];
  assign t[14] = t[18] ^ t[20];
  assign t[15] = (t[21]);
  assign t[16] = (t[22]);
  assign t[17] = (t[23]);
  assign t[18] = (t[24]);
  assign t[19] = (t[25]);
  assign t[1] = ~(t[2] ^ t[15]);
  assign t[20] = (t[26]);
  assign t[21] = t[27] ^ x[6];
  assign t[22] = t[28] ^ x[11];
  assign t[23] = t[29] ^ x[16];
  assign t[24] = t[30] ^ x[21];
  assign t[25] = t[31] ^ x[26];
  assign t[26] = t[32] ^ x[31];
  assign t[27] = (~t[33] & t[34] & t[35] & t[36]) | (t[33] & ~t[35] & ~t[36]) | (t[33] & ~t[34] & ~t[36]) | (t[33] & ~t[34] & ~t[35]);
  assign t[28] = (~t[37] & t[38] & t[39] & t[40]) | (t[37] & ~t[39] & ~t[40]) | (t[37] & ~t[38] & ~t[40]) | (t[37] & ~t[38] & ~t[39]);
  assign t[29] = (~t[41] & t[42] & t[43] & t[44]) | (t[41] & ~t[43] & ~t[44]) | (t[41] & ~t[42] & ~t[44]) | (t[41] & ~t[42] & ~t[43]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[45] & t[46] & t[47] & t[48]) | (t[45] & ~t[47] & ~t[48]) | (t[45] & ~t[46] & ~t[48]) | (t[45] & ~t[46] & ~t[47]);
  assign t[31] = (~t[49] & t[50] & t[51] & t[52]) | (t[49] & ~t[51] & ~t[52]) | (t[49] & ~t[50] & ~t[52]) | (t[49] & ~t[50] & ~t[51]);
  assign t[32] = (~t[53] & t[54] & t[55] & t[56]) | (t[53] & ~t[55] & ~t[56]) | (t[53] & ~t[54] & ~t[56]) | (t[53] & ~t[54] & ~t[55]);
  assign t[33] = t[57] ^ x[6];
  assign t[34] = t[58] ^ x[3];
  assign t[35] = t[59] ^ x[4];
  assign t[36] = t[60] ^ x[5];
  assign t[37] = t[61] ^ x[11];
  assign t[38] = t[62] ^ x[8];
  assign t[39] = t[63] ^ x[9];
  assign t[3] = ~(t[4] ^ t[16]);
  assign t[40] = t[64] ^ x[10];
  assign t[41] = t[65] ^ x[16];
  assign t[42] = t[66] ^ x[13];
  assign t[43] = t[67] ^ x[14];
  assign t[44] = t[68] ^ x[15];
  assign t[45] = t[69] ^ x[21];
  assign t[46] = t[70] ^ x[18];
  assign t[47] = t[71] ^ x[19];
  assign t[48] = t[72] ^ x[20];
  assign t[49] = t[73] ^ x[26];
  assign t[4] = ~t[5];
  assign t[50] = t[74] ^ x[23];
  assign t[51] = t[75] ^ x[24];
  assign t[52] = t[76] ^ x[25];
  assign t[53] = t[77] ^ x[31];
  assign t[54] = t[78] ^ x[28];
  assign t[55] = t[79] ^ x[29];
  assign t[56] = t[80] ^ x[30];
  assign t[57] = (x[2]);
  assign t[58] = (x[2]);
  assign t[59] = (x[2]);
  assign t[5] = ~(t[6]);
  assign t[60] = (x[2]);
  assign t[61] = (x[7]);
  assign t[62] = (x[7]);
  assign t[63] = (x[7]);
  assign t[64] = (x[7]);
  assign t[65] = (x[12]);
  assign t[66] = (x[12]);
  assign t[67] = (x[12]);
  assign t[68] = (x[12]);
  assign t[69] = (x[17]);
  assign t[6] = t[7] ^ t[8];
  assign t[70] = (x[17]);
  assign t[71] = (x[17]);
  assign t[72] = (x[17]);
  assign t[73] = (x[22]);
  assign t[74] = (x[22]);
  assign t[75] = (x[22]);
  assign t[76] = (x[22]);
  assign t[77] = (x[27]);
  assign t[78] = (x[27]);
  assign t[79] = (x[27]);
  assign t[7] = t[9] ^ t[10];
  assign t[80] = (x[27]);
  assign t[8] = t[11] & t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = (t[0]);
endmodule

module R2ind221(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[11] & t[13];
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] ^ t[14];
  assign t[14] = t[18] ^ t[20];
  assign t[15] = (t[21]);
  assign t[16] = (t[22]);
  assign t[17] = (t[23]);
  assign t[18] = (t[24]);
  assign t[19] = (t[25]);
  assign t[1] = ~(t[2] ^ t[15]);
  assign t[20] = (t[26]);
  assign t[21] = t[27] ^ x[6];
  assign t[22] = t[28] ^ x[11];
  assign t[23] = t[29] ^ x[16];
  assign t[24] = t[30] ^ x[21];
  assign t[25] = t[31] ^ x[26];
  assign t[26] = t[32] ^ x[31];
  assign t[27] = (~t[33] & t[34] & t[35] & t[36]) | (t[33] & ~t[35] & ~t[36]) | (t[33] & ~t[34] & ~t[36]) | (t[33] & ~t[34] & ~t[35]);
  assign t[28] = (~t[37] & t[38] & t[39] & t[40]) | (t[37] & ~t[39] & ~t[40]) | (t[37] & ~t[38] & ~t[40]) | (t[37] & ~t[38] & ~t[39]);
  assign t[29] = (~t[41] & t[42] & t[43] & t[44]) | (t[41] & ~t[43] & ~t[44]) | (t[41] & ~t[42] & ~t[44]) | (t[41] & ~t[42] & ~t[43]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[45] & t[46] & t[47] & t[48]) | (t[45] & ~t[47] & ~t[48]) | (t[45] & ~t[46] & ~t[48]) | (t[45] & ~t[46] & ~t[47]);
  assign t[31] = (~t[49] & t[50] & t[51] & t[52]) | (t[49] & ~t[51] & ~t[52]) | (t[49] & ~t[50] & ~t[52]) | (t[49] & ~t[50] & ~t[51]);
  assign t[32] = (~t[53] & t[54] & t[55] & t[56]) | (t[53] & ~t[55] & ~t[56]) | (t[53] & ~t[54] & ~t[56]) | (t[53] & ~t[54] & ~t[55]);
  assign t[33] = t[57] ^ x[6];
  assign t[34] = t[58] ^ x[3];
  assign t[35] = t[59] ^ x[4];
  assign t[36] = t[60] ^ x[5];
  assign t[37] = t[61] ^ x[11];
  assign t[38] = t[62] ^ x[8];
  assign t[39] = t[63] ^ x[9];
  assign t[3] = ~(t[4] ^ t[16]);
  assign t[40] = t[64] ^ x[10];
  assign t[41] = t[65] ^ x[16];
  assign t[42] = t[66] ^ x[13];
  assign t[43] = t[67] ^ x[14];
  assign t[44] = t[68] ^ x[15];
  assign t[45] = t[69] ^ x[21];
  assign t[46] = t[70] ^ x[18];
  assign t[47] = t[71] ^ x[19];
  assign t[48] = t[72] ^ x[20];
  assign t[49] = t[73] ^ x[26];
  assign t[4] = ~t[5];
  assign t[50] = t[74] ^ x[23];
  assign t[51] = t[75] ^ x[24];
  assign t[52] = t[76] ^ x[25];
  assign t[53] = t[77] ^ x[31];
  assign t[54] = t[78] ^ x[28];
  assign t[55] = t[79] ^ x[29];
  assign t[56] = t[80] ^ x[30];
  assign t[57] = (x[2]);
  assign t[58] = (x[2]);
  assign t[59] = (x[2]);
  assign t[5] = ~(t[6]);
  assign t[60] = (x[2]);
  assign t[61] = (x[7]);
  assign t[62] = (x[7]);
  assign t[63] = (x[7]);
  assign t[64] = (x[7]);
  assign t[65] = (x[12]);
  assign t[66] = (x[12]);
  assign t[67] = (x[12]);
  assign t[68] = (x[12]);
  assign t[69] = (x[17]);
  assign t[6] = t[7] ^ t[8];
  assign t[70] = (x[17]);
  assign t[71] = (x[17]);
  assign t[72] = (x[17]);
  assign t[73] = (x[22]);
  assign t[74] = (x[22]);
  assign t[75] = (x[22]);
  assign t[76] = (x[22]);
  assign t[77] = (x[27]);
  assign t[78] = (x[27]);
  assign t[79] = (x[27]);
  assign t[7] = t[9] ^ t[10];
  assign t[80] = (x[27]);
  assign t[8] = t[11] & t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = (t[0]);
endmodule

module R2ind222(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[11] & t[13];
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] ^ t[14];
  assign t[14] = t[18] ^ t[20];
  assign t[15] = (t[21]);
  assign t[16] = (t[22]);
  assign t[17] = (t[23]);
  assign t[18] = (t[24]);
  assign t[19] = (t[25]);
  assign t[1] = ~(t[2] ^ t[15]);
  assign t[20] = (t[26]);
  assign t[21] = t[27] ^ x[6];
  assign t[22] = t[28] ^ x[11];
  assign t[23] = t[29] ^ x[16];
  assign t[24] = t[30] ^ x[21];
  assign t[25] = t[31] ^ x[26];
  assign t[26] = t[32] ^ x[31];
  assign t[27] = (~t[33] & t[34] & t[35] & t[36]) | (t[33] & ~t[35] & ~t[36]) | (t[33] & ~t[34] & ~t[36]) | (t[33] & ~t[34] & ~t[35]);
  assign t[28] = (~t[37] & t[38] & t[39] & t[40]) | (t[37] & ~t[39] & ~t[40]) | (t[37] & ~t[38] & ~t[40]) | (t[37] & ~t[38] & ~t[39]);
  assign t[29] = (~t[41] & t[42] & t[43] & t[44]) | (t[41] & ~t[43] & ~t[44]) | (t[41] & ~t[42] & ~t[44]) | (t[41] & ~t[42] & ~t[43]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[45] & t[46] & t[47] & t[48]) | (t[45] & ~t[47] & ~t[48]) | (t[45] & ~t[46] & ~t[48]) | (t[45] & ~t[46] & ~t[47]);
  assign t[31] = (~t[49] & t[50] & t[51] & t[52]) | (t[49] & ~t[51] & ~t[52]) | (t[49] & ~t[50] & ~t[52]) | (t[49] & ~t[50] & ~t[51]);
  assign t[32] = (~t[53] & t[54] & t[55] & t[56]) | (t[53] & ~t[55] & ~t[56]) | (t[53] & ~t[54] & ~t[56]) | (t[53] & ~t[54] & ~t[55]);
  assign t[33] = t[57] ^ x[6];
  assign t[34] = t[58] ^ x[3];
  assign t[35] = t[59] ^ x[4];
  assign t[36] = t[60] ^ x[5];
  assign t[37] = t[61] ^ x[11];
  assign t[38] = t[62] ^ x[8];
  assign t[39] = t[63] ^ x[9];
  assign t[3] = ~(t[4] ^ t[16]);
  assign t[40] = t[64] ^ x[10];
  assign t[41] = t[65] ^ x[16];
  assign t[42] = t[66] ^ x[13];
  assign t[43] = t[67] ^ x[14];
  assign t[44] = t[68] ^ x[15];
  assign t[45] = t[69] ^ x[21];
  assign t[46] = t[70] ^ x[18];
  assign t[47] = t[71] ^ x[19];
  assign t[48] = t[72] ^ x[20];
  assign t[49] = t[73] ^ x[26];
  assign t[4] = ~t[5];
  assign t[50] = t[74] ^ x[23];
  assign t[51] = t[75] ^ x[24];
  assign t[52] = t[76] ^ x[25];
  assign t[53] = t[77] ^ x[31];
  assign t[54] = t[78] ^ x[28];
  assign t[55] = t[79] ^ x[29];
  assign t[56] = t[80] ^ x[30];
  assign t[57] = (x[2]);
  assign t[58] = (x[2]);
  assign t[59] = (x[2]);
  assign t[5] = ~(t[6]);
  assign t[60] = (x[2]);
  assign t[61] = (x[7]);
  assign t[62] = (x[7]);
  assign t[63] = (x[7]);
  assign t[64] = (x[7]);
  assign t[65] = (x[12]);
  assign t[66] = (x[12]);
  assign t[67] = (x[12]);
  assign t[68] = (x[12]);
  assign t[69] = (x[17]);
  assign t[6] = t[7] ^ t[8];
  assign t[70] = (x[17]);
  assign t[71] = (x[17]);
  assign t[72] = (x[17]);
  assign t[73] = (x[22]);
  assign t[74] = (x[22]);
  assign t[75] = (x[22]);
  assign t[76] = (x[22]);
  assign t[77] = (x[27]);
  assign t[78] = (x[27]);
  assign t[79] = (x[27]);
  assign t[7] = t[9] ^ t[10];
  assign t[80] = (x[27]);
  assign t[8] = t[11] & t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = (t[0]);
endmodule

module R2ind223(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[11] & t[13];
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] ^ t[14];
  assign t[14] = t[18] ^ t[20];
  assign t[15] = (t[21]);
  assign t[16] = (t[22]);
  assign t[17] = (t[23]);
  assign t[18] = (t[24]);
  assign t[19] = (t[25]);
  assign t[1] = ~(t[2] ^ t[15]);
  assign t[20] = (t[26]);
  assign t[21] = t[27] ^ x[6];
  assign t[22] = t[28] ^ x[11];
  assign t[23] = t[29] ^ x[16];
  assign t[24] = t[30] ^ x[21];
  assign t[25] = t[31] ^ x[26];
  assign t[26] = t[32] ^ x[31];
  assign t[27] = (~t[33] & t[34] & t[35] & t[36]) | (t[33] & ~t[35] & ~t[36]) | (t[33] & ~t[34] & ~t[36]) | (t[33] & ~t[34] & ~t[35]);
  assign t[28] = (~t[37] & t[38] & t[39] & t[40]) | (t[37] & ~t[39] & ~t[40]) | (t[37] & ~t[38] & ~t[40]) | (t[37] & ~t[38] & ~t[39]);
  assign t[29] = (~t[41] & t[42] & t[43] & t[44]) | (t[41] & ~t[43] & ~t[44]) | (t[41] & ~t[42] & ~t[44]) | (t[41] & ~t[42] & ~t[43]);
  assign t[2] = ~t[3];
  assign t[30] = (~t[45] & t[46] & t[47] & t[48]) | (t[45] & ~t[47] & ~t[48]) | (t[45] & ~t[46] & ~t[48]) | (t[45] & ~t[46] & ~t[47]);
  assign t[31] = (~t[49] & t[50] & t[51] & t[52]) | (t[49] & ~t[51] & ~t[52]) | (t[49] & ~t[50] & ~t[52]) | (t[49] & ~t[50] & ~t[51]);
  assign t[32] = (~t[53] & t[54] & t[55] & t[56]) | (t[53] & ~t[55] & ~t[56]) | (t[53] & ~t[54] & ~t[56]) | (t[53] & ~t[54] & ~t[55]);
  assign t[33] = t[57] ^ x[6];
  assign t[34] = t[58] ^ x[3];
  assign t[35] = t[59] ^ x[4];
  assign t[36] = t[60] ^ x[5];
  assign t[37] = t[61] ^ x[11];
  assign t[38] = t[62] ^ x[8];
  assign t[39] = t[63] ^ x[9];
  assign t[3] = ~(t[4] ^ t[16]);
  assign t[40] = t[64] ^ x[10];
  assign t[41] = t[65] ^ x[16];
  assign t[42] = t[66] ^ x[13];
  assign t[43] = t[67] ^ x[14];
  assign t[44] = t[68] ^ x[15];
  assign t[45] = t[69] ^ x[21];
  assign t[46] = t[70] ^ x[18];
  assign t[47] = t[71] ^ x[19];
  assign t[48] = t[72] ^ x[20];
  assign t[49] = t[73] ^ x[26];
  assign t[4] = ~t[5];
  assign t[50] = t[74] ^ x[23];
  assign t[51] = t[75] ^ x[24];
  assign t[52] = t[76] ^ x[25];
  assign t[53] = t[77] ^ x[31];
  assign t[54] = t[78] ^ x[28];
  assign t[55] = t[79] ^ x[29];
  assign t[56] = t[80] ^ x[30];
  assign t[57] = (x[2]);
  assign t[58] = (x[2]);
  assign t[59] = (x[2]);
  assign t[5] = ~(t[6]);
  assign t[60] = (x[2]);
  assign t[61] = (x[7]);
  assign t[62] = (x[7]);
  assign t[63] = (x[7]);
  assign t[64] = (x[7]);
  assign t[65] = (x[12]);
  assign t[66] = (x[12]);
  assign t[67] = (x[12]);
  assign t[68] = (x[12]);
  assign t[69] = (x[17]);
  assign t[6] = t[7] ^ t[8];
  assign t[70] = (x[17]);
  assign t[71] = (x[17]);
  assign t[72] = (x[17]);
  assign t[73] = (x[22]);
  assign t[74] = (x[22]);
  assign t[75] = (x[22]);
  assign t[76] = (x[22]);
  assign t[77] = (x[27]);
  assign t[78] = (x[27]);
  assign t[79] = (x[27]);
  assign t[7] = t[9] ^ t[10];
  assign t[80] = (x[27]);
  assign t[8] = t[11] & t[12];
  assign t[9] = t[17] ^ t[18];
  assign y = (t[0]);
endmodule

module R2ind224(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[54] & t[26];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[55] & t[31];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[56] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[54] ^ t[27]);
  assign t[29] = t[58] ^ t[57];
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[55] ^ t[32]);
  assign t[34] = t[60] ^ t[59];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[56] ^ t[37]);
  assign t[39] = t[62] ^ t[61];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[54] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[54] ^ t[50];
  assign t[44] = t[55] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[55] ^ t[51];
  assign t[47] = t[56] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[56] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[57] ^ t[63];
  assign t[51] = t[59] ^ t[64];
  assign t[52] = t[61] ^ t[65];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] & t[17];
  assign y = (t[0]);
endmodule

module R2ind225(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[54] & t[26];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[55] & t[31];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[56] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[54] ^ t[27]);
  assign t[29] = t[58] ^ t[57];
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[55] ^ t[32]);
  assign t[34] = t[60] ^ t[59];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[56] ^ t[37]);
  assign t[39] = t[62] ^ t[61];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[54] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[54] ^ t[50];
  assign t[44] = t[55] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[55] ^ t[51];
  assign t[47] = t[56] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[56] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[57] ^ t[63];
  assign t[51] = t[59] ^ t[64];
  assign t[52] = t[61] ^ t[65];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] & t[17];
  assign y = (t[0]);
endmodule

module R2ind226(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[54] & t[26];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[55] & t[31];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[56] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[54] ^ t[27]);
  assign t[29] = t[58] ^ t[57];
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[55] ^ t[32]);
  assign t[34] = t[60] ^ t[59];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[56] ^ t[37]);
  assign t[39] = t[62] ^ t[61];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[54] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[54] ^ t[50];
  assign t[44] = t[55] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[55] ^ t[51];
  assign t[47] = t[56] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[56] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[57] ^ t[63];
  assign t[51] = t[59] ^ t[64];
  assign t[52] = t[61] ^ t[65];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] & t[17];
  assign y = (t[0]);
endmodule

module R2ind227(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[54] & t[26];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[55] & t[31];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[56] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[54] ^ t[27]);
  assign t[29] = t[58] ^ t[57];
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[55] ^ t[32]);
  assign t[34] = t[60] ^ t[59];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[56] ^ t[37]);
  assign t[39] = t[62] ^ t[61];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[54] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[54] ^ t[50];
  assign t[44] = t[55] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[55] ^ t[51];
  assign t[47] = t[56] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[56] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[57] ^ t[63];
  assign t[51] = t[59] ^ t[64];
  assign t[52] = t[61] ^ t[65];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] & t[17];
  assign y = (t[0]);
endmodule

module R2ind228(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[26] ^ t[27];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[28] & t[29];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[30] ^ t[15];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[54] ^ t[28];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[31] ^ t[32];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[55] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[56] ^ t[38];
  assign t[26] = t[57] ^ t[58];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[58]);
  assign t[29] = ~(t[54] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = t[54] & t[42];
  assign t[31] = t[59] ^ t[60];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[60]);
  assign t[34] = ~(t[55] ^ t[33]);
  assign t[35] = t[55] & t[44];
  assign t[36] = t[61] ^ t[62];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[62]);
  assign t[39] = ~(t[56] ^ t[38]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[56] & t[46];
  assign t[41] = t[54] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[55] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[56] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[58] ^ t[63];
  assign t[48] = t[54] ^ t[26];
  assign t[49] = t[60] ^ t[64];
  assign t[4] = ~t[7];
  assign t[50] = t[55] ^ t[31];
  assign t[51] = t[62] ^ t[65];
  assign t[52] = t[56] ^ t[36];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind229(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[26] ^ t[27];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[28] & t[29];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[30] ^ t[15];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[54] ^ t[28];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[31] ^ t[32];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[55] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[56] ^ t[38];
  assign t[26] = t[57] ^ t[58];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[58]);
  assign t[29] = ~(t[54] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = t[54] & t[42];
  assign t[31] = t[59] ^ t[60];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[60]);
  assign t[34] = ~(t[55] ^ t[33]);
  assign t[35] = t[55] & t[44];
  assign t[36] = t[61] ^ t[62];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[62]);
  assign t[39] = ~(t[56] ^ t[38]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[56] & t[46];
  assign t[41] = t[54] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[55] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[56] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[58] ^ t[63];
  assign t[48] = t[54] ^ t[26];
  assign t[49] = t[60] ^ t[64];
  assign t[4] = ~t[7];
  assign t[50] = t[55] ^ t[31];
  assign t[51] = t[62] ^ t[65];
  assign t[52] = t[56] ^ t[36];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind230(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[26] ^ t[27];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[28] & t[29];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[30] ^ t[15];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[54] ^ t[28];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[31] ^ t[32];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[55] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[56] ^ t[38];
  assign t[26] = t[57] ^ t[58];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[58]);
  assign t[29] = ~(t[54] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = t[54] & t[42];
  assign t[31] = t[59] ^ t[60];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[60]);
  assign t[34] = ~(t[55] ^ t[33]);
  assign t[35] = t[55] & t[44];
  assign t[36] = t[61] ^ t[62];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[62]);
  assign t[39] = ~(t[56] ^ t[38]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[56] & t[46];
  assign t[41] = t[54] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[55] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[56] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[58] ^ t[63];
  assign t[48] = t[54] ^ t[26];
  assign t[49] = t[60] ^ t[64];
  assign t[4] = ~t[7];
  assign t[50] = t[55] ^ t[31];
  assign t[51] = t[62] ^ t[65];
  assign t[52] = t[56] ^ t[36];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind231(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[26] ^ t[27];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[28] & t[29];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[30] ^ t[15];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[54] ^ t[28];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[31] ^ t[32];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[55] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[56] ^ t[38];
  assign t[26] = t[57] ^ t[58];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[58]);
  assign t[29] = ~(t[54] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = t[54] & t[42];
  assign t[31] = t[59] ^ t[60];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[60]);
  assign t[34] = ~(t[55] ^ t[33]);
  assign t[35] = t[55] & t[44];
  assign t[36] = t[61] ^ t[62];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[62]);
  assign t[39] = ~(t[56] ^ t[38]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[56] & t[46];
  assign t[41] = t[54] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[55] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[56] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[58] ^ t[63];
  assign t[48] = t[54] ^ t[26];
  assign t[49] = t[60] ^ t[64];
  assign t[4] = ~t[7];
  assign t[50] = t[55] ^ t[31];
  assign t[51] = t[62] ^ t[65];
  assign t[52] = t[56] ^ t[36];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind232(x, y);
 input [51:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[7]);
  assign t[101] = (x[12]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[17]);
  assign t[106] = (x[17]);
  assign t[107] = (x[17]);
  assign t[108] = (x[17]);
  assign t[109] = (x[22]);
  assign t[10] = t[15] ^ t[16];
  assign t[110] = (x[22]);
  assign t[111] = (x[22]);
  assign t[112] = (x[22]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[32]);
  assign t[118] = (x[32]);
  assign t[119] = (x[32]);
  assign t[11] = t[24] ^ t[25];
  assign t[120] = (x[32]);
  assign t[121] = (x[37]);
  assign t[122] = (x[37]);
  assign t[123] = (x[37]);
  assign t[124] = (x[37]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[127] = (x[42]);
  assign t[128] = (x[42]);
  assign t[129] = (x[47]);
  assign t[12] = t[17] & t[18];
  assign t[130] = (x[47]);
  assign t[131] = (x[47]);
  assign t[132] = (x[47]);
  assign t[13] = t[26] ^ t[27];
  assign t[14] = t[19] & t[20];
  assign t[15] = t[28] ^ t[29];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[30] ^ t[17]);
  assign t[19] = ~(t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] ^ t[19]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[23]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = t[43] ^ x[6];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[21];
  assign t[37] = t[47] ^ x[26];
  assign t[38] = t[48] ^ x[31];
  assign t[39] = t[49] ^ x[36];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[41];
  assign t[41] = t[51] ^ x[46];
  assign t[42] = t[52] ^ x[51];
  assign t[43] = (~t[53] & t[54] & t[55] & t[56]) | (t[53] & ~t[55] & ~t[56]) | (t[53] & ~t[54] & ~t[56]) | (t[53] & ~t[54] & ~t[55]);
  assign t[44] = (~t[57] & t[58] & t[59] & t[60]) | (t[57] & ~t[59] & ~t[60]) | (t[57] & ~t[58] & ~t[60]) | (t[57] & ~t[58] & ~t[59]);
  assign t[45] = (~t[61] & t[62] & t[63] & t[64]) | (t[61] & ~t[63] & ~t[64]) | (t[61] & ~t[62] & ~t[64]) | (t[61] & ~t[62] & ~t[63]);
  assign t[46] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[47] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[48] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[49] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[51] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[52] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[53] = t[93] ^ x[6];
  assign t[54] = t[94] ^ x[3];
  assign t[55] = t[95] ^ x[4];
  assign t[56] = t[96] ^ x[5];
  assign t[57] = t[97] ^ x[11];
  assign t[58] = t[98] ^ x[8];
  assign t[59] = t[99] ^ x[9];
  assign t[5] = ~(t[8]);
  assign t[60] = t[100] ^ x[10];
  assign t[61] = t[101] ^ x[16];
  assign t[62] = t[102] ^ x[13];
  assign t[63] = t[103] ^ x[14];
  assign t[64] = t[104] ^ x[15];
  assign t[65] = t[105] ^ x[21];
  assign t[66] = t[106] ^ x[18];
  assign t[67] = t[107] ^ x[19];
  assign t[68] = t[108] ^ x[20];
  assign t[69] = t[109] ^ x[26];
  assign t[6] = ~(t[9]);
  assign t[70] = t[110] ^ x[23];
  assign t[71] = t[111] ^ x[24];
  assign t[72] = t[112] ^ x[25];
  assign t[73] = t[113] ^ x[31];
  assign t[74] = t[114] ^ x[28];
  assign t[75] = t[115] ^ x[29];
  assign t[76] = t[116] ^ x[30];
  assign t[77] = t[117] ^ x[36];
  assign t[78] = t[118] ^ x[33];
  assign t[79] = t[119] ^ x[34];
  assign t[7] = ~(t[10]);
  assign t[80] = t[120] ^ x[35];
  assign t[81] = t[121] ^ x[41];
  assign t[82] = t[122] ^ x[38];
  assign t[83] = t[123] ^ x[39];
  assign t[84] = t[124] ^ x[40];
  assign t[85] = t[125] ^ x[46];
  assign t[86] = t[126] ^ x[43];
  assign t[87] = t[127] ^ x[44];
  assign t[88] = t[128] ^ x[45];
  assign t[89] = t[129] ^ x[51];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[130] ^ x[48];
  assign t[91] = t[131] ^ x[49];
  assign t[92] = t[132] ^ x[50];
  assign t[93] = (x[2]);
  assign t[94] = (x[2]);
  assign t[95] = (x[2]);
  assign t[96] = (x[2]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[7]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind233(x, y);
 input [51:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[7]);
  assign t[101] = (x[12]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[17]);
  assign t[106] = (x[17]);
  assign t[107] = (x[17]);
  assign t[108] = (x[17]);
  assign t[109] = (x[22]);
  assign t[10] = t[15] ^ t[16];
  assign t[110] = (x[22]);
  assign t[111] = (x[22]);
  assign t[112] = (x[22]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[32]);
  assign t[118] = (x[32]);
  assign t[119] = (x[32]);
  assign t[11] = t[24] ^ t[25];
  assign t[120] = (x[32]);
  assign t[121] = (x[37]);
  assign t[122] = (x[37]);
  assign t[123] = (x[37]);
  assign t[124] = (x[37]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[127] = (x[42]);
  assign t[128] = (x[42]);
  assign t[129] = (x[47]);
  assign t[12] = t[17] & t[18];
  assign t[130] = (x[47]);
  assign t[131] = (x[47]);
  assign t[132] = (x[47]);
  assign t[13] = t[26] ^ t[27];
  assign t[14] = t[19] & t[20];
  assign t[15] = t[28] ^ t[29];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[30] ^ t[17]);
  assign t[19] = ~(t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] ^ t[19]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[23]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = t[43] ^ x[6];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[21];
  assign t[37] = t[47] ^ x[26];
  assign t[38] = t[48] ^ x[31];
  assign t[39] = t[49] ^ x[36];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[41];
  assign t[41] = t[51] ^ x[46];
  assign t[42] = t[52] ^ x[51];
  assign t[43] = (~t[53] & t[54] & t[55] & t[56]) | (t[53] & ~t[55] & ~t[56]) | (t[53] & ~t[54] & ~t[56]) | (t[53] & ~t[54] & ~t[55]);
  assign t[44] = (~t[57] & t[58] & t[59] & t[60]) | (t[57] & ~t[59] & ~t[60]) | (t[57] & ~t[58] & ~t[60]) | (t[57] & ~t[58] & ~t[59]);
  assign t[45] = (~t[61] & t[62] & t[63] & t[64]) | (t[61] & ~t[63] & ~t[64]) | (t[61] & ~t[62] & ~t[64]) | (t[61] & ~t[62] & ~t[63]);
  assign t[46] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[47] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[48] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[49] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[51] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[52] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[53] = t[93] ^ x[6];
  assign t[54] = t[94] ^ x[3];
  assign t[55] = t[95] ^ x[4];
  assign t[56] = t[96] ^ x[5];
  assign t[57] = t[97] ^ x[11];
  assign t[58] = t[98] ^ x[8];
  assign t[59] = t[99] ^ x[9];
  assign t[5] = ~(t[8]);
  assign t[60] = t[100] ^ x[10];
  assign t[61] = t[101] ^ x[16];
  assign t[62] = t[102] ^ x[13];
  assign t[63] = t[103] ^ x[14];
  assign t[64] = t[104] ^ x[15];
  assign t[65] = t[105] ^ x[21];
  assign t[66] = t[106] ^ x[18];
  assign t[67] = t[107] ^ x[19];
  assign t[68] = t[108] ^ x[20];
  assign t[69] = t[109] ^ x[26];
  assign t[6] = ~(t[9]);
  assign t[70] = t[110] ^ x[23];
  assign t[71] = t[111] ^ x[24];
  assign t[72] = t[112] ^ x[25];
  assign t[73] = t[113] ^ x[31];
  assign t[74] = t[114] ^ x[28];
  assign t[75] = t[115] ^ x[29];
  assign t[76] = t[116] ^ x[30];
  assign t[77] = t[117] ^ x[36];
  assign t[78] = t[118] ^ x[33];
  assign t[79] = t[119] ^ x[34];
  assign t[7] = ~(t[10]);
  assign t[80] = t[120] ^ x[35];
  assign t[81] = t[121] ^ x[41];
  assign t[82] = t[122] ^ x[38];
  assign t[83] = t[123] ^ x[39];
  assign t[84] = t[124] ^ x[40];
  assign t[85] = t[125] ^ x[46];
  assign t[86] = t[126] ^ x[43];
  assign t[87] = t[127] ^ x[44];
  assign t[88] = t[128] ^ x[45];
  assign t[89] = t[129] ^ x[51];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[130] ^ x[48];
  assign t[91] = t[131] ^ x[49];
  assign t[92] = t[132] ^ x[50];
  assign t[93] = (x[2]);
  assign t[94] = (x[2]);
  assign t[95] = (x[2]);
  assign t[96] = (x[2]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[7]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind234(x, y);
 input [51:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[7]);
  assign t[101] = (x[12]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[17]);
  assign t[106] = (x[17]);
  assign t[107] = (x[17]);
  assign t[108] = (x[17]);
  assign t[109] = (x[22]);
  assign t[10] = t[15] ^ t[16];
  assign t[110] = (x[22]);
  assign t[111] = (x[22]);
  assign t[112] = (x[22]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[32]);
  assign t[118] = (x[32]);
  assign t[119] = (x[32]);
  assign t[11] = t[24] ^ t[25];
  assign t[120] = (x[32]);
  assign t[121] = (x[37]);
  assign t[122] = (x[37]);
  assign t[123] = (x[37]);
  assign t[124] = (x[37]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[127] = (x[42]);
  assign t[128] = (x[42]);
  assign t[129] = (x[47]);
  assign t[12] = t[17] & t[18];
  assign t[130] = (x[47]);
  assign t[131] = (x[47]);
  assign t[132] = (x[47]);
  assign t[13] = t[26] ^ t[27];
  assign t[14] = t[19] & t[20];
  assign t[15] = t[28] ^ t[29];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[30] ^ t[17]);
  assign t[19] = ~(t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] ^ t[19]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[23]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = t[43] ^ x[6];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[21];
  assign t[37] = t[47] ^ x[26];
  assign t[38] = t[48] ^ x[31];
  assign t[39] = t[49] ^ x[36];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[41];
  assign t[41] = t[51] ^ x[46];
  assign t[42] = t[52] ^ x[51];
  assign t[43] = (~t[53] & t[54] & t[55] & t[56]) | (t[53] & ~t[55] & ~t[56]) | (t[53] & ~t[54] & ~t[56]) | (t[53] & ~t[54] & ~t[55]);
  assign t[44] = (~t[57] & t[58] & t[59] & t[60]) | (t[57] & ~t[59] & ~t[60]) | (t[57] & ~t[58] & ~t[60]) | (t[57] & ~t[58] & ~t[59]);
  assign t[45] = (~t[61] & t[62] & t[63] & t[64]) | (t[61] & ~t[63] & ~t[64]) | (t[61] & ~t[62] & ~t[64]) | (t[61] & ~t[62] & ~t[63]);
  assign t[46] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[47] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[48] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[49] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[51] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[52] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[53] = t[93] ^ x[6];
  assign t[54] = t[94] ^ x[3];
  assign t[55] = t[95] ^ x[4];
  assign t[56] = t[96] ^ x[5];
  assign t[57] = t[97] ^ x[11];
  assign t[58] = t[98] ^ x[8];
  assign t[59] = t[99] ^ x[9];
  assign t[5] = ~(t[8]);
  assign t[60] = t[100] ^ x[10];
  assign t[61] = t[101] ^ x[16];
  assign t[62] = t[102] ^ x[13];
  assign t[63] = t[103] ^ x[14];
  assign t[64] = t[104] ^ x[15];
  assign t[65] = t[105] ^ x[21];
  assign t[66] = t[106] ^ x[18];
  assign t[67] = t[107] ^ x[19];
  assign t[68] = t[108] ^ x[20];
  assign t[69] = t[109] ^ x[26];
  assign t[6] = ~(t[9]);
  assign t[70] = t[110] ^ x[23];
  assign t[71] = t[111] ^ x[24];
  assign t[72] = t[112] ^ x[25];
  assign t[73] = t[113] ^ x[31];
  assign t[74] = t[114] ^ x[28];
  assign t[75] = t[115] ^ x[29];
  assign t[76] = t[116] ^ x[30];
  assign t[77] = t[117] ^ x[36];
  assign t[78] = t[118] ^ x[33];
  assign t[79] = t[119] ^ x[34];
  assign t[7] = ~(t[10]);
  assign t[80] = t[120] ^ x[35];
  assign t[81] = t[121] ^ x[41];
  assign t[82] = t[122] ^ x[38];
  assign t[83] = t[123] ^ x[39];
  assign t[84] = t[124] ^ x[40];
  assign t[85] = t[125] ^ x[46];
  assign t[86] = t[126] ^ x[43];
  assign t[87] = t[127] ^ x[44];
  assign t[88] = t[128] ^ x[45];
  assign t[89] = t[129] ^ x[51];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[130] ^ x[48];
  assign t[91] = t[131] ^ x[49];
  assign t[92] = t[132] ^ x[50];
  assign t[93] = (x[2]);
  assign t[94] = (x[2]);
  assign t[95] = (x[2]);
  assign t[96] = (x[2]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[7]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind235(x, y);
 input [51:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[7]);
  assign t[101] = (x[12]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[17]);
  assign t[106] = (x[17]);
  assign t[107] = (x[17]);
  assign t[108] = (x[17]);
  assign t[109] = (x[22]);
  assign t[10] = t[15] ^ t[16];
  assign t[110] = (x[22]);
  assign t[111] = (x[22]);
  assign t[112] = (x[22]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[32]);
  assign t[118] = (x[32]);
  assign t[119] = (x[32]);
  assign t[11] = t[24] ^ t[25];
  assign t[120] = (x[32]);
  assign t[121] = (x[37]);
  assign t[122] = (x[37]);
  assign t[123] = (x[37]);
  assign t[124] = (x[37]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[127] = (x[42]);
  assign t[128] = (x[42]);
  assign t[129] = (x[47]);
  assign t[12] = t[17] & t[18];
  assign t[130] = (x[47]);
  assign t[131] = (x[47]);
  assign t[132] = (x[47]);
  assign t[13] = t[26] ^ t[27];
  assign t[14] = t[19] & t[20];
  assign t[15] = t[28] ^ t[29];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[30] ^ t[17]);
  assign t[19] = ~(t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] ^ t[19]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[23]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = t[43] ^ x[6];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[21];
  assign t[37] = t[47] ^ x[26];
  assign t[38] = t[48] ^ x[31];
  assign t[39] = t[49] ^ x[36];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[41];
  assign t[41] = t[51] ^ x[46];
  assign t[42] = t[52] ^ x[51];
  assign t[43] = (~t[53] & t[54] & t[55] & t[56]) | (t[53] & ~t[55] & ~t[56]) | (t[53] & ~t[54] & ~t[56]) | (t[53] & ~t[54] & ~t[55]);
  assign t[44] = (~t[57] & t[58] & t[59] & t[60]) | (t[57] & ~t[59] & ~t[60]) | (t[57] & ~t[58] & ~t[60]) | (t[57] & ~t[58] & ~t[59]);
  assign t[45] = (~t[61] & t[62] & t[63] & t[64]) | (t[61] & ~t[63] & ~t[64]) | (t[61] & ~t[62] & ~t[64]) | (t[61] & ~t[62] & ~t[63]);
  assign t[46] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[47] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[48] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[49] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[51] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[52] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[53] = t[93] ^ x[6];
  assign t[54] = t[94] ^ x[3];
  assign t[55] = t[95] ^ x[4];
  assign t[56] = t[96] ^ x[5];
  assign t[57] = t[97] ^ x[11];
  assign t[58] = t[98] ^ x[8];
  assign t[59] = t[99] ^ x[9];
  assign t[5] = ~(t[8]);
  assign t[60] = t[100] ^ x[10];
  assign t[61] = t[101] ^ x[16];
  assign t[62] = t[102] ^ x[13];
  assign t[63] = t[103] ^ x[14];
  assign t[64] = t[104] ^ x[15];
  assign t[65] = t[105] ^ x[21];
  assign t[66] = t[106] ^ x[18];
  assign t[67] = t[107] ^ x[19];
  assign t[68] = t[108] ^ x[20];
  assign t[69] = t[109] ^ x[26];
  assign t[6] = ~(t[9]);
  assign t[70] = t[110] ^ x[23];
  assign t[71] = t[111] ^ x[24];
  assign t[72] = t[112] ^ x[25];
  assign t[73] = t[113] ^ x[31];
  assign t[74] = t[114] ^ x[28];
  assign t[75] = t[115] ^ x[29];
  assign t[76] = t[116] ^ x[30];
  assign t[77] = t[117] ^ x[36];
  assign t[78] = t[118] ^ x[33];
  assign t[79] = t[119] ^ x[34];
  assign t[7] = ~(t[10]);
  assign t[80] = t[120] ^ x[35];
  assign t[81] = t[121] ^ x[41];
  assign t[82] = t[122] ^ x[38];
  assign t[83] = t[123] ^ x[39];
  assign t[84] = t[124] ^ x[40];
  assign t[85] = t[125] ^ x[46];
  assign t[86] = t[126] ^ x[43];
  assign t[87] = t[127] ^ x[44];
  assign t[88] = t[128] ^ x[45];
  assign t[89] = t[129] ^ x[51];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[130] ^ x[48];
  assign t[91] = t[131] ^ x[49];
  assign t[92] = t[132] ^ x[50];
  assign t[93] = (x[2]);
  assign t[94] = (x[2]);
  assign t[95] = (x[2]);
  assign t[96] = (x[2]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[7]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind236(x, y);
 input [66:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[34];
  assign t[101] = t[153] ^ x[35];
  assign t[102] = t[154] ^ x[41];
  assign t[103] = t[155] ^ x[38];
  assign t[104] = t[156] ^ x[39];
  assign t[105] = t[157] ^ x[40];
  assign t[106] = t[158] ^ x[46];
  assign t[107] = t[159] ^ x[43];
  assign t[108] = t[160] ^ x[44];
  assign t[109] = t[161] ^ x[45];
  assign t[10] = t[15] ^ t[16];
  assign t[110] = t[162] ^ x[51];
  assign t[111] = t[163] ^ x[48];
  assign t[112] = t[164] ^ x[49];
  assign t[113] = t[165] ^ x[50];
  assign t[114] = t[166] ^ x[56];
  assign t[115] = t[167] ^ x[53];
  assign t[116] = t[168] ^ x[54];
  assign t[117] = t[169] ^ x[55];
  assign t[118] = t[170] ^ x[61];
  assign t[119] = t[171] ^ x[58];
  assign t[11] = t[17] ^ t[18];
  assign t[120] = t[172] ^ x[59];
  assign t[121] = t[173] ^ x[60];
  assign t[122] = t[174] ^ x[66];
  assign t[123] = t[175] ^ x[63];
  assign t[124] = t[176] ^ x[64];
  assign t[125] = t[177] ^ x[65];
  assign t[126] = (x[2]);
  assign t[127] = (x[2]);
  assign t[128] = (x[2]);
  assign t[129] = (x[2]);
  assign t[12] = t[19] & t[20];
  assign t[130] = (x[7]);
  assign t[131] = (x[7]);
  assign t[132] = (x[7]);
  assign t[133] = (x[7]);
  assign t[134] = (x[12]);
  assign t[135] = (x[12]);
  assign t[136] = (x[12]);
  assign t[137] = (x[12]);
  assign t[138] = (x[17]);
  assign t[139] = (x[17]);
  assign t[13] = t[21] ^ t[22];
  assign t[140] = (x[17]);
  assign t[141] = (x[17]);
  assign t[142] = (x[22]);
  assign t[143] = (x[22]);
  assign t[144] = (x[22]);
  assign t[145] = (x[22]);
  assign t[146] = (x[27]);
  assign t[147] = (x[27]);
  assign t[148] = (x[27]);
  assign t[149] = (x[27]);
  assign t[14] = t[23] & t[24];
  assign t[150] = (x[32]);
  assign t[151] = (x[32]);
  assign t[152] = (x[32]);
  assign t[153] = (x[32]);
  assign t[154] = (x[37]);
  assign t[155] = (x[37]);
  assign t[156] = (x[37]);
  assign t[157] = (x[37]);
  assign t[158] = (x[42]);
  assign t[159] = (x[42]);
  assign t[15] = t[25] ^ t[26];
  assign t[160] = (x[42]);
  assign t[161] = (x[42]);
  assign t[162] = (x[47]);
  assign t[163] = (x[47]);
  assign t[164] = (x[47]);
  assign t[165] = (x[47]);
  assign t[166] = (x[52]);
  assign t[167] = (x[52]);
  assign t[168] = (x[52]);
  assign t[169] = (x[52]);
  assign t[16] = t[27] & t[28];
  assign t[170] = (x[57]);
  assign t[171] = (x[57]);
  assign t[172] = (x[57]);
  assign t[173] = (x[57]);
  assign t[174] = (x[62]);
  assign t[175] = (x[62]);
  assign t[176] = (x[62]);
  assign t[177] = (x[62]);
  assign t[17] = t[36] ^ t[37];
  assign t[18] = t[19] & t[29];
  assign t[19] = ~(t[37]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[38] ^ t[19]);
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[23] & t[30];
  assign t[23] = ~(t[40]);
  assign t[24] = ~(t[41] ^ t[23]);
  assign t[25] = t[42] ^ t[43];
  assign t[26] = t[27] & t[31];
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[44] ^ t[27]);
  assign t[29] = t[38] ^ t[32];
  assign t[2] = ~(t[4] ^ t[35]);
  assign t[30] = t[41] ^ t[33];
  assign t[31] = t[44] ^ t[34];
  assign t[32] = t[37] ^ t[45];
  assign t[33] = t[40] ^ t[46];
  assign t[34] = t[43] ^ t[47];
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = t[61] ^ x[6];
  assign t[49] = t[62] ^ x[11];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ x[16];
  assign t[51] = t[64] ^ x[21];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[31];
  assign t[54] = t[67] ^ x[36];
  assign t[55] = t[68] ^ x[41];
  assign t[56] = t[69] ^ x[46];
  assign t[57] = t[70] ^ x[51];
  assign t[58] = t[71] ^ x[56];
  assign t[59] = t[72] ^ x[61];
  assign t[5] = ~(t[8]);
  assign t[60] = t[73] ^ x[66];
  assign t[61] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[62] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[63] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[64] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[65] = (~t[90] & t[91] & t[92] & t[93]) | (t[90] & ~t[92] & ~t[93]) | (t[90] & ~t[91] & ~t[93]) | (t[90] & ~t[91] & ~t[92]);
  assign t[66] = (~t[94] & t[95] & t[96] & t[97]) | (t[94] & ~t[96] & ~t[97]) | (t[94] & ~t[95] & ~t[97]) | (t[94] & ~t[95] & ~t[96]);
  assign t[67] = (~t[98] & t[99] & t[100] & t[101]) | (t[98] & ~t[100] & ~t[101]) | (t[98] & ~t[99] & ~t[101]) | (t[98] & ~t[99] & ~t[100]);
  assign t[68] = (~t[102] & t[103] & t[104] & t[105]) | (t[102] & ~t[104] & ~t[105]) | (t[102] & ~t[103] & ~t[105]) | (t[102] & ~t[103] & ~t[104]);
  assign t[69] = (~t[106] & t[107] & t[108] & t[109]) | (t[106] & ~t[108] & ~t[109]) | (t[106] & ~t[107] & ~t[109]) | (t[106] & ~t[107] & ~t[108]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[110] & t[111] & t[112] & t[113]) | (t[110] & ~t[112] & ~t[113]) | (t[110] & ~t[111] & ~t[113]) | (t[110] & ~t[111] & ~t[112]);
  assign t[71] = (~t[114] & t[115] & t[116] & t[117]) | (t[114] & ~t[116] & ~t[117]) | (t[114] & ~t[115] & ~t[117]) | (t[114] & ~t[115] & ~t[116]);
  assign t[72] = (~t[118] & t[119] & t[120] & t[121]) | (t[118] & ~t[120] & ~t[121]) | (t[118] & ~t[119] & ~t[121]) | (t[118] & ~t[119] & ~t[120]);
  assign t[73] = (~t[122] & t[123] & t[124] & t[125]) | (t[122] & ~t[124] & ~t[125]) | (t[122] & ~t[123] & ~t[125]) | (t[122] & ~t[123] & ~t[124]);
  assign t[74] = t[126] ^ x[6];
  assign t[75] = t[127] ^ x[3];
  assign t[76] = t[128] ^ x[4];
  assign t[77] = t[129] ^ x[5];
  assign t[78] = t[130] ^ x[11];
  assign t[79] = t[131] ^ x[8];
  assign t[7] = ~(t[10]);
  assign t[80] = t[132] ^ x[9];
  assign t[81] = t[133] ^ x[10];
  assign t[82] = t[134] ^ x[16];
  assign t[83] = t[135] ^ x[13];
  assign t[84] = t[136] ^ x[14];
  assign t[85] = t[137] ^ x[15];
  assign t[86] = t[138] ^ x[21];
  assign t[87] = t[139] ^ x[18];
  assign t[88] = t[140] ^ x[19];
  assign t[89] = t[141] ^ x[20];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[142] ^ x[26];
  assign t[91] = t[143] ^ x[23];
  assign t[92] = t[144] ^ x[24];
  assign t[93] = t[145] ^ x[25];
  assign t[94] = t[146] ^ x[31];
  assign t[95] = t[147] ^ x[28];
  assign t[96] = t[148] ^ x[29];
  assign t[97] = t[149] ^ x[30];
  assign t[98] = t[150] ^ x[36];
  assign t[99] = t[151] ^ x[33];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind237(x, y);
 input [66:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[34];
  assign t[101] = t[153] ^ x[35];
  assign t[102] = t[154] ^ x[41];
  assign t[103] = t[155] ^ x[38];
  assign t[104] = t[156] ^ x[39];
  assign t[105] = t[157] ^ x[40];
  assign t[106] = t[158] ^ x[46];
  assign t[107] = t[159] ^ x[43];
  assign t[108] = t[160] ^ x[44];
  assign t[109] = t[161] ^ x[45];
  assign t[10] = t[15] ^ t[16];
  assign t[110] = t[162] ^ x[51];
  assign t[111] = t[163] ^ x[48];
  assign t[112] = t[164] ^ x[49];
  assign t[113] = t[165] ^ x[50];
  assign t[114] = t[166] ^ x[56];
  assign t[115] = t[167] ^ x[53];
  assign t[116] = t[168] ^ x[54];
  assign t[117] = t[169] ^ x[55];
  assign t[118] = t[170] ^ x[61];
  assign t[119] = t[171] ^ x[58];
  assign t[11] = t[17] ^ t[18];
  assign t[120] = t[172] ^ x[59];
  assign t[121] = t[173] ^ x[60];
  assign t[122] = t[174] ^ x[66];
  assign t[123] = t[175] ^ x[63];
  assign t[124] = t[176] ^ x[64];
  assign t[125] = t[177] ^ x[65];
  assign t[126] = (x[2]);
  assign t[127] = (x[2]);
  assign t[128] = (x[2]);
  assign t[129] = (x[2]);
  assign t[12] = t[19] & t[20];
  assign t[130] = (x[7]);
  assign t[131] = (x[7]);
  assign t[132] = (x[7]);
  assign t[133] = (x[7]);
  assign t[134] = (x[12]);
  assign t[135] = (x[12]);
  assign t[136] = (x[12]);
  assign t[137] = (x[12]);
  assign t[138] = (x[17]);
  assign t[139] = (x[17]);
  assign t[13] = t[21] ^ t[22];
  assign t[140] = (x[17]);
  assign t[141] = (x[17]);
  assign t[142] = (x[22]);
  assign t[143] = (x[22]);
  assign t[144] = (x[22]);
  assign t[145] = (x[22]);
  assign t[146] = (x[27]);
  assign t[147] = (x[27]);
  assign t[148] = (x[27]);
  assign t[149] = (x[27]);
  assign t[14] = t[23] & t[24];
  assign t[150] = (x[32]);
  assign t[151] = (x[32]);
  assign t[152] = (x[32]);
  assign t[153] = (x[32]);
  assign t[154] = (x[37]);
  assign t[155] = (x[37]);
  assign t[156] = (x[37]);
  assign t[157] = (x[37]);
  assign t[158] = (x[42]);
  assign t[159] = (x[42]);
  assign t[15] = t[25] ^ t[26];
  assign t[160] = (x[42]);
  assign t[161] = (x[42]);
  assign t[162] = (x[47]);
  assign t[163] = (x[47]);
  assign t[164] = (x[47]);
  assign t[165] = (x[47]);
  assign t[166] = (x[52]);
  assign t[167] = (x[52]);
  assign t[168] = (x[52]);
  assign t[169] = (x[52]);
  assign t[16] = t[27] & t[28];
  assign t[170] = (x[57]);
  assign t[171] = (x[57]);
  assign t[172] = (x[57]);
  assign t[173] = (x[57]);
  assign t[174] = (x[62]);
  assign t[175] = (x[62]);
  assign t[176] = (x[62]);
  assign t[177] = (x[62]);
  assign t[17] = t[36] ^ t[37];
  assign t[18] = t[19] & t[29];
  assign t[19] = ~(t[37]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[38] ^ t[19]);
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[23] & t[30];
  assign t[23] = ~(t[40]);
  assign t[24] = ~(t[41] ^ t[23]);
  assign t[25] = t[42] ^ t[43];
  assign t[26] = t[27] & t[31];
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[44] ^ t[27]);
  assign t[29] = t[38] ^ t[32];
  assign t[2] = ~(t[4] ^ t[35]);
  assign t[30] = t[41] ^ t[33];
  assign t[31] = t[44] ^ t[34];
  assign t[32] = t[37] ^ t[45];
  assign t[33] = t[40] ^ t[46];
  assign t[34] = t[43] ^ t[47];
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = t[61] ^ x[6];
  assign t[49] = t[62] ^ x[11];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ x[16];
  assign t[51] = t[64] ^ x[21];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[31];
  assign t[54] = t[67] ^ x[36];
  assign t[55] = t[68] ^ x[41];
  assign t[56] = t[69] ^ x[46];
  assign t[57] = t[70] ^ x[51];
  assign t[58] = t[71] ^ x[56];
  assign t[59] = t[72] ^ x[61];
  assign t[5] = ~(t[8]);
  assign t[60] = t[73] ^ x[66];
  assign t[61] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[62] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[63] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[64] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[65] = (~t[90] & t[91] & t[92] & t[93]) | (t[90] & ~t[92] & ~t[93]) | (t[90] & ~t[91] & ~t[93]) | (t[90] & ~t[91] & ~t[92]);
  assign t[66] = (~t[94] & t[95] & t[96] & t[97]) | (t[94] & ~t[96] & ~t[97]) | (t[94] & ~t[95] & ~t[97]) | (t[94] & ~t[95] & ~t[96]);
  assign t[67] = (~t[98] & t[99] & t[100] & t[101]) | (t[98] & ~t[100] & ~t[101]) | (t[98] & ~t[99] & ~t[101]) | (t[98] & ~t[99] & ~t[100]);
  assign t[68] = (~t[102] & t[103] & t[104] & t[105]) | (t[102] & ~t[104] & ~t[105]) | (t[102] & ~t[103] & ~t[105]) | (t[102] & ~t[103] & ~t[104]);
  assign t[69] = (~t[106] & t[107] & t[108] & t[109]) | (t[106] & ~t[108] & ~t[109]) | (t[106] & ~t[107] & ~t[109]) | (t[106] & ~t[107] & ~t[108]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[110] & t[111] & t[112] & t[113]) | (t[110] & ~t[112] & ~t[113]) | (t[110] & ~t[111] & ~t[113]) | (t[110] & ~t[111] & ~t[112]);
  assign t[71] = (~t[114] & t[115] & t[116] & t[117]) | (t[114] & ~t[116] & ~t[117]) | (t[114] & ~t[115] & ~t[117]) | (t[114] & ~t[115] & ~t[116]);
  assign t[72] = (~t[118] & t[119] & t[120] & t[121]) | (t[118] & ~t[120] & ~t[121]) | (t[118] & ~t[119] & ~t[121]) | (t[118] & ~t[119] & ~t[120]);
  assign t[73] = (~t[122] & t[123] & t[124] & t[125]) | (t[122] & ~t[124] & ~t[125]) | (t[122] & ~t[123] & ~t[125]) | (t[122] & ~t[123] & ~t[124]);
  assign t[74] = t[126] ^ x[6];
  assign t[75] = t[127] ^ x[3];
  assign t[76] = t[128] ^ x[4];
  assign t[77] = t[129] ^ x[5];
  assign t[78] = t[130] ^ x[11];
  assign t[79] = t[131] ^ x[8];
  assign t[7] = ~(t[10]);
  assign t[80] = t[132] ^ x[9];
  assign t[81] = t[133] ^ x[10];
  assign t[82] = t[134] ^ x[16];
  assign t[83] = t[135] ^ x[13];
  assign t[84] = t[136] ^ x[14];
  assign t[85] = t[137] ^ x[15];
  assign t[86] = t[138] ^ x[21];
  assign t[87] = t[139] ^ x[18];
  assign t[88] = t[140] ^ x[19];
  assign t[89] = t[141] ^ x[20];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[142] ^ x[26];
  assign t[91] = t[143] ^ x[23];
  assign t[92] = t[144] ^ x[24];
  assign t[93] = t[145] ^ x[25];
  assign t[94] = t[146] ^ x[31];
  assign t[95] = t[147] ^ x[28];
  assign t[96] = t[148] ^ x[29];
  assign t[97] = t[149] ^ x[30];
  assign t[98] = t[150] ^ x[36];
  assign t[99] = t[151] ^ x[33];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind238(x, y);
 input [66:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[34];
  assign t[101] = t[153] ^ x[35];
  assign t[102] = t[154] ^ x[41];
  assign t[103] = t[155] ^ x[38];
  assign t[104] = t[156] ^ x[39];
  assign t[105] = t[157] ^ x[40];
  assign t[106] = t[158] ^ x[46];
  assign t[107] = t[159] ^ x[43];
  assign t[108] = t[160] ^ x[44];
  assign t[109] = t[161] ^ x[45];
  assign t[10] = t[15] ^ t[16];
  assign t[110] = t[162] ^ x[51];
  assign t[111] = t[163] ^ x[48];
  assign t[112] = t[164] ^ x[49];
  assign t[113] = t[165] ^ x[50];
  assign t[114] = t[166] ^ x[56];
  assign t[115] = t[167] ^ x[53];
  assign t[116] = t[168] ^ x[54];
  assign t[117] = t[169] ^ x[55];
  assign t[118] = t[170] ^ x[61];
  assign t[119] = t[171] ^ x[58];
  assign t[11] = t[17] ^ t[18];
  assign t[120] = t[172] ^ x[59];
  assign t[121] = t[173] ^ x[60];
  assign t[122] = t[174] ^ x[66];
  assign t[123] = t[175] ^ x[63];
  assign t[124] = t[176] ^ x[64];
  assign t[125] = t[177] ^ x[65];
  assign t[126] = (x[2]);
  assign t[127] = (x[2]);
  assign t[128] = (x[2]);
  assign t[129] = (x[2]);
  assign t[12] = t[19] & t[20];
  assign t[130] = (x[7]);
  assign t[131] = (x[7]);
  assign t[132] = (x[7]);
  assign t[133] = (x[7]);
  assign t[134] = (x[12]);
  assign t[135] = (x[12]);
  assign t[136] = (x[12]);
  assign t[137] = (x[12]);
  assign t[138] = (x[17]);
  assign t[139] = (x[17]);
  assign t[13] = t[21] ^ t[22];
  assign t[140] = (x[17]);
  assign t[141] = (x[17]);
  assign t[142] = (x[22]);
  assign t[143] = (x[22]);
  assign t[144] = (x[22]);
  assign t[145] = (x[22]);
  assign t[146] = (x[27]);
  assign t[147] = (x[27]);
  assign t[148] = (x[27]);
  assign t[149] = (x[27]);
  assign t[14] = t[23] & t[24];
  assign t[150] = (x[32]);
  assign t[151] = (x[32]);
  assign t[152] = (x[32]);
  assign t[153] = (x[32]);
  assign t[154] = (x[37]);
  assign t[155] = (x[37]);
  assign t[156] = (x[37]);
  assign t[157] = (x[37]);
  assign t[158] = (x[42]);
  assign t[159] = (x[42]);
  assign t[15] = t[25] ^ t[26];
  assign t[160] = (x[42]);
  assign t[161] = (x[42]);
  assign t[162] = (x[47]);
  assign t[163] = (x[47]);
  assign t[164] = (x[47]);
  assign t[165] = (x[47]);
  assign t[166] = (x[52]);
  assign t[167] = (x[52]);
  assign t[168] = (x[52]);
  assign t[169] = (x[52]);
  assign t[16] = t[27] & t[28];
  assign t[170] = (x[57]);
  assign t[171] = (x[57]);
  assign t[172] = (x[57]);
  assign t[173] = (x[57]);
  assign t[174] = (x[62]);
  assign t[175] = (x[62]);
  assign t[176] = (x[62]);
  assign t[177] = (x[62]);
  assign t[17] = t[36] ^ t[37];
  assign t[18] = t[19] & t[29];
  assign t[19] = ~(t[37]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[38] ^ t[19]);
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[23] & t[30];
  assign t[23] = ~(t[40]);
  assign t[24] = ~(t[41] ^ t[23]);
  assign t[25] = t[42] ^ t[43];
  assign t[26] = t[27] & t[31];
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[44] ^ t[27]);
  assign t[29] = t[38] ^ t[32];
  assign t[2] = ~(t[4] ^ t[35]);
  assign t[30] = t[41] ^ t[33];
  assign t[31] = t[44] ^ t[34];
  assign t[32] = t[37] ^ t[45];
  assign t[33] = t[40] ^ t[46];
  assign t[34] = t[43] ^ t[47];
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = t[61] ^ x[6];
  assign t[49] = t[62] ^ x[11];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ x[16];
  assign t[51] = t[64] ^ x[21];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[31];
  assign t[54] = t[67] ^ x[36];
  assign t[55] = t[68] ^ x[41];
  assign t[56] = t[69] ^ x[46];
  assign t[57] = t[70] ^ x[51];
  assign t[58] = t[71] ^ x[56];
  assign t[59] = t[72] ^ x[61];
  assign t[5] = ~(t[8]);
  assign t[60] = t[73] ^ x[66];
  assign t[61] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[62] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[63] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[64] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[65] = (~t[90] & t[91] & t[92] & t[93]) | (t[90] & ~t[92] & ~t[93]) | (t[90] & ~t[91] & ~t[93]) | (t[90] & ~t[91] & ~t[92]);
  assign t[66] = (~t[94] & t[95] & t[96] & t[97]) | (t[94] & ~t[96] & ~t[97]) | (t[94] & ~t[95] & ~t[97]) | (t[94] & ~t[95] & ~t[96]);
  assign t[67] = (~t[98] & t[99] & t[100] & t[101]) | (t[98] & ~t[100] & ~t[101]) | (t[98] & ~t[99] & ~t[101]) | (t[98] & ~t[99] & ~t[100]);
  assign t[68] = (~t[102] & t[103] & t[104] & t[105]) | (t[102] & ~t[104] & ~t[105]) | (t[102] & ~t[103] & ~t[105]) | (t[102] & ~t[103] & ~t[104]);
  assign t[69] = (~t[106] & t[107] & t[108] & t[109]) | (t[106] & ~t[108] & ~t[109]) | (t[106] & ~t[107] & ~t[109]) | (t[106] & ~t[107] & ~t[108]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[110] & t[111] & t[112] & t[113]) | (t[110] & ~t[112] & ~t[113]) | (t[110] & ~t[111] & ~t[113]) | (t[110] & ~t[111] & ~t[112]);
  assign t[71] = (~t[114] & t[115] & t[116] & t[117]) | (t[114] & ~t[116] & ~t[117]) | (t[114] & ~t[115] & ~t[117]) | (t[114] & ~t[115] & ~t[116]);
  assign t[72] = (~t[118] & t[119] & t[120] & t[121]) | (t[118] & ~t[120] & ~t[121]) | (t[118] & ~t[119] & ~t[121]) | (t[118] & ~t[119] & ~t[120]);
  assign t[73] = (~t[122] & t[123] & t[124] & t[125]) | (t[122] & ~t[124] & ~t[125]) | (t[122] & ~t[123] & ~t[125]) | (t[122] & ~t[123] & ~t[124]);
  assign t[74] = t[126] ^ x[6];
  assign t[75] = t[127] ^ x[3];
  assign t[76] = t[128] ^ x[4];
  assign t[77] = t[129] ^ x[5];
  assign t[78] = t[130] ^ x[11];
  assign t[79] = t[131] ^ x[8];
  assign t[7] = ~(t[10]);
  assign t[80] = t[132] ^ x[9];
  assign t[81] = t[133] ^ x[10];
  assign t[82] = t[134] ^ x[16];
  assign t[83] = t[135] ^ x[13];
  assign t[84] = t[136] ^ x[14];
  assign t[85] = t[137] ^ x[15];
  assign t[86] = t[138] ^ x[21];
  assign t[87] = t[139] ^ x[18];
  assign t[88] = t[140] ^ x[19];
  assign t[89] = t[141] ^ x[20];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[142] ^ x[26];
  assign t[91] = t[143] ^ x[23];
  assign t[92] = t[144] ^ x[24];
  assign t[93] = t[145] ^ x[25];
  assign t[94] = t[146] ^ x[31];
  assign t[95] = t[147] ^ x[28];
  assign t[96] = t[148] ^ x[29];
  assign t[97] = t[149] ^ x[30];
  assign t[98] = t[150] ^ x[36];
  assign t[99] = t[151] ^ x[33];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind239(x, y);
 input [66:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[34];
  assign t[101] = t[153] ^ x[35];
  assign t[102] = t[154] ^ x[41];
  assign t[103] = t[155] ^ x[38];
  assign t[104] = t[156] ^ x[39];
  assign t[105] = t[157] ^ x[40];
  assign t[106] = t[158] ^ x[46];
  assign t[107] = t[159] ^ x[43];
  assign t[108] = t[160] ^ x[44];
  assign t[109] = t[161] ^ x[45];
  assign t[10] = t[15] ^ t[16];
  assign t[110] = t[162] ^ x[51];
  assign t[111] = t[163] ^ x[48];
  assign t[112] = t[164] ^ x[49];
  assign t[113] = t[165] ^ x[50];
  assign t[114] = t[166] ^ x[56];
  assign t[115] = t[167] ^ x[53];
  assign t[116] = t[168] ^ x[54];
  assign t[117] = t[169] ^ x[55];
  assign t[118] = t[170] ^ x[61];
  assign t[119] = t[171] ^ x[58];
  assign t[11] = t[17] ^ t[18];
  assign t[120] = t[172] ^ x[59];
  assign t[121] = t[173] ^ x[60];
  assign t[122] = t[174] ^ x[66];
  assign t[123] = t[175] ^ x[63];
  assign t[124] = t[176] ^ x[64];
  assign t[125] = t[177] ^ x[65];
  assign t[126] = (x[2]);
  assign t[127] = (x[2]);
  assign t[128] = (x[2]);
  assign t[129] = (x[2]);
  assign t[12] = t[19] & t[20];
  assign t[130] = (x[7]);
  assign t[131] = (x[7]);
  assign t[132] = (x[7]);
  assign t[133] = (x[7]);
  assign t[134] = (x[12]);
  assign t[135] = (x[12]);
  assign t[136] = (x[12]);
  assign t[137] = (x[12]);
  assign t[138] = (x[17]);
  assign t[139] = (x[17]);
  assign t[13] = t[21] ^ t[22];
  assign t[140] = (x[17]);
  assign t[141] = (x[17]);
  assign t[142] = (x[22]);
  assign t[143] = (x[22]);
  assign t[144] = (x[22]);
  assign t[145] = (x[22]);
  assign t[146] = (x[27]);
  assign t[147] = (x[27]);
  assign t[148] = (x[27]);
  assign t[149] = (x[27]);
  assign t[14] = t[23] & t[24];
  assign t[150] = (x[32]);
  assign t[151] = (x[32]);
  assign t[152] = (x[32]);
  assign t[153] = (x[32]);
  assign t[154] = (x[37]);
  assign t[155] = (x[37]);
  assign t[156] = (x[37]);
  assign t[157] = (x[37]);
  assign t[158] = (x[42]);
  assign t[159] = (x[42]);
  assign t[15] = t[25] ^ t[26];
  assign t[160] = (x[42]);
  assign t[161] = (x[42]);
  assign t[162] = (x[47]);
  assign t[163] = (x[47]);
  assign t[164] = (x[47]);
  assign t[165] = (x[47]);
  assign t[166] = (x[52]);
  assign t[167] = (x[52]);
  assign t[168] = (x[52]);
  assign t[169] = (x[52]);
  assign t[16] = t[27] & t[28];
  assign t[170] = (x[57]);
  assign t[171] = (x[57]);
  assign t[172] = (x[57]);
  assign t[173] = (x[57]);
  assign t[174] = (x[62]);
  assign t[175] = (x[62]);
  assign t[176] = (x[62]);
  assign t[177] = (x[62]);
  assign t[17] = t[36] ^ t[37];
  assign t[18] = t[19] & t[29];
  assign t[19] = ~(t[37]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[38] ^ t[19]);
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[23] & t[30];
  assign t[23] = ~(t[40]);
  assign t[24] = ~(t[41] ^ t[23]);
  assign t[25] = t[42] ^ t[43];
  assign t[26] = t[27] & t[31];
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[44] ^ t[27]);
  assign t[29] = t[38] ^ t[32];
  assign t[2] = ~(t[4] ^ t[35]);
  assign t[30] = t[41] ^ t[33];
  assign t[31] = t[44] ^ t[34];
  assign t[32] = t[37] ^ t[45];
  assign t[33] = t[40] ^ t[46];
  assign t[34] = t[43] ^ t[47];
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = t[61] ^ x[6];
  assign t[49] = t[62] ^ x[11];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ x[16];
  assign t[51] = t[64] ^ x[21];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[31];
  assign t[54] = t[67] ^ x[36];
  assign t[55] = t[68] ^ x[41];
  assign t[56] = t[69] ^ x[46];
  assign t[57] = t[70] ^ x[51];
  assign t[58] = t[71] ^ x[56];
  assign t[59] = t[72] ^ x[61];
  assign t[5] = ~(t[8]);
  assign t[60] = t[73] ^ x[66];
  assign t[61] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[62] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[63] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[64] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[65] = (~t[90] & t[91] & t[92] & t[93]) | (t[90] & ~t[92] & ~t[93]) | (t[90] & ~t[91] & ~t[93]) | (t[90] & ~t[91] & ~t[92]);
  assign t[66] = (~t[94] & t[95] & t[96] & t[97]) | (t[94] & ~t[96] & ~t[97]) | (t[94] & ~t[95] & ~t[97]) | (t[94] & ~t[95] & ~t[96]);
  assign t[67] = (~t[98] & t[99] & t[100] & t[101]) | (t[98] & ~t[100] & ~t[101]) | (t[98] & ~t[99] & ~t[101]) | (t[98] & ~t[99] & ~t[100]);
  assign t[68] = (~t[102] & t[103] & t[104] & t[105]) | (t[102] & ~t[104] & ~t[105]) | (t[102] & ~t[103] & ~t[105]) | (t[102] & ~t[103] & ~t[104]);
  assign t[69] = (~t[106] & t[107] & t[108] & t[109]) | (t[106] & ~t[108] & ~t[109]) | (t[106] & ~t[107] & ~t[109]) | (t[106] & ~t[107] & ~t[108]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[110] & t[111] & t[112] & t[113]) | (t[110] & ~t[112] & ~t[113]) | (t[110] & ~t[111] & ~t[113]) | (t[110] & ~t[111] & ~t[112]);
  assign t[71] = (~t[114] & t[115] & t[116] & t[117]) | (t[114] & ~t[116] & ~t[117]) | (t[114] & ~t[115] & ~t[117]) | (t[114] & ~t[115] & ~t[116]);
  assign t[72] = (~t[118] & t[119] & t[120] & t[121]) | (t[118] & ~t[120] & ~t[121]) | (t[118] & ~t[119] & ~t[121]) | (t[118] & ~t[119] & ~t[120]);
  assign t[73] = (~t[122] & t[123] & t[124] & t[125]) | (t[122] & ~t[124] & ~t[125]) | (t[122] & ~t[123] & ~t[125]) | (t[122] & ~t[123] & ~t[124]);
  assign t[74] = t[126] ^ x[6];
  assign t[75] = t[127] ^ x[3];
  assign t[76] = t[128] ^ x[4];
  assign t[77] = t[129] ^ x[5];
  assign t[78] = t[130] ^ x[11];
  assign t[79] = t[131] ^ x[8];
  assign t[7] = ~(t[10]);
  assign t[80] = t[132] ^ x[9];
  assign t[81] = t[133] ^ x[10];
  assign t[82] = t[134] ^ x[16];
  assign t[83] = t[135] ^ x[13];
  assign t[84] = t[136] ^ x[14];
  assign t[85] = t[137] ^ x[15];
  assign t[86] = t[138] ^ x[21];
  assign t[87] = t[139] ^ x[18];
  assign t[88] = t[140] ^ x[19];
  assign t[89] = t[141] ^ x[20];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[142] ^ x[26];
  assign t[91] = t[143] ^ x[23];
  assign t[92] = t[144] ^ x[24];
  assign t[93] = t[145] ^ x[25];
  assign t[94] = t[146] ^ x[31];
  assign t[95] = t[147] ^ x[28];
  assign t[96] = t[148] ^ x[29];
  assign t[97] = t[149] ^ x[30];
  assign t[98] = t[150] ^ x[36];
  assign t[99] = t[151] ^ x[33];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind240(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[54] & t[26];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[55] & t[31];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[56] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[54] ^ t[27]);
  assign t[29] = t[58] ^ t[57];
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[55] ^ t[32]);
  assign t[34] = t[60] ^ t[59];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[56] ^ t[37]);
  assign t[39] = t[62] ^ t[61];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[54] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[54] ^ t[50];
  assign t[44] = t[55] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[55] ^ t[51];
  assign t[47] = t[56] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[56] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[57] ^ t[63];
  assign t[51] = t[59] ^ t[64];
  assign t[52] = t[61] ^ t[65];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] & t[17];
  assign y = (t[0]);
endmodule

module R2ind241(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[54] & t[26];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[55] & t[31];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[56] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[54] ^ t[27]);
  assign t[29] = t[58] ^ t[57];
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[55] ^ t[32]);
  assign t[34] = t[60] ^ t[59];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[56] ^ t[37]);
  assign t[39] = t[62] ^ t[61];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[54] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[54] ^ t[50];
  assign t[44] = t[55] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[55] ^ t[51];
  assign t[47] = t[56] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[56] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[57] ^ t[63];
  assign t[51] = t[59] ^ t[64];
  assign t[52] = t[61] ^ t[65];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] & t[17];
  assign y = (t[0]);
endmodule

module R2ind242(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[54] & t[26];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[55] & t[31];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[56] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[54] ^ t[27]);
  assign t[29] = t[58] ^ t[57];
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[55] ^ t[32]);
  assign t[34] = t[60] ^ t[59];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[56] ^ t[37]);
  assign t[39] = t[62] ^ t[61];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[54] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[54] ^ t[50];
  assign t[44] = t[55] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[55] ^ t[51];
  assign t[47] = t[56] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[56] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[57] ^ t[63];
  assign t[51] = t[59] ^ t[64];
  assign t[52] = t[61] ^ t[65];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] & t[17];
  assign y = (t[0]);
endmodule

module R2ind243(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[54] & t[26];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[55] & t[31];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[56] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[54] ^ t[27]);
  assign t[29] = t[58] ^ t[57];
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[55] ^ t[32]);
  assign t[34] = t[60] ^ t[59];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[56] ^ t[37]);
  assign t[39] = t[62] ^ t[61];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[54] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[54] ^ t[50];
  assign t[44] = t[55] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[55] ^ t[51];
  assign t[47] = t[56] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[56] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[57] ^ t[63];
  assign t[51] = t[59] ^ t[64];
  assign t[52] = t[61] ^ t[65];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] & t[17];
  assign y = (t[0]);
endmodule

module R2ind244(x, y);
 input [66:0] x;
 output y;

 wire [196:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[10];
  assign t[101] = t[153] ^ x[16];
  assign t[102] = t[154] ^ x[13];
  assign t[103] = t[155] ^ x[14];
  assign t[104] = t[156] ^ x[15];
  assign t[105] = t[157] ^ x[21];
  assign t[106] = t[158] ^ x[18];
  assign t[107] = t[159] ^ x[19];
  assign t[108] = t[160] ^ x[20];
  assign t[109] = t[161] ^ x[26];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[162] ^ x[23];
  assign t[111] = t[163] ^ x[24];
  assign t[112] = t[164] ^ x[25];
  assign t[113] = t[165] ^ x[31];
  assign t[114] = t[166] ^ x[28];
  assign t[115] = t[167] ^ x[29];
  assign t[116] = t[168] ^ x[30];
  assign t[117] = t[169] ^ x[36];
  assign t[118] = t[170] ^ x[33];
  assign t[119] = t[171] ^ x[34];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[172] ^ x[35];
  assign t[121] = t[173] ^ x[41];
  assign t[122] = t[174] ^ x[38];
  assign t[123] = t[175] ^ x[39];
  assign t[124] = t[176] ^ x[40];
  assign t[125] = t[177] ^ x[46];
  assign t[126] = t[178] ^ x[43];
  assign t[127] = t[179] ^ x[44];
  assign t[128] = t[180] ^ x[45];
  assign t[129] = t[181] ^ x[51];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[182] ^ x[48];
  assign t[131] = t[183] ^ x[49];
  assign t[132] = t[184] ^ x[50];
  assign t[133] = t[185] ^ x[56];
  assign t[134] = t[186] ^ x[53];
  assign t[135] = t[187] ^ x[54];
  assign t[136] = t[188] ^ x[55];
  assign t[137] = t[189] ^ x[61];
  assign t[138] = t[190] ^ x[58];
  assign t[139] = t[191] ^ x[59];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[192] ^ x[60];
  assign t[141] = t[193] ^ x[66];
  assign t[142] = t[194] ^ x[63];
  assign t[143] = t[195] ^ x[64];
  assign t[144] = t[196] ^ x[65];
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[2]);
  assign t[149] = (x[7]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[7]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[12]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[27] ^ t[28];
  assign t[160] = (x[17]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[22]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[27]);
  assign t[169] = (x[32]);
  assign t[16] = t[29] & t[30];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[32]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[37]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[31] ^ t[16];
  assign t[180] = (x[42]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[47]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[52]);
  assign t[189] = (x[57]);
  assign t[18] = t[55] ^ t[29];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[57]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[196] = (x[62]);
  assign t[19] = t[32] ^ t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] & t[35];
  assign t[21] = t[36] ^ t[20];
  assign t[22] = t[56] ^ t[34];
  assign t[23] = t[37] ^ t[38];
  assign t[24] = t[39] & t[40];
  assign t[25] = t[41] ^ t[24];
  assign t[26] = t[57] ^ t[39];
  assign t[27] = t[58] ^ t[59];
  assign t[28] = t[29] & t[42];
  assign t[29] = ~(t[59]);
  assign t[2] = ~(t[4] ^ t[54]);
  assign t[30] = ~(t[55] ^ t[29]);
  assign t[31] = t[55] & t[43];
  assign t[32] = t[60] ^ t[61];
  assign t[33] = t[34] & t[44];
  assign t[34] = ~(t[61]);
  assign t[35] = ~(t[56] ^ t[34]);
  assign t[36] = t[56] & t[45];
  assign t[37] = t[62] ^ t[63];
  assign t[38] = t[39] & t[46];
  assign t[39] = ~(t[63]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[57] ^ t[39]);
  assign t[41] = t[57] & t[47];
  assign t[42] = t[55] ^ t[48];
  assign t[43] = t[49] ^ t[28];
  assign t[44] = t[56] ^ t[50];
  assign t[45] = t[51] ^ t[33];
  assign t[46] = t[57] ^ t[52];
  assign t[47] = t[53] ^ t[38];
  assign t[48] = t[59] ^ t[64];
  assign t[49] = t[55] ^ t[27];
  assign t[4] = ~t[7];
  assign t[50] = t[61] ^ t[65];
  assign t[51] = t[56] ^ t[32];
  assign t[52] = t[63] ^ t[66];
  assign t[53] = t[57] ^ t[37];
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = ~(t[8]);
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = (t[79]);
  assign t[67] = t[80] ^ x[6];
  assign t[68] = t[81] ^ x[11];
  assign t[69] = t[82] ^ x[16];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[83] ^ x[21];
  assign t[71] = t[84] ^ x[26];
  assign t[72] = t[85] ^ x[31];
  assign t[73] = t[86] ^ x[36];
  assign t[74] = t[87] ^ x[41];
  assign t[75] = t[88] ^ x[46];
  assign t[76] = t[89] ^ x[51];
  assign t[77] = t[90] ^ x[56];
  assign t[78] = t[91] ^ x[61];
  assign t[79] = t[92] ^ x[66];
  assign t[7] = ~(t[11] ^ t[12]);
  assign t[80] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[81] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[82] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[83] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[84] = (~t[109] & t[110] & t[111] & t[112]) | (t[109] & ~t[111] & ~t[112]) | (t[109] & ~t[110] & ~t[112]) | (t[109] & ~t[110] & ~t[111]);
  assign t[85] = (~t[113] & t[114] & t[115] & t[116]) | (t[113] & ~t[115] & ~t[116]) | (t[113] & ~t[114] & ~t[116]) | (t[113] & ~t[114] & ~t[115]);
  assign t[86] = (~t[117] & t[118] & t[119] & t[120]) | (t[117] & ~t[119] & ~t[120]) | (t[117] & ~t[118] & ~t[120]) | (t[117] & ~t[118] & ~t[119]);
  assign t[87] = (~t[121] & t[122] & t[123] & t[124]) | (t[121] & ~t[123] & ~t[124]) | (t[121] & ~t[122] & ~t[124]) | (t[121] & ~t[122] & ~t[123]);
  assign t[88] = (~t[125] & t[126] & t[127] & t[128]) | (t[125] & ~t[127] & ~t[128]) | (t[125] & ~t[126] & ~t[128]) | (t[125] & ~t[126] & ~t[127]);
  assign t[89] = (~t[129] & t[130] & t[131] & t[132]) | (t[129] & ~t[131] & ~t[132]) | (t[129] & ~t[130] & ~t[132]) | (t[129] & ~t[130] & ~t[131]);
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = (~t[133] & t[134] & t[135] & t[136]) | (t[133] & ~t[135] & ~t[136]) | (t[133] & ~t[134] & ~t[136]) | (t[133] & ~t[134] & ~t[135]);
  assign t[91] = (~t[137] & t[138] & t[139] & t[140]) | (t[137] & ~t[139] & ~t[140]) | (t[137] & ~t[138] & ~t[140]) | (t[137] & ~t[138] & ~t[139]);
  assign t[92] = (~t[141] & t[142] & t[143] & t[144]) | (t[141] & ~t[143] & ~t[144]) | (t[141] & ~t[142] & ~t[144]) | (t[141] & ~t[142] & ~t[143]);
  assign t[93] = t[145] ^ x[6];
  assign t[94] = t[146] ^ x[3];
  assign t[95] = t[147] ^ x[4];
  assign t[96] = t[148] ^ x[5];
  assign t[97] = t[149] ^ x[11];
  assign t[98] = t[150] ^ x[8];
  assign t[99] = t[151] ^ x[9];
  assign t[9] = t[15] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind245(x, y);
 input [66:0] x;
 output y;

 wire [196:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[10];
  assign t[101] = t[153] ^ x[16];
  assign t[102] = t[154] ^ x[13];
  assign t[103] = t[155] ^ x[14];
  assign t[104] = t[156] ^ x[15];
  assign t[105] = t[157] ^ x[21];
  assign t[106] = t[158] ^ x[18];
  assign t[107] = t[159] ^ x[19];
  assign t[108] = t[160] ^ x[20];
  assign t[109] = t[161] ^ x[26];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[162] ^ x[23];
  assign t[111] = t[163] ^ x[24];
  assign t[112] = t[164] ^ x[25];
  assign t[113] = t[165] ^ x[31];
  assign t[114] = t[166] ^ x[28];
  assign t[115] = t[167] ^ x[29];
  assign t[116] = t[168] ^ x[30];
  assign t[117] = t[169] ^ x[36];
  assign t[118] = t[170] ^ x[33];
  assign t[119] = t[171] ^ x[34];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[172] ^ x[35];
  assign t[121] = t[173] ^ x[41];
  assign t[122] = t[174] ^ x[38];
  assign t[123] = t[175] ^ x[39];
  assign t[124] = t[176] ^ x[40];
  assign t[125] = t[177] ^ x[46];
  assign t[126] = t[178] ^ x[43];
  assign t[127] = t[179] ^ x[44];
  assign t[128] = t[180] ^ x[45];
  assign t[129] = t[181] ^ x[51];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[182] ^ x[48];
  assign t[131] = t[183] ^ x[49];
  assign t[132] = t[184] ^ x[50];
  assign t[133] = t[185] ^ x[56];
  assign t[134] = t[186] ^ x[53];
  assign t[135] = t[187] ^ x[54];
  assign t[136] = t[188] ^ x[55];
  assign t[137] = t[189] ^ x[61];
  assign t[138] = t[190] ^ x[58];
  assign t[139] = t[191] ^ x[59];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[192] ^ x[60];
  assign t[141] = t[193] ^ x[66];
  assign t[142] = t[194] ^ x[63];
  assign t[143] = t[195] ^ x[64];
  assign t[144] = t[196] ^ x[65];
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[2]);
  assign t[149] = (x[7]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[7]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[12]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[27] ^ t[28];
  assign t[160] = (x[17]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[22]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[27]);
  assign t[169] = (x[32]);
  assign t[16] = t[29] & t[30];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[32]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[37]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[31] ^ t[16];
  assign t[180] = (x[42]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[47]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[52]);
  assign t[189] = (x[57]);
  assign t[18] = t[55] ^ t[29];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[57]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[196] = (x[62]);
  assign t[19] = t[32] ^ t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] & t[35];
  assign t[21] = t[36] ^ t[20];
  assign t[22] = t[56] ^ t[34];
  assign t[23] = t[37] ^ t[38];
  assign t[24] = t[39] & t[40];
  assign t[25] = t[41] ^ t[24];
  assign t[26] = t[57] ^ t[39];
  assign t[27] = t[58] ^ t[59];
  assign t[28] = t[29] & t[42];
  assign t[29] = ~(t[59]);
  assign t[2] = ~(t[4] ^ t[54]);
  assign t[30] = ~(t[55] ^ t[29]);
  assign t[31] = t[55] & t[43];
  assign t[32] = t[60] ^ t[61];
  assign t[33] = t[34] & t[44];
  assign t[34] = ~(t[61]);
  assign t[35] = ~(t[56] ^ t[34]);
  assign t[36] = t[56] & t[45];
  assign t[37] = t[62] ^ t[63];
  assign t[38] = t[39] & t[46];
  assign t[39] = ~(t[63]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[57] ^ t[39]);
  assign t[41] = t[57] & t[47];
  assign t[42] = t[55] ^ t[48];
  assign t[43] = t[49] ^ t[28];
  assign t[44] = t[56] ^ t[50];
  assign t[45] = t[51] ^ t[33];
  assign t[46] = t[57] ^ t[52];
  assign t[47] = t[53] ^ t[38];
  assign t[48] = t[59] ^ t[64];
  assign t[49] = t[55] ^ t[27];
  assign t[4] = ~t[7];
  assign t[50] = t[61] ^ t[65];
  assign t[51] = t[56] ^ t[32];
  assign t[52] = t[63] ^ t[66];
  assign t[53] = t[57] ^ t[37];
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = ~(t[8]);
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = (t[79]);
  assign t[67] = t[80] ^ x[6];
  assign t[68] = t[81] ^ x[11];
  assign t[69] = t[82] ^ x[16];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[83] ^ x[21];
  assign t[71] = t[84] ^ x[26];
  assign t[72] = t[85] ^ x[31];
  assign t[73] = t[86] ^ x[36];
  assign t[74] = t[87] ^ x[41];
  assign t[75] = t[88] ^ x[46];
  assign t[76] = t[89] ^ x[51];
  assign t[77] = t[90] ^ x[56];
  assign t[78] = t[91] ^ x[61];
  assign t[79] = t[92] ^ x[66];
  assign t[7] = ~(t[11] ^ t[12]);
  assign t[80] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[81] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[82] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[83] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[84] = (~t[109] & t[110] & t[111] & t[112]) | (t[109] & ~t[111] & ~t[112]) | (t[109] & ~t[110] & ~t[112]) | (t[109] & ~t[110] & ~t[111]);
  assign t[85] = (~t[113] & t[114] & t[115] & t[116]) | (t[113] & ~t[115] & ~t[116]) | (t[113] & ~t[114] & ~t[116]) | (t[113] & ~t[114] & ~t[115]);
  assign t[86] = (~t[117] & t[118] & t[119] & t[120]) | (t[117] & ~t[119] & ~t[120]) | (t[117] & ~t[118] & ~t[120]) | (t[117] & ~t[118] & ~t[119]);
  assign t[87] = (~t[121] & t[122] & t[123] & t[124]) | (t[121] & ~t[123] & ~t[124]) | (t[121] & ~t[122] & ~t[124]) | (t[121] & ~t[122] & ~t[123]);
  assign t[88] = (~t[125] & t[126] & t[127] & t[128]) | (t[125] & ~t[127] & ~t[128]) | (t[125] & ~t[126] & ~t[128]) | (t[125] & ~t[126] & ~t[127]);
  assign t[89] = (~t[129] & t[130] & t[131] & t[132]) | (t[129] & ~t[131] & ~t[132]) | (t[129] & ~t[130] & ~t[132]) | (t[129] & ~t[130] & ~t[131]);
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = (~t[133] & t[134] & t[135] & t[136]) | (t[133] & ~t[135] & ~t[136]) | (t[133] & ~t[134] & ~t[136]) | (t[133] & ~t[134] & ~t[135]);
  assign t[91] = (~t[137] & t[138] & t[139] & t[140]) | (t[137] & ~t[139] & ~t[140]) | (t[137] & ~t[138] & ~t[140]) | (t[137] & ~t[138] & ~t[139]);
  assign t[92] = (~t[141] & t[142] & t[143] & t[144]) | (t[141] & ~t[143] & ~t[144]) | (t[141] & ~t[142] & ~t[144]) | (t[141] & ~t[142] & ~t[143]);
  assign t[93] = t[145] ^ x[6];
  assign t[94] = t[146] ^ x[3];
  assign t[95] = t[147] ^ x[4];
  assign t[96] = t[148] ^ x[5];
  assign t[97] = t[149] ^ x[11];
  assign t[98] = t[150] ^ x[8];
  assign t[99] = t[151] ^ x[9];
  assign t[9] = t[15] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind246(x, y);
 input [66:0] x;
 output y;

 wire [196:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[10];
  assign t[101] = t[153] ^ x[16];
  assign t[102] = t[154] ^ x[13];
  assign t[103] = t[155] ^ x[14];
  assign t[104] = t[156] ^ x[15];
  assign t[105] = t[157] ^ x[21];
  assign t[106] = t[158] ^ x[18];
  assign t[107] = t[159] ^ x[19];
  assign t[108] = t[160] ^ x[20];
  assign t[109] = t[161] ^ x[26];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[162] ^ x[23];
  assign t[111] = t[163] ^ x[24];
  assign t[112] = t[164] ^ x[25];
  assign t[113] = t[165] ^ x[31];
  assign t[114] = t[166] ^ x[28];
  assign t[115] = t[167] ^ x[29];
  assign t[116] = t[168] ^ x[30];
  assign t[117] = t[169] ^ x[36];
  assign t[118] = t[170] ^ x[33];
  assign t[119] = t[171] ^ x[34];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[172] ^ x[35];
  assign t[121] = t[173] ^ x[41];
  assign t[122] = t[174] ^ x[38];
  assign t[123] = t[175] ^ x[39];
  assign t[124] = t[176] ^ x[40];
  assign t[125] = t[177] ^ x[46];
  assign t[126] = t[178] ^ x[43];
  assign t[127] = t[179] ^ x[44];
  assign t[128] = t[180] ^ x[45];
  assign t[129] = t[181] ^ x[51];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[182] ^ x[48];
  assign t[131] = t[183] ^ x[49];
  assign t[132] = t[184] ^ x[50];
  assign t[133] = t[185] ^ x[56];
  assign t[134] = t[186] ^ x[53];
  assign t[135] = t[187] ^ x[54];
  assign t[136] = t[188] ^ x[55];
  assign t[137] = t[189] ^ x[61];
  assign t[138] = t[190] ^ x[58];
  assign t[139] = t[191] ^ x[59];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[192] ^ x[60];
  assign t[141] = t[193] ^ x[66];
  assign t[142] = t[194] ^ x[63];
  assign t[143] = t[195] ^ x[64];
  assign t[144] = t[196] ^ x[65];
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[2]);
  assign t[149] = (x[7]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[7]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[12]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[27] ^ t[28];
  assign t[160] = (x[17]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[22]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[27]);
  assign t[169] = (x[32]);
  assign t[16] = t[29] & t[30];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[32]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[37]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[31] ^ t[16];
  assign t[180] = (x[42]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[47]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[52]);
  assign t[189] = (x[57]);
  assign t[18] = t[55] ^ t[29];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[57]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[196] = (x[62]);
  assign t[19] = t[32] ^ t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] & t[35];
  assign t[21] = t[36] ^ t[20];
  assign t[22] = t[56] ^ t[34];
  assign t[23] = t[37] ^ t[38];
  assign t[24] = t[39] & t[40];
  assign t[25] = t[41] ^ t[24];
  assign t[26] = t[57] ^ t[39];
  assign t[27] = t[58] ^ t[59];
  assign t[28] = t[29] & t[42];
  assign t[29] = ~(t[59]);
  assign t[2] = ~(t[4] ^ t[54]);
  assign t[30] = ~(t[55] ^ t[29]);
  assign t[31] = t[55] & t[43];
  assign t[32] = t[60] ^ t[61];
  assign t[33] = t[34] & t[44];
  assign t[34] = ~(t[61]);
  assign t[35] = ~(t[56] ^ t[34]);
  assign t[36] = t[56] & t[45];
  assign t[37] = t[62] ^ t[63];
  assign t[38] = t[39] & t[46];
  assign t[39] = ~(t[63]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[57] ^ t[39]);
  assign t[41] = t[57] & t[47];
  assign t[42] = t[55] ^ t[48];
  assign t[43] = t[49] ^ t[28];
  assign t[44] = t[56] ^ t[50];
  assign t[45] = t[51] ^ t[33];
  assign t[46] = t[57] ^ t[52];
  assign t[47] = t[53] ^ t[38];
  assign t[48] = t[59] ^ t[64];
  assign t[49] = t[55] ^ t[27];
  assign t[4] = ~t[7];
  assign t[50] = t[61] ^ t[65];
  assign t[51] = t[56] ^ t[32];
  assign t[52] = t[63] ^ t[66];
  assign t[53] = t[57] ^ t[37];
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = ~(t[8]);
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = (t[79]);
  assign t[67] = t[80] ^ x[6];
  assign t[68] = t[81] ^ x[11];
  assign t[69] = t[82] ^ x[16];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[83] ^ x[21];
  assign t[71] = t[84] ^ x[26];
  assign t[72] = t[85] ^ x[31];
  assign t[73] = t[86] ^ x[36];
  assign t[74] = t[87] ^ x[41];
  assign t[75] = t[88] ^ x[46];
  assign t[76] = t[89] ^ x[51];
  assign t[77] = t[90] ^ x[56];
  assign t[78] = t[91] ^ x[61];
  assign t[79] = t[92] ^ x[66];
  assign t[7] = ~(t[11] ^ t[12]);
  assign t[80] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[81] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[82] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[83] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[84] = (~t[109] & t[110] & t[111] & t[112]) | (t[109] & ~t[111] & ~t[112]) | (t[109] & ~t[110] & ~t[112]) | (t[109] & ~t[110] & ~t[111]);
  assign t[85] = (~t[113] & t[114] & t[115] & t[116]) | (t[113] & ~t[115] & ~t[116]) | (t[113] & ~t[114] & ~t[116]) | (t[113] & ~t[114] & ~t[115]);
  assign t[86] = (~t[117] & t[118] & t[119] & t[120]) | (t[117] & ~t[119] & ~t[120]) | (t[117] & ~t[118] & ~t[120]) | (t[117] & ~t[118] & ~t[119]);
  assign t[87] = (~t[121] & t[122] & t[123] & t[124]) | (t[121] & ~t[123] & ~t[124]) | (t[121] & ~t[122] & ~t[124]) | (t[121] & ~t[122] & ~t[123]);
  assign t[88] = (~t[125] & t[126] & t[127] & t[128]) | (t[125] & ~t[127] & ~t[128]) | (t[125] & ~t[126] & ~t[128]) | (t[125] & ~t[126] & ~t[127]);
  assign t[89] = (~t[129] & t[130] & t[131] & t[132]) | (t[129] & ~t[131] & ~t[132]) | (t[129] & ~t[130] & ~t[132]) | (t[129] & ~t[130] & ~t[131]);
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = (~t[133] & t[134] & t[135] & t[136]) | (t[133] & ~t[135] & ~t[136]) | (t[133] & ~t[134] & ~t[136]) | (t[133] & ~t[134] & ~t[135]);
  assign t[91] = (~t[137] & t[138] & t[139] & t[140]) | (t[137] & ~t[139] & ~t[140]) | (t[137] & ~t[138] & ~t[140]) | (t[137] & ~t[138] & ~t[139]);
  assign t[92] = (~t[141] & t[142] & t[143] & t[144]) | (t[141] & ~t[143] & ~t[144]) | (t[141] & ~t[142] & ~t[144]) | (t[141] & ~t[142] & ~t[143]);
  assign t[93] = t[145] ^ x[6];
  assign t[94] = t[146] ^ x[3];
  assign t[95] = t[147] ^ x[4];
  assign t[96] = t[148] ^ x[5];
  assign t[97] = t[149] ^ x[11];
  assign t[98] = t[150] ^ x[8];
  assign t[99] = t[151] ^ x[9];
  assign t[9] = t[15] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind247(x, y);
 input [66:0] x;
 output y;

 wire [196:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[10];
  assign t[101] = t[153] ^ x[16];
  assign t[102] = t[154] ^ x[13];
  assign t[103] = t[155] ^ x[14];
  assign t[104] = t[156] ^ x[15];
  assign t[105] = t[157] ^ x[21];
  assign t[106] = t[158] ^ x[18];
  assign t[107] = t[159] ^ x[19];
  assign t[108] = t[160] ^ x[20];
  assign t[109] = t[161] ^ x[26];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[162] ^ x[23];
  assign t[111] = t[163] ^ x[24];
  assign t[112] = t[164] ^ x[25];
  assign t[113] = t[165] ^ x[31];
  assign t[114] = t[166] ^ x[28];
  assign t[115] = t[167] ^ x[29];
  assign t[116] = t[168] ^ x[30];
  assign t[117] = t[169] ^ x[36];
  assign t[118] = t[170] ^ x[33];
  assign t[119] = t[171] ^ x[34];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[172] ^ x[35];
  assign t[121] = t[173] ^ x[41];
  assign t[122] = t[174] ^ x[38];
  assign t[123] = t[175] ^ x[39];
  assign t[124] = t[176] ^ x[40];
  assign t[125] = t[177] ^ x[46];
  assign t[126] = t[178] ^ x[43];
  assign t[127] = t[179] ^ x[44];
  assign t[128] = t[180] ^ x[45];
  assign t[129] = t[181] ^ x[51];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[182] ^ x[48];
  assign t[131] = t[183] ^ x[49];
  assign t[132] = t[184] ^ x[50];
  assign t[133] = t[185] ^ x[56];
  assign t[134] = t[186] ^ x[53];
  assign t[135] = t[187] ^ x[54];
  assign t[136] = t[188] ^ x[55];
  assign t[137] = t[189] ^ x[61];
  assign t[138] = t[190] ^ x[58];
  assign t[139] = t[191] ^ x[59];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[192] ^ x[60];
  assign t[141] = t[193] ^ x[66];
  assign t[142] = t[194] ^ x[63];
  assign t[143] = t[195] ^ x[64];
  assign t[144] = t[196] ^ x[65];
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[2]);
  assign t[149] = (x[7]);
  assign t[14] = t[25] ^ t[26];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[7]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[12]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[27] ^ t[28];
  assign t[160] = (x[17]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[22]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[27]);
  assign t[169] = (x[32]);
  assign t[16] = t[29] & t[30];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[32]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[37]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[31] ^ t[16];
  assign t[180] = (x[42]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[47]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[52]);
  assign t[189] = (x[57]);
  assign t[18] = t[55] ^ t[29];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[57]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[196] = (x[62]);
  assign t[19] = t[32] ^ t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] & t[35];
  assign t[21] = t[36] ^ t[20];
  assign t[22] = t[56] ^ t[34];
  assign t[23] = t[37] ^ t[38];
  assign t[24] = t[39] & t[40];
  assign t[25] = t[41] ^ t[24];
  assign t[26] = t[57] ^ t[39];
  assign t[27] = t[58] ^ t[59];
  assign t[28] = t[29] & t[42];
  assign t[29] = ~(t[59]);
  assign t[2] = ~(t[4] ^ t[54]);
  assign t[30] = ~(t[55] ^ t[29]);
  assign t[31] = t[55] & t[43];
  assign t[32] = t[60] ^ t[61];
  assign t[33] = t[34] & t[44];
  assign t[34] = ~(t[61]);
  assign t[35] = ~(t[56] ^ t[34]);
  assign t[36] = t[56] & t[45];
  assign t[37] = t[62] ^ t[63];
  assign t[38] = t[39] & t[46];
  assign t[39] = ~(t[63]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[57] ^ t[39]);
  assign t[41] = t[57] & t[47];
  assign t[42] = t[55] ^ t[48];
  assign t[43] = t[49] ^ t[28];
  assign t[44] = t[56] ^ t[50];
  assign t[45] = t[51] ^ t[33];
  assign t[46] = t[57] ^ t[52];
  assign t[47] = t[53] ^ t[38];
  assign t[48] = t[59] ^ t[64];
  assign t[49] = t[55] ^ t[27];
  assign t[4] = ~t[7];
  assign t[50] = t[61] ^ t[65];
  assign t[51] = t[56] ^ t[32];
  assign t[52] = t[63] ^ t[66];
  assign t[53] = t[57] ^ t[37];
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = ~(t[8]);
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = (t[79]);
  assign t[67] = t[80] ^ x[6];
  assign t[68] = t[81] ^ x[11];
  assign t[69] = t[82] ^ x[16];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[83] ^ x[21];
  assign t[71] = t[84] ^ x[26];
  assign t[72] = t[85] ^ x[31];
  assign t[73] = t[86] ^ x[36];
  assign t[74] = t[87] ^ x[41];
  assign t[75] = t[88] ^ x[46];
  assign t[76] = t[89] ^ x[51];
  assign t[77] = t[90] ^ x[56];
  assign t[78] = t[91] ^ x[61];
  assign t[79] = t[92] ^ x[66];
  assign t[7] = ~(t[11] ^ t[12]);
  assign t[80] = (~t[93] & t[94] & t[95] & t[96]) | (t[93] & ~t[95] & ~t[96]) | (t[93] & ~t[94] & ~t[96]) | (t[93] & ~t[94] & ~t[95]);
  assign t[81] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[82] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[83] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[84] = (~t[109] & t[110] & t[111] & t[112]) | (t[109] & ~t[111] & ~t[112]) | (t[109] & ~t[110] & ~t[112]) | (t[109] & ~t[110] & ~t[111]);
  assign t[85] = (~t[113] & t[114] & t[115] & t[116]) | (t[113] & ~t[115] & ~t[116]) | (t[113] & ~t[114] & ~t[116]) | (t[113] & ~t[114] & ~t[115]);
  assign t[86] = (~t[117] & t[118] & t[119] & t[120]) | (t[117] & ~t[119] & ~t[120]) | (t[117] & ~t[118] & ~t[120]) | (t[117] & ~t[118] & ~t[119]);
  assign t[87] = (~t[121] & t[122] & t[123] & t[124]) | (t[121] & ~t[123] & ~t[124]) | (t[121] & ~t[122] & ~t[124]) | (t[121] & ~t[122] & ~t[123]);
  assign t[88] = (~t[125] & t[126] & t[127] & t[128]) | (t[125] & ~t[127] & ~t[128]) | (t[125] & ~t[126] & ~t[128]) | (t[125] & ~t[126] & ~t[127]);
  assign t[89] = (~t[129] & t[130] & t[131] & t[132]) | (t[129] & ~t[131] & ~t[132]) | (t[129] & ~t[130] & ~t[132]) | (t[129] & ~t[130] & ~t[131]);
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = (~t[133] & t[134] & t[135] & t[136]) | (t[133] & ~t[135] & ~t[136]) | (t[133] & ~t[134] & ~t[136]) | (t[133] & ~t[134] & ~t[135]);
  assign t[91] = (~t[137] & t[138] & t[139] & t[140]) | (t[137] & ~t[139] & ~t[140]) | (t[137] & ~t[138] & ~t[140]) | (t[137] & ~t[138] & ~t[139]);
  assign t[92] = (~t[141] & t[142] & t[143] & t[144]) | (t[141] & ~t[143] & ~t[144]) | (t[141] & ~t[142] & ~t[144]) | (t[141] & ~t[142] & ~t[143]);
  assign t[93] = t[145] ^ x[6];
  assign t[94] = t[146] ^ x[3];
  assign t[95] = t[147] ^ x[4];
  assign t[96] = t[148] ^ x[5];
  assign t[97] = t[149] ^ x[11];
  assign t[98] = t[150] ^ x[8];
  assign t[99] = t[151] ^ x[9];
  assign t[9] = t[15] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind248(x, y);
 input [51:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[7]);
  assign t[101] = (x[12]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[17]);
  assign t[106] = (x[17]);
  assign t[107] = (x[17]);
  assign t[108] = (x[17]);
  assign t[109] = (x[22]);
  assign t[10] = t[15] ^ t[16];
  assign t[110] = (x[22]);
  assign t[111] = (x[22]);
  assign t[112] = (x[22]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[32]);
  assign t[118] = (x[32]);
  assign t[119] = (x[32]);
  assign t[11] = t[24] ^ t[25];
  assign t[120] = (x[32]);
  assign t[121] = (x[37]);
  assign t[122] = (x[37]);
  assign t[123] = (x[37]);
  assign t[124] = (x[37]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[127] = (x[42]);
  assign t[128] = (x[42]);
  assign t[129] = (x[47]);
  assign t[12] = t[17] & t[18];
  assign t[130] = (x[47]);
  assign t[131] = (x[47]);
  assign t[132] = (x[47]);
  assign t[13] = t[26] ^ t[27];
  assign t[14] = t[19] & t[20];
  assign t[15] = t[28] ^ t[29];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[30] ^ t[17]);
  assign t[19] = ~(t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] ^ t[19]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[23]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = t[43] ^ x[6];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[21];
  assign t[37] = t[47] ^ x[26];
  assign t[38] = t[48] ^ x[31];
  assign t[39] = t[49] ^ x[36];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[41];
  assign t[41] = t[51] ^ x[46];
  assign t[42] = t[52] ^ x[51];
  assign t[43] = (~t[53] & t[54] & t[55] & t[56]) | (t[53] & ~t[55] & ~t[56]) | (t[53] & ~t[54] & ~t[56]) | (t[53] & ~t[54] & ~t[55]);
  assign t[44] = (~t[57] & t[58] & t[59] & t[60]) | (t[57] & ~t[59] & ~t[60]) | (t[57] & ~t[58] & ~t[60]) | (t[57] & ~t[58] & ~t[59]);
  assign t[45] = (~t[61] & t[62] & t[63] & t[64]) | (t[61] & ~t[63] & ~t[64]) | (t[61] & ~t[62] & ~t[64]) | (t[61] & ~t[62] & ~t[63]);
  assign t[46] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[47] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[48] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[49] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[51] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[52] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[53] = t[93] ^ x[6];
  assign t[54] = t[94] ^ x[3];
  assign t[55] = t[95] ^ x[4];
  assign t[56] = t[96] ^ x[5];
  assign t[57] = t[97] ^ x[11];
  assign t[58] = t[98] ^ x[8];
  assign t[59] = t[99] ^ x[9];
  assign t[5] = ~(t[8]);
  assign t[60] = t[100] ^ x[10];
  assign t[61] = t[101] ^ x[16];
  assign t[62] = t[102] ^ x[13];
  assign t[63] = t[103] ^ x[14];
  assign t[64] = t[104] ^ x[15];
  assign t[65] = t[105] ^ x[21];
  assign t[66] = t[106] ^ x[18];
  assign t[67] = t[107] ^ x[19];
  assign t[68] = t[108] ^ x[20];
  assign t[69] = t[109] ^ x[26];
  assign t[6] = ~(t[9]);
  assign t[70] = t[110] ^ x[23];
  assign t[71] = t[111] ^ x[24];
  assign t[72] = t[112] ^ x[25];
  assign t[73] = t[113] ^ x[31];
  assign t[74] = t[114] ^ x[28];
  assign t[75] = t[115] ^ x[29];
  assign t[76] = t[116] ^ x[30];
  assign t[77] = t[117] ^ x[36];
  assign t[78] = t[118] ^ x[33];
  assign t[79] = t[119] ^ x[34];
  assign t[7] = ~(t[10]);
  assign t[80] = t[120] ^ x[35];
  assign t[81] = t[121] ^ x[41];
  assign t[82] = t[122] ^ x[38];
  assign t[83] = t[123] ^ x[39];
  assign t[84] = t[124] ^ x[40];
  assign t[85] = t[125] ^ x[46];
  assign t[86] = t[126] ^ x[43];
  assign t[87] = t[127] ^ x[44];
  assign t[88] = t[128] ^ x[45];
  assign t[89] = t[129] ^ x[51];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[130] ^ x[48];
  assign t[91] = t[131] ^ x[49];
  assign t[92] = t[132] ^ x[50];
  assign t[93] = (x[2]);
  assign t[94] = (x[2]);
  assign t[95] = (x[2]);
  assign t[96] = (x[2]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[7]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind249(x, y);
 input [51:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[7]);
  assign t[101] = (x[12]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[17]);
  assign t[106] = (x[17]);
  assign t[107] = (x[17]);
  assign t[108] = (x[17]);
  assign t[109] = (x[22]);
  assign t[10] = t[15] ^ t[16];
  assign t[110] = (x[22]);
  assign t[111] = (x[22]);
  assign t[112] = (x[22]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[32]);
  assign t[118] = (x[32]);
  assign t[119] = (x[32]);
  assign t[11] = t[24] ^ t[25];
  assign t[120] = (x[32]);
  assign t[121] = (x[37]);
  assign t[122] = (x[37]);
  assign t[123] = (x[37]);
  assign t[124] = (x[37]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[127] = (x[42]);
  assign t[128] = (x[42]);
  assign t[129] = (x[47]);
  assign t[12] = t[17] & t[18];
  assign t[130] = (x[47]);
  assign t[131] = (x[47]);
  assign t[132] = (x[47]);
  assign t[13] = t[26] ^ t[27];
  assign t[14] = t[19] & t[20];
  assign t[15] = t[28] ^ t[29];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[30] ^ t[17]);
  assign t[19] = ~(t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] ^ t[19]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[23]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = t[43] ^ x[6];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[21];
  assign t[37] = t[47] ^ x[26];
  assign t[38] = t[48] ^ x[31];
  assign t[39] = t[49] ^ x[36];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[41];
  assign t[41] = t[51] ^ x[46];
  assign t[42] = t[52] ^ x[51];
  assign t[43] = (~t[53] & t[54] & t[55] & t[56]) | (t[53] & ~t[55] & ~t[56]) | (t[53] & ~t[54] & ~t[56]) | (t[53] & ~t[54] & ~t[55]);
  assign t[44] = (~t[57] & t[58] & t[59] & t[60]) | (t[57] & ~t[59] & ~t[60]) | (t[57] & ~t[58] & ~t[60]) | (t[57] & ~t[58] & ~t[59]);
  assign t[45] = (~t[61] & t[62] & t[63] & t[64]) | (t[61] & ~t[63] & ~t[64]) | (t[61] & ~t[62] & ~t[64]) | (t[61] & ~t[62] & ~t[63]);
  assign t[46] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[47] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[48] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[49] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[51] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[52] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[53] = t[93] ^ x[6];
  assign t[54] = t[94] ^ x[3];
  assign t[55] = t[95] ^ x[4];
  assign t[56] = t[96] ^ x[5];
  assign t[57] = t[97] ^ x[11];
  assign t[58] = t[98] ^ x[8];
  assign t[59] = t[99] ^ x[9];
  assign t[5] = ~(t[8]);
  assign t[60] = t[100] ^ x[10];
  assign t[61] = t[101] ^ x[16];
  assign t[62] = t[102] ^ x[13];
  assign t[63] = t[103] ^ x[14];
  assign t[64] = t[104] ^ x[15];
  assign t[65] = t[105] ^ x[21];
  assign t[66] = t[106] ^ x[18];
  assign t[67] = t[107] ^ x[19];
  assign t[68] = t[108] ^ x[20];
  assign t[69] = t[109] ^ x[26];
  assign t[6] = ~(t[9]);
  assign t[70] = t[110] ^ x[23];
  assign t[71] = t[111] ^ x[24];
  assign t[72] = t[112] ^ x[25];
  assign t[73] = t[113] ^ x[31];
  assign t[74] = t[114] ^ x[28];
  assign t[75] = t[115] ^ x[29];
  assign t[76] = t[116] ^ x[30];
  assign t[77] = t[117] ^ x[36];
  assign t[78] = t[118] ^ x[33];
  assign t[79] = t[119] ^ x[34];
  assign t[7] = ~(t[10]);
  assign t[80] = t[120] ^ x[35];
  assign t[81] = t[121] ^ x[41];
  assign t[82] = t[122] ^ x[38];
  assign t[83] = t[123] ^ x[39];
  assign t[84] = t[124] ^ x[40];
  assign t[85] = t[125] ^ x[46];
  assign t[86] = t[126] ^ x[43];
  assign t[87] = t[127] ^ x[44];
  assign t[88] = t[128] ^ x[45];
  assign t[89] = t[129] ^ x[51];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[130] ^ x[48];
  assign t[91] = t[131] ^ x[49];
  assign t[92] = t[132] ^ x[50];
  assign t[93] = (x[2]);
  assign t[94] = (x[2]);
  assign t[95] = (x[2]);
  assign t[96] = (x[2]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[7]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind250(x, y);
 input [51:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[7]);
  assign t[101] = (x[12]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[17]);
  assign t[106] = (x[17]);
  assign t[107] = (x[17]);
  assign t[108] = (x[17]);
  assign t[109] = (x[22]);
  assign t[10] = t[15] ^ t[16];
  assign t[110] = (x[22]);
  assign t[111] = (x[22]);
  assign t[112] = (x[22]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[32]);
  assign t[118] = (x[32]);
  assign t[119] = (x[32]);
  assign t[11] = t[24] ^ t[25];
  assign t[120] = (x[32]);
  assign t[121] = (x[37]);
  assign t[122] = (x[37]);
  assign t[123] = (x[37]);
  assign t[124] = (x[37]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[127] = (x[42]);
  assign t[128] = (x[42]);
  assign t[129] = (x[47]);
  assign t[12] = t[17] & t[18];
  assign t[130] = (x[47]);
  assign t[131] = (x[47]);
  assign t[132] = (x[47]);
  assign t[13] = t[26] ^ t[27];
  assign t[14] = t[19] & t[20];
  assign t[15] = t[28] ^ t[29];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[30] ^ t[17]);
  assign t[19] = ~(t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] ^ t[19]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[23]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = t[43] ^ x[6];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[21];
  assign t[37] = t[47] ^ x[26];
  assign t[38] = t[48] ^ x[31];
  assign t[39] = t[49] ^ x[36];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[41];
  assign t[41] = t[51] ^ x[46];
  assign t[42] = t[52] ^ x[51];
  assign t[43] = (~t[53] & t[54] & t[55] & t[56]) | (t[53] & ~t[55] & ~t[56]) | (t[53] & ~t[54] & ~t[56]) | (t[53] & ~t[54] & ~t[55]);
  assign t[44] = (~t[57] & t[58] & t[59] & t[60]) | (t[57] & ~t[59] & ~t[60]) | (t[57] & ~t[58] & ~t[60]) | (t[57] & ~t[58] & ~t[59]);
  assign t[45] = (~t[61] & t[62] & t[63] & t[64]) | (t[61] & ~t[63] & ~t[64]) | (t[61] & ~t[62] & ~t[64]) | (t[61] & ~t[62] & ~t[63]);
  assign t[46] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[47] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[48] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[49] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[51] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[52] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[53] = t[93] ^ x[6];
  assign t[54] = t[94] ^ x[3];
  assign t[55] = t[95] ^ x[4];
  assign t[56] = t[96] ^ x[5];
  assign t[57] = t[97] ^ x[11];
  assign t[58] = t[98] ^ x[8];
  assign t[59] = t[99] ^ x[9];
  assign t[5] = ~(t[8]);
  assign t[60] = t[100] ^ x[10];
  assign t[61] = t[101] ^ x[16];
  assign t[62] = t[102] ^ x[13];
  assign t[63] = t[103] ^ x[14];
  assign t[64] = t[104] ^ x[15];
  assign t[65] = t[105] ^ x[21];
  assign t[66] = t[106] ^ x[18];
  assign t[67] = t[107] ^ x[19];
  assign t[68] = t[108] ^ x[20];
  assign t[69] = t[109] ^ x[26];
  assign t[6] = ~(t[9]);
  assign t[70] = t[110] ^ x[23];
  assign t[71] = t[111] ^ x[24];
  assign t[72] = t[112] ^ x[25];
  assign t[73] = t[113] ^ x[31];
  assign t[74] = t[114] ^ x[28];
  assign t[75] = t[115] ^ x[29];
  assign t[76] = t[116] ^ x[30];
  assign t[77] = t[117] ^ x[36];
  assign t[78] = t[118] ^ x[33];
  assign t[79] = t[119] ^ x[34];
  assign t[7] = ~(t[10]);
  assign t[80] = t[120] ^ x[35];
  assign t[81] = t[121] ^ x[41];
  assign t[82] = t[122] ^ x[38];
  assign t[83] = t[123] ^ x[39];
  assign t[84] = t[124] ^ x[40];
  assign t[85] = t[125] ^ x[46];
  assign t[86] = t[126] ^ x[43];
  assign t[87] = t[127] ^ x[44];
  assign t[88] = t[128] ^ x[45];
  assign t[89] = t[129] ^ x[51];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[130] ^ x[48];
  assign t[91] = t[131] ^ x[49];
  assign t[92] = t[132] ^ x[50];
  assign t[93] = (x[2]);
  assign t[94] = (x[2]);
  assign t[95] = (x[2]);
  assign t[96] = (x[2]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[7]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind251(x, y);
 input [51:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[7]);
  assign t[101] = (x[12]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[17]);
  assign t[106] = (x[17]);
  assign t[107] = (x[17]);
  assign t[108] = (x[17]);
  assign t[109] = (x[22]);
  assign t[10] = t[15] ^ t[16];
  assign t[110] = (x[22]);
  assign t[111] = (x[22]);
  assign t[112] = (x[22]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[32]);
  assign t[118] = (x[32]);
  assign t[119] = (x[32]);
  assign t[11] = t[24] ^ t[25];
  assign t[120] = (x[32]);
  assign t[121] = (x[37]);
  assign t[122] = (x[37]);
  assign t[123] = (x[37]);
  assign t[124] = (x[37]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[127] = (x[42]);
  assign t[128] = (x[42]);
  assign t[129] = (x[47]);
  assign t[12] = t[17] & t[18];
  assign t[130] = (x[47]);
  assign t[131] = (x[47]);
  assign t[132] = (x[47]);
  assign t[13] = t[26] ^ t[27];
  assign t[14] = t[19] & t[20];
  assign t[15] = t[28] ^ t[29];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[30] ^ t[17]);
  assign t[19] = ~(t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] ^ t[19]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[23]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = t[43] ^ x[6];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[21];
  assign t[37] = t[47] ^ x[26];
  assign t[38] = t[48] ^ x[31];
  assign t[39] = t[49] ^ x[36];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[41];
  assign t[41] = t[51] ^ x[46];
  assign t[42] = t[52] ^ x[51];
  assign t[43] = (~t[53] & t[54] & t[55] & t[56]) | (t[53] & ~t[55] & ~t[56]) | (t[53] & ~t[54] & ~t[56]) | (t[53] & ~t[54] & ~t[55]);
  assign t[44] = (~t[57] & t[58] & t[59] & t[60]) | (t[57] & ~t[59] & ~t[60]) | (t[57] & ~t[58] & ~t[60]) | (t[57] & ~t[58] & ~t[59]);
  assign t[45] = (~t[61] & t[62] & t[63] & t[64]) | (t[61] & ~t[63] & ~t[64]) | (t[61] & ~t[62] & ~t[64]) | (t[61] & ~t[62] & ~t[63]);
  assign t[46] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[47] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[48] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[49] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[51] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[52] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[53] = t[93] ^ x[6];
  assign t[54] = t[94] ^ x[3];
  assign t[55] = t[95] ^ x[4];
  assign t[56] = t[96] ^ x[5];
  assign t[57] = t[97] ^ x[11];
  assign t[58] = t[98] ^ x[8];
  assign t[59] = t[99] ^ x[9];
  assign t[5] = ~(t[8]);
  assign t[60] = t[100] ^ x[10];
  assign t[61] = t[101] ^ x[16];
  assign t[62] = t[102] ^ x[13];
  assign t[63] = t[103] ^ x[14];
  assign t[64] = t[104] ^ x[15];
  assign t[65] = t[105] ^ x[21];
  assign t[66] = t[106] ^ x[18];
  assign t[67] = t[107] ^ x[19];
  assign t[68] = t[108] ^ x[20];
  assign t[69] = t[109] ^ x[26];
  assign t[6] = ~(t[9]);
  assign t[70] = t[110] ^ x[23];
  assign t[71] = t[111] ^ x[24];
  assign t[72] = t[112] ^ x[25];
  assign t[73] = t[113] ^ x[31];
  assign t[74] = t[114] ^ x[28];
  assign t[75] = t[115] ^ x[29];
  assign t[76] = t[116] ^ x[30];
  assign t[77] = t[117] ^ x[36];
  assign t[78] = t[118] ^ x[33];
  assign t[79] = t[119] ^ x[34];
  assign t[7] = ~(t[10]);
  assign t[80] = t[120] ^ x[35];
  assign t[81] = t[121] ^ x[41];
  assign t[82] = t[122] ^ x[38];
  assign t[83] = t[123] ^ x[39];
  assign t[84] = t[124] ^ x[40];
  assign t[85] = t[125] ^ x[46];
  assign t[86] = t[126] ^ x[43];
  assign t[87] = t[127] ^ x[44];
  assign t[88] = t[128] ^ x[45];
  assign t[89] = t[129] ^ x[51];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[130] ^ x[48];
  assign t[91] = t[131] ^ x[49];
  assign t[92] = t[132] ^ x[50];
  assign t[93] = (x[2]);
  assign t[94] = (x[2]);
  assign t[95] = (x[2]);
  assign t[96] = (x[2]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[7]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind252(x, y);
 input [66:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[34];
  assign t[101] = t[153] ^ x[35];
  assign t[102] = t[154] ^ x[41];
  assign t[103] = t[155] ^ x[38];
  assign t[104] = t[156] ^ x[39];
  assign t[105] = t[157] ^ x[40];
  assign t[106] = t[158] ^ x[46];
  assign t[107] = t[159] ^ x[43];
  assign t[108] = t[160] ^ x[44];
  assign t[109] = t[161] ^ x[45];
  assign t[10] = t[15] ^ t[16];
  assign t[110] = t[162] ^ x[51];
  assign t[111] = t[163] ^ x[48];
  assign t[112] = t[164] ^ x[49];
  assign t[113] = t[165] ^ x[50];
  assign t[114] = t[166] ^ x[56];
  assign t[115] = t[167] ^ x[53];
  assign t[116] = t[168] ^ x[54];
  assign t[117] = t[169] ^ x[55];
  assign t[118] = t[170] ^ x[61];
  assign t[119] = t[171] ^ x[58];
  assign t[11] = t[17] ^ t[18];
  assign t[120] = t[172] ^ x[59];
  assign t[121] = t[173] ^ x[60];
  assign t[122] = t[174] ^ x[66];
  assign t[123] = t[175] ^ x[63];
  assign t[124] = t[176] ^ x[64];
  assign t[125] = t[177] ^ x[65];
  assign t[126] = (x[2]);
  assign t[127] = (x[2]);
  assign t[128] = (x[2]);
  assign t[129] = (x[2]);
  assign t[12] = t[19] & t[20];
  assign t[130] = (x[7]);
  assign t[131] = (x[7]);
  assign t[132] = (x[7]);
  assign t[133] = (x[7]);
  assign t[134] = (x[12]);
  assign t[135] = (x[12]);
  assign t[136] = (x[12]);
  assign t[137] = (x[12]);
  assign t[138] = (x[17]);
  assign t[139] = (x[17]);
  assign t[13] = t[21] ^ t[22];
  assign t[140] = (x[17]);
  assign t[141] = (x[17]);
  assign t[142] = (x[22]);
  assign t[143] = (x[22]);
  assign t[144] = (x[22]);
  assign t[145] = (x[22]);
  assign t[146] = (x[27]);
  assign t[147] = (x[27]);
  assign t[148] = (x[27]);
  assign t[149] = (x[27]);
  assign t[14] = t[23] & t[24];
  assign t[150] = (x[32]);
  assign t[151] = (x[32]);
  assign t[152] = (x[32]);
  assign t[153] = (x[32]);
  assign t[154] = (x[37]);
  assign t[155] = (x[37]);
  assign t[156] = (x[37]);
  assign t[157] = (x[37]);
  assign t[158] = (x[42]);
  assign t[159] = (x[42]);
  assign t[15] = t[25] ^ t[26];
  assign t[160] = (x[42]);
  assign t[161] = (x[42]);
  assign t[162] = (x[47]);
  assign t[163] = (x[47]);
  assign t[164] = (x[47]);
  assign t[165] = (x[47]);
  assign t[166] = (x[52]);
  assign t[167] = (x[52]);
  assign t[168] = (x[52]);
  assign t[169] = (x[52]);
  assign t[16] = t[27] & t[28];
  assign t[170] = (x[57]);
  assign t[171] = (x[57]);
  assign t[172] = (x[57]);
  assign t[173] = (x[57]);
  assign t[174] = (x[62]);
  assign t[175] = (x[62]);
  assign t[176] = (x[62]);
  assign t[177] = (x[62]);
  assign t[17] = t[36] ^ t[37];
  assign t[18] = t[19] & t[29];
  assign t[19] = ~(t[37]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[38] ^ t[19]);
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[23] & t[30];
  assign t[23] = ~(t[40]);
  assign t[24] = ~(t[41] ^ t[23]);
  assign t[25] = t[42] ^ t[43];
  assign t[26] = t[27] & t[31];
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[44] ^ t[27]);
  assign t[29] = t[38] ^ t[32];
  assign t[2] = ~(t[4] ^ t[35]);
  assign t[30] = t[41] ^ t[33];
  assign t[31] = t[44] ^ t[34];
  assign t[32] = t[37] ^ t[45];
  assign t[33] = t[40] ^ t[46];
  assign t[34] = t[43] ^ t[47];
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = t[61] ^ x[6];
  assign t[49] = t[62] ^ x[11];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ x[16];
  assign t[51] = t[64] ^ x[21];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[31];
  assign t[54] = t[67] ^ x[36];
  assign t[55] = t[68] ^ x[41];
  assign t[56] = t[69] ^ x[46];
  assign t[57] = t[70] ^ x[51];
  assign t[58] = t[71] ^ x[56];
  assign t[59] = t[72] ^ x[61];
  assign t[5] = ~(t[8]);
  assign t[60] = t[73] ^ x[66];
  assign t[61] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[62] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[63] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[64] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[65] = (~t[90] & t[91] & t[92] & t[93]) | (t[90] & ~t[92] & ~t[93]) | (t[90] & ~t[91] & ~t[93]) | (t[90] & ~t[91] & ~t[92]);
  assign t[66] = (~t[94] & t[95] & t[96] & t[97]) | (t[94] & ~t[96] & ~t[97]) | (t[94] & ~t[95] & ~t[97]) | (t[94] & ~t[95] & ~t[96]);
  assign t[67] = (~t[98] & t[99] & t[100] & t[101]) | (t[98] & ~t[100] & ~t[101]) | (t[98] & ~t[99] & ~t[101]) | (t[98] & ~t[99] & ~t[100]);
  assign t[68] = (~t[102] & t[103] & t[104] & t[105]) | (t[102] & ~t[104] & ~t[105]) | (t[102] & ~t[103] & ~t[105]) | (t[102] & ~t[103] & ~t[104]);
  assign t[69] = (~t[106] & t[107] & t[108] & t[109]) | (t[106] & ~t[108] & ~t[109]) | (t[106] & ~t[107] & ~t[109]) | (t[106] & ~t[107] & ~t[108]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[110] & t[111] & t[112] & t[113]) | (t[110] & ~t[112] & ~t[113]) | (t[110] & ~t[111] & ~t[113]) | (t[110] & ~t[111] & ~t[112]);
  assign t[71] = (~t[114] & t[115] & t[116] & t[117]) | (t[114] & ~t[116] & ~t[117]) | (t[114] & ~t[115] & ~t[117]) | (t[114] & ~t[115] & ~t[116]);
  assign t[72] = (~t[118] & t[119] & t[120] & t[121]) | (t[118] & ~t[120] & ~t[121]) | (t[118] & ~t[119] & ~t[121]) | (t[118] & ~t[119] & ~t[120]);
  assign t[73] = (~t[122] & t[123] & t[124] & t[125]) | (t[122] & ~t[124] & ~t[125]) | (t[122] & ~t[123] & ~t[125]) | (t[122] & ~t[123] & ~t[124]);
  assign t[74] = t[126] ^ x[6];
  assign t[75] = t[127] ^ x[3];
  assign t[76] = t[128] ^ x[4];
  assign t[77] = t[129] ^ x[5];
  assign t[78] = t[130] ^ x[11];
  assign t[79] = t[131] ^ x[8];
  assign t[7] = ~(t[10]);
  assign t[80] = t[132] ^ x[9];
  assign t[81] = t[133] ^ x[10];
  assign t[82] = t[134] ^ x[16];
  assign t[83] = t[135] ^ x[13];
  assign t[84] = t[136] ^ x[14];
  assign t[85] = t[137] ^ x[15];
  assign t[86] = t[138] ^ x[21];
  assign t[87] = t[139] ^ x[18];
  assign t[88] = t[140] ^ x[19];
  assign t[89] = t[141] ^ x[20];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[142] ^ x[26];
  assign t[91] = t[143] ^ x[23];
  assign t[92] = t[144] ^ x[24];
  assign t[93] = t[145] ^ x[25];
  assign t[94] = t[146] ^ x[31];
  assign t[95] = t[147] ^ x[28];
  assign t[96] = t[148] ^ x[29];
  assign t[97] = t[149] ^ x[30];
  assign t[98] = t[150] ^ x[36];
  assign t[99] = t[151] ^ x[33];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind253(x, y);
 input [66:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[34];
  assign t[101] = t[153] ^ x[35];
  assign t[102] = t[154] ^ x[41];
  assign t[103] = t[155] ^ x[38];
  assign t[104] = t[156] ^ x[39];
  assign t[105] = t[157] ^ x[40];
  assign t[106] = t[158] ^ x[46];
  assign t[107] = t[159] ^ x[43];
  assign t[108] = t[160] ^ x[44];
  assign t[109] = t[161] ^ x[45];
  assign t[10] = t[15] ^ t[16];
  assign t[110] = t[162] ^ x[51];
  assign t[111] = t[163] ^ x[48];
  assign t[112] = t[164] ^ x[49];
  assign t[113] = t[165] ^ x[50];
  assign t[114] = t[166] ^ x[56];
  assign t[115] = t[167] ^ x[53];
  assign t[116] = t[168] ^ x[54];
  assign t[117] = t[169] ^ x[55];
  assign t[118] = t[170] ^ x[61];
  assign t[119] = t[171] ^ x[58];
  assign t[11] = t[17] ^ t[18];
  assign t[120] = t[172] ^ x[59];
  assign t[121] = t[173] ^ x[60];
  assign t[122] = t[174] ^ x[66];
  assign t[123] = t[175] ^ x[63];
  assign t[124] = t[176] ^ x[64];
  assign t[125] = t[177] ^ x[65];
  assign t[126] = (x[2]);
  assign t[127] = (x[2]);
  assign t[128] = (x[2]);
  assign t[129] = (x[2]);
  assign t[12] = t[19] & t[20];
  assign t[130] = (x[7]);
  assign t[131] = (x[7]);
  assign t[132] = (x[7]);
  assign t[133] = (x[7]);
  assign t[134] = (x[12]);
  assign t[135] = (x[12]);
  assign t[136] = (x[12]);
  assign t[137] = (x[12]);
  assign t[138] = (x[17]);
  assign t[139] = (x[17]);
  assign t[13] = t[21] ^ t[22];
  assign t[140] = (x[17]);
  assign t[141] = (x[17]);
  assign t[142] = (x[22]);
  assign t[143] = (x[22]);
  assign t[144] = (x[22]);
  assign t[145] = (x[22]);
  assign t[146] = (x[27]);
  assign t[147] = (x[27]);
  assign t[148] = (x[27]);
  assign t[149] = (x[27]);
  assign t[14] = t[23] & t[24];
  assign t[150] = (x[32]);
  assign t[151] = (x[32]);
  assign t[152] = (x[32]);
  assign t[153] = (x[32]);
  assign t[154] = (x[37]);
  assign t[155] = (x[37]);
  assign t[156] = (x[37]);
  assign t[157] = (x[37]);
  assign t[158] = (x[42]);
  assign t[159] = (x[42]);
  assign t[15] = t[25] ^ t[26];
  assign t[160] = (x[42]);
  assign t[161] = (x[42]);
  assign t[162] = (x[47]);
  assign t[163] = (x[47]);
  assign t[164] = (x[47]);
  assign t[165] = (x[47]);
  assign t[166] = (x[52]);
  assign t[167] = (x[52]);
  assign t[168] = (x[52]);
  assign t[169] = (x[52]);
  assign t[16] = t[27] & t[28];
  assign t[170] = (x[57]);
  assign t[171] = (x[57]);
  assign t[172] = (x[57]);
  assign t[173] = (x[57]);
  assign t[174] = (x[62]);
  assign t[175] = (x[62]);
  assign t[176] = (x[62]);
  assign t[177] = (x[62]);
  assign t[17] = t[36] ^ t[37];
  assign t[18] = t[19] & t[29];
  assign t[19] = ~(t[37]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[38] ^ t[19]);
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[23] & t[30];
  assign t[23] = ~(t[40]);
  assign t[24] = ~(t[41] ^ t[23]);
  assign t[25] = t[42] ^ t[43];
  assign t[26] = t[27] & t[31];
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[44] ^ t[27]);
  assign t[29] = t[38] ^ t[32];
  assign t[2] = ~(t[4] ^ t[35]);
  assign t[30] = t[41] ^ t[33];
  assign t[31] = t[44] ^ t[34];
  assign t[32] = t[37] ^ t[45];
  assign t[33] = t[40] ^ t[46];
  assign t[34] = t[43] ^ t[47];
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = t[61] ^ x[6];
  assign t[49] = t[62] ^ x[11];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ x[16];
  assign t[51] = t[64] ^ x[21];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[31];
  assign t[54] = t[67] ^ x[36];
  assign t[55] = t[68] ^ x[41];
  assign t[56] = t[69] ^ x[46];
  assign t[57] = t[70] ^ x[51];
  assign t[58] = t[71] ^ x[56];
  assign t[59] = t[72] ^ x[61];
  assign t[5] = ~(t[8]);
  assign t[60] = t[73] ^ x[66];
  assign t[61] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[62] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[63] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[64] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[65] = (~t[90] & t[91] & t[92] & t[93]) | (t[90] & ~t[92] & ~t[93]) | (t[90] & ~t[91] & ~t[93]) | (t[90] & ~t[91] & ~t[92]);
  assign t[66] = (~t[94] & t[95] & t[96] & t[97]) | (t[94] & ~t[96] & ~t[97]) | (t[94] & ~t[95] & ~t[97]) | (t[94] & ~t[95] & ~t[96]);
  assign t[67] = (~t[98] & t[99] & t[100] & t[101]) | (t[98] & ~t[100] & ~t[101]) | (t[98] & ~t[99] & ~t[101]) | (t[98] & ~t[99] & ~t[100]);
  assign t[68] = (~t[102] & t[103] & t[104] & t[105]) | (t[102] & ~t[104] & ~t[105]) | (t[102] & ~t[103] & ~t[105]) | (t[102] & ~t[103] & ~t[104]);
  assign t[69] = (~t[106] & t[107] & t[108] & t[109]) | (t[106] & ~t[108] & ~t[109]) | (t[106] & ~t[107] & ~t[109]) | (t[106] & ~t[107] & ~t[108]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[110] & t[111] & t[112] & t[113]) | (t[110] & ~t[112] & ~t[113]) | (t[110] & ~t[111] & ~t[113]) | (t[110] & ~t[111] & ~t[112]);
  assign t[71] = (~t[114] & t[115] & t[116] & t[117]) | (t[114] & ~t[116] & ~t[117]) | (t[114] & ~t[115] & ~t[117]) | (t[114] & ~t[115] & ~t[116]);
  assign t[72] = (~t[118] & t[119] & t[120] & t[121]) | (t[118] & ~t[120] & ~t[121]) | (t[118] & ~t[119] & ~t[121]) | (t[118] & ~t[119] & ~t[120]);
  assign t[73] = (~t[122] & t[123] & t[124] & t[125]) | (t[122] & ~t[124] & ~t[125]) | (t[122] & ~t[123] & ~t[125]) | (t[122] & ~t[123] & ~t[124]);
  assign t[74] = t[126] ^ x[6];
  assign t[75] = t[127] ^ x[3];
  assign t[76] = t[128] ^ x[4];
  assign t[77] = t[129] ^ x[5];
  assign t[78] = t[130] ^ x[11];
  assign t[79] = t[131] ^ x[8];
  assign t[7] = ~(t[10]);
  assign t[80] = t[132] ^ x[9];
  assign t[81] = t[133] ^ x[10];
  assign t[82] = t[134] ^ x[16];
  assign t[83] = t[135] ^ x[13];
  assign t[84] = t[136] ^ x[14];
  assign t[85] = t[137] ^ x[15];
  assign t[86] = t[138] ^ x[21];
  assign t[87] = t[139] ^ x[18];
  assign t[88] = t[140] ^ x[19];
  assign t[89] = t[141] ^ x[20];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[142] ^ x[26];
  assign t[91] = t[143] ^ x[23];
  assign t[92] = t[144] ^ x[24];
  assign t[93] = t[145] ^ x[25];
  assign t[94] = t[146] ^ x[31];
  assign t[95] = t[147] ^ x[28];
  assign t[96] = t[148] ^ x[29];
  assign t[97] = t[149] ^ x[30];
  assign t[98] = t[150] ^ x[36];
  assign t[99] = t[151] ^ x[33];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind254(x, y);
 input [66:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[34];
  assign t[101] = t[153] ^ x[35];
  assign t[102] = t[154] ^ x[41];
  assign t[103] = t[155] ^ x[38];
  assign t[104] = t[156] ^ x[39];
  assign t[105] = t[157] ^ x[40];
  assign t[106] = t[158] ^ x[46];
  assign t[107] = t[159] ^ x[43];
  assign t[108] = t[160] ^ x[44];
  assign t[109] = t[161] ^ x[45];
  assign t[10] = t[15] ^ t[16];
  assign t[110] = t[162] ^ x[51];
  assign t[111] = t[163] ^ x[48];
  assign t[112] = t[164] ^ x[49];
  assign t[113] = t[165] ^ x[50];
  assign t[114] = t[166] ^ x[56];
  assign t[115] = t[167] ^ x[53];
  assign t[116] = t[168] ^ x[54];
  assign t[117] = t[169] ^ x[55];
  assign t[118] = t[170] ^ x[61];
  assign t[119] = t[171] ^ x[58];
  assign t[11] = t[17] ^ t[18];
  assign t[120] = t[172] ^ x[59];
  assign t[121] = t[173] ^ x[60];
  assign t[122] = t[174] ^ x[66];
  assign t[123] = t[175] ^ x[63];
  assign t[124] = t[176] ^ x[64];
  assign t[125] = t[177] ^ x[65];
  assign t[126] = (x[2]);
  assign t[127] = (x[2]);
  assign t[128] = (x[2]);
  assign t[129] = (x[2]);
  assign t[12] = t[19] & t[20];
  assign t[130] = (x[7]);
  assign t[131] = (x[7]);
  assign t[132] = (x[7]);
  assign t[133] = (x[7]);
  assign t[134] = (x[12]);
  assign t[135] = (x[12]);
  assign t[136] = (x[12]);
  assign t[137] = (x[12]);
  assign t[138] = (x[17]);
  assign t[139] = (x[17]);
  assign t[13] = t[21] ^ t[22];
  assign t[140] = (x[17]);
  assign t[141] = (x[17]);
  assign t[142] = (x[22]);
  assign t[143] = (x[22]);
  assign t[144] = (x[22]);
  assign t[145] = (x[22]);
  assign t[146] = (x[27]);
  assign t[147] = (x[27]);
  assign t[148] = (x[27]);
  assign t[149] = (x[27]);
  assign t[14] = t[23] & t[24];
  assign t[150] = (x[32]);
  assign t[151] = (x[32]);
  assign t[152] = (x[32]);
  assign t[153] = (x[32]);
  assign t[154] = (x[37]);
  assign t[155] = (x[37]);
  assign t[156] = (x[37]);
  assign t[157] = (x[37]);
  assign t[158] = (x[42]);
  assign t[159] = (x[42]);
  assign t[15] = t[25] ^ t[26];
  assign t[160] = (x[42]);
  assign t[161] = (x[42]);
  assign t[162] = (x[47]);
  assign t[163] = (x[47]);
  assign t[164] = (x[47]);
  assign t[165] = (x[47]);
  assign t[166] = (x[52]);
  assign t[167] = (x[52]);
  assign t[168] = (x[52]);
  assign t[169] = (x[52]);
  assign t[16] = t[27] & t[28];
  assign t[170] = (x[57]);
  assign t[171] = (x[57]);
  assign t[172] = (x[57]);
  assign t[173] = (x[57]);
  assign t[174] = (x[62]);
  assign t[175] = (x[62]);
  assign t[176] = (x[62]);
  assign t[177] = (x[62]);
  assign t[17] = t[36] ^ t[37];
  assign t[18] = t[19] & t[29];
  assign t[19] = ~(t[37]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[38] ^ t[19]);
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[23] & t[30];
  assign t[23] = ~(t[40]);
  assign t[24] = ~(t[41] ^ t[23]);
  assign t[25] = t[42] ^ t[43];
  assign t[26] = t[27] & t[31];
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[44] ^ t[27]);
  assign t[29] = t[38] ^ t[32];
  assign t[2] = ~(t[4] ^ t[35]);
  assign t[30] = t[41] ^ t[33];
  assign t[31] = t[44] ^ t[34];
  assign t[32] = t[37] ^ t[45];
  assign t[33] = t[40] ^ t[46];
  assign t[34] = t[43] ^ t[47];
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = t[61] ^ x[6];
  assign t[49] = t[62] ^ x[11];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ x[16];
  assign t[51] = t[64] ^ x[21];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[31];
  assign t[54] = t[67] ^ x[36];
  assign t[55] = t[68] ^ x[41];
  assign t[56] = t[69] ^ x[46];
  assign t[57] = t[70] ^ x[51];
  assign t[58] = t[71] ^ x[56];
  assign t[59] = t[72] ^ x[61];
  assign t[5] = ~(t[8]);
  assign t[60] = t[73] ^ x[66];
  assign t[61] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[62] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[63] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[64] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[65] = (~t[90] & t[91] & t[92] & t[93]) | (t[90] & ~t[92] & ~t[93]) | (t[90] & ~t[91] & ~t[93]) | (t[90] & ~t[91] & ~t[92]);
  assign t[66] = (~t[94] & t[95] & t[96] & t[97]) | (t[94] & ~t[96] & ~t[97]) | (t[94] & ~t[95] & ~t[97]) | (t[94] & ~t[95] & ~t[96]);
  assign t[67] = (~t[98] & t[99] & t[100] & t[101]) | (t[98] & ~t[100] & ~t[101]) | (t[98] & ~t[99] & ~t[101]) | (t[98] & ~t[99] & ~t[100]);
  assign t[68] = (~t[102] & t[103] & t[104] & t[105]) | (t[102] & ~t[104] & ~t[105]) | (t[102] & ~t[103] & ~t[105]) | (t[102] & ~t[103] & ~t[104]);
  assign t[69] = (~t[106] & t[107] & t[108] & t[109]) | (t[106] & ~t[108] & ~t[109]) | (t[106] & ~t[107] & ~t[109]) | (t[106] & ~t[107] & ~t[108]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[110] & t[111] & t[112] & t[113]) | (t[110] & ~t[112] & ~t[113]) | (t[110] & ~t[111] & ~t[113]) | (t[110] & ~t[111] & ~t[112]);
  assign t[71] = (~t[114] & t[115] & t[116] & t[117]) | (t[114] & ~t[116] & ~t[117]) | (t[114] & ~t[115] & ~t[117]) | (t[114] & ~t[115] & ~t[116]);
  assign t[72] = (~t[118] & t[119] & t[120] & t[121]) | (t[118] & ~t[120] & ~t[121]) | (t[118] & ~t[119] & ~t[121]) | (t[118] & ~t[119] & ~t[120]);
  assign t[73] = (~t[122] & t[123] & t[124] & t[125]) | (t[122] & ~t[124] & ~t[125]) | (t[122] & ~t[123] & ~t[125]) | (t[122] & ~t[123] & ~t[124]);
  assign t[74] = t[126] ^ x[6];
  assign t[75] = t[127] ^ x[3];
  assign t[76] = t[128] ^ x[4];
  assign t[77] = t[129] ^ x[5];
  assign t[78] = t[130] ^ x[11];
  assign t[79] = t[131] ^ x[8];
  assign t[7] = ~(t[10]);
  assign t[80] = t[132] ^ x[9];
  assign t[81] = t[133] ^ x[10];
  assign t[82] = t[134] ^ x[16];
  assign t[83] = t[135] ^ x[13];
  assign t[84] = t[136] ^ x[14];
  assign t[85] = t[137] ^ x[15];
  assign t[86] = t[138] ^ x[21];
  assign t[87] = t[139] ^ x[18];
  assign t[88] = t[140] ^ x[19];
  assign t[89] = t[141] ^ x[20];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[142] ^ x[26];
  assign t[91] = t[143] ^ x[23];
  assign t[92] = t[144] ^ x[24];
  assign t[93] = t[145] ^ x[25];
  assign t[94] = t[146] ^ x[31];
  assign t[95] = t[147] ^ x[28];
  assign t[96] = t[148] ^ x[29];
  assign t[97] = t[149] ^ x[30];
  assign t[98] = t[150] ^ x[36];
  assign t[99] = t[151] ^ x[33];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind255(x, y);
 input [66:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[34];
  assign t[101] = t[153] ^ x[35];
  assign t[102] = t[154] ^ x[41];
  assign t[103] = t[155] ^ x[38];
  assign t[104] = t[156] ^ x[39];
  assign t[105] = t[157] ^ x[40];
  assign t[106] = t[158] ^ x[46];
  assign t[107] = t[159] ^ x[43];
  assign t[108] = t[160] ^ x[44];
  assign t[109] = t[161] ^ x[45];
  assign t[10] = t[15] ^ t[16];
  assign t[110] = t[162] ^ x[51];
  assign t[111] = t[163] ^ x[48];
  assign t[112] = t[164] ^ x[49];
  assign t[113] = t[165] ^ x[50];
  assign t[114] = t[166] ^ x[56];
  assign t[115] = t[167] ^ x[53];
  assign t[116] = t[168] ^ x[54];
  assign t[117] = t[169] ^ x[55];
  assign t[118] = t[170] ^ x[61];
  assign t[119] = t[171] ^ x[58];
  assign t[11] = t[17] ^ t[18];
  assign t[120] = t[172] ^ x[59];
  assign t[121] = t[173] ^ x[60];
  assign t[122] = t[174] ^ x[66];
  assign t[123] = t[175] ^ x[63];
  assign t[124] = t[176] ^ x[64];
  assign t[125] = t[177] ^ x[65];
  assign t[126] = (x[2]);
  assign t[127] = (x[2]);
  assign t[128] = (x[2]);
  assign t[129] = (x[2]);
  assign t[12] = t[19] & t[20];
  assign t[130] = (x[7]);
  assign t[131] = (x[7]);
  assign t[132] = (x[7]);
  assign t[133] = (x[7]);
  assign t[134] = (x[12]);
  assign t[135] = (x[12]);
  assign t[136] = (x[12]);
  assign t[137] = (x[12]);
  assign t[138] = (x[17]);
  assign t[139] = (x[17]);
  assign t[13] = t[21] ^ t[22];
  assign t[140] = (x[17]);
  assign t[141] = (x[17]);
  assign t[142] = (x[22]);
  assign t[143] = (x[22]);
  assign t[144] = (x[22]);
  assign t[145] = (x[22]);
  assign t[146] = (x[27]);
  assign t[147] = (x[27]);
  assign t[148] = (x[27]);
  assign t[149] = (x[27]);
  assign t[14] = t[23] & t[24];
  assign t[150] = (x[32]);
  assign t[151] = (x[32]);
  assign t[152] = (x[32]);
  assign t[153] = (x[32]);
  assign t[154] = (x[37]);
  assign t[155] = (x[37]);
  assign t[156] = (x[37]);
  assign t[157] = (x[37]);
  assign t[158] = (x[42]);
  assign t[159] = (x[42]);
  assign t[15] = t[25] ^ t[26];
  assign t[160] = (x[42]);
  assign t[161] = (x[42]);
  assign t[162] = (x[47]);
  assign t[163] = (x[47]);
  assign t[164] = (x[47]);
  assign t[165] = (x[47]);
  assign t[166] = (x[52]);
  assign t[167] = (x[52]);
  assign t[168] = (x[52]);
  assign t[169] = (x[52]);
  assign t[16] = t[27] & t[28];
  assign t[170] = (x[57]);
  assign t[171] = (x[57]);
  assign t[172] = (x[57]);
  assign t[173] = (x[57]);
  assign t[174] = (x[62]);
  assign t[175] = (x[62]);
  assign t[176] = (x[62]);
  assign t[177] = (x[62]);
  assign t[17] = t[36] ^ t[37];
  assign t[18] = t[19] & t[29];
  assign t[19] = ~(t[37]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[38] ^ t[19]);
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[23] & t[30];
  assign t[23] = ~(t[40]);
  assign t[24] = ~(t[41] ^ t[23]);
  assign t[25] = t[42] ^ t[43];
  assign t[26] = t[27] & t[31];
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[44] ^ t[27]);
  assign t[29] = t[38] ^ t[32];
  assign t[2] = ~(t[4] ^ t[35]);
  assign t[30] = t[41] ^ t[33];
  assign t[31] = t[44] ^ t[34];
  assign t[32] = t[37] ^ t[45];
  assign t[33] = t[40] ^ t[46];
  assign t[34] = t[43] ^ t[47];
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = t[61] ^ x[6];
  assign t[49] = t[62] ^ x[11];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ x[16];
  assign t[51] = t[64] ^ x[21];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[31];
  assign t[54] = t[67] ^ x[36];
  assign t[55] = t[68] ^ x[41];
  assign t[56] = t[69] ^ x[46];
  assign t[57] = t[70] ^ x[51];
  assign t[58] = t[71] ^ x[56];
  assign t[59] = t[72] ^ x[61];
  assign t[5] = ~(t[8]);
  assign t[60] = t[73] ^ x[66];
  assign t[61] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[62] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[63] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[64] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[65] = (~t[90] & t[91] & t[92] & t[93]) | (t[90] & ~t[92] & ~t[93]) | (t[90] & ~t[91] & ~t[93]) | (t[90] & ~t[91] & ~t[92]);
  assign t[66] = (~t[94] & t[95] & t[96] & t[97]) | (t[94] & ~t[96] & ~t[97]) | (t[94] & ~t[95] & ~t[97]) | (t[94] & ~t[95] & ~t[96]);
  assign t[67] = (~t[98] & t[99] & t[100] & t[101]) | (t[98] & ~t[100] & ~t[101]) | (t[98] & ~t[99] & ~t[101]) | (t[98] & ~t[99] & ~t[100]);
  assign t[68] = (~t[102] & t[103] & t[104] & t[105]) | (t[102] & ~t[104] & ~t[105]) | (t[102] & ~t[103] & ~t[105]) | (t[102] & ~t[103] & ~t[104]);
  assign t[69] = (~t[106] & t[107] & t[108] & t[109]) | (t[106] & ~t[108] & ~t[109]) | (t[106] & ~t[107] & ~t[109]) | (t[106] & ~t[107] & ~t[108]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[110] & t[111] & t[112] & t[113]) | (t[110] & ~t[112] & ~t[113]) | (t[110] & ~t[111] & ~t[113]) | (t[110] & ~t[111] & ~t[112]);
  assign t[71] = (~t[114] & t[115] & t[116] & t[117]) | (t[114] & ~t[116] & ~t[117]) | (t[114] & ~t[115] & ~t[117]) | (t[114] & ~t[115] & ~t[116]);
  assign t[72] = (~t[118] & t[119] & t[120] & t[121]) | (t[118] & ~t[120] & ~t[121]) | (t[118] & ~t[119] & ~t[121]) | (t[118] & ~t[119] & ~t[120]);
  assign t[73] = (~t[122] & t[123] & t[124] & t[125]) | (t[122] & ~t[124] & ~t[125]) | (t[122] & ~t[123] & ~t[125]) | (t[122] & ~t[123] & ~t[124]);
  assign t[74] = t[126] ^ x[6];
  assign t[75] = t[127] ^ x[3];
  assign t[76] = t[128] ^ x[4];
  assign t[77] = t[129] ^ x[5];
  assign t[78] = t[130] ^ x[11];
  assign t[79] = t[131] ^ x[8];
  assign t[7] = ~(t[10]);
  assign t[80] = t[132] ^ x[9];
  assign t[81] = t[133] ^ x[10];
  assign t[82] = t[134] ^ x[16];
  assign t[83] = t[135] ^ x[13];
  assign t[84] = t[136] ^ x[14];
  assign t[85] = t[137] ^ x[15];
  assign t[86] = t[138] ^ x[21];
  assign t[87] = t[139] ^ x[18];
  assign t[88] = t[140] ^ x[19];
  assign t[89] = t[141] ^ x[20];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[142] ^ x[26];
  assign t[91] = t[143] ^ x[23];
  assign t[92] = t[144] ^ x[24];
  assign t[93] = t[145] ^ x[25];
  assign t[94] = t[146] ^ x[31];
  assign t[95] = t[147] ^ x[28];
  assign t[96] = t[148] ^ x[29];
  assign t[97] = t[149] ^ x[30];
  assign t[98] = t[150] ^ x[36];
  assign t[99] = t[151] ^ x[33];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind256(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[54] & t[26];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[55] & t[31];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[56] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[54] ^ t[27]);
  assign t[29] = t[58] ^ t[57];
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[55] ^ t[32]);
  assign t[34] = t[60] ^ t[59];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[56] ^ t[37]);
  assign t[39] = t[62] ^ t[61];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[54] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[54] ^ t[50];
  assign t[44] = t[55] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[55] ^ t[51];
  assign t[47] = t[56] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[56] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[57] ^ t[63];
  assign t[51] = t[59] ^ t[64];
  assign t[52] = t[61] ^ t[65];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] & t[17];
  assign y = (t[0]);
endmodule

module R2ind257(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[54] & t[26];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[55] & t[31];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[56] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[54] ^ t[27]);
  assign t[29] = t[58] ^ t[57];
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[55] ^ t[32]);
  assign t[34] = t[60] ^ t[59];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[56] ^ t[37]);
  assign t[39] = t[62] ^ t[61];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[54] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[54] ^ t[50];
  assign t[44] = t[55] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[55] ^ t[51];
  assign t[47] = t[56] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[56] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[57] ^ t[63];
  assign t[51] = t[59] ^ t[64];
  assign t[52] = t[61] ^ t[65];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] & t[17];
  assign y = (t[0]);
endmodule

module R2ind258(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[54] & t[26];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[55] & t[31];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[56] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[54] ^ t[27]);
  assign t[29] = t[58] ^ t[57];
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[55] ^ t[32]);
  assign t[34] = t[60] ^ t[59];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[56] ^ t[37]);
  assign t[39] = t[62] ^ t[61];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[54] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[54] ^ t[50];
  assign t[44] = t[55] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[55] ^ t[51];
  assign t[47] = t[56] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[56] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[57] ^ t[63];
  assign t[51] = t[59] ^ t[64];
  assign t[52] = t[61] ^ t[65];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] & t[17];
  assign y = (t[0]);
endmodule

module R2ind259(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[54] & t[26];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[55] & t[31];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[56] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[54] ^ t[27]);
  assign t[29] = t[58] ^ t[57];
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[55] ^ t[32]);
  assign t[34] = t[60] ^ t[59];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[56] ^ t[37]);
  assign t[39] = t[62] ^ t[61];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[54] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[54] ^ t[50];
  assign t[44] = t[55] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[55] ^ t[51];
  assign t[47] = t[56] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[56] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[57] ^ t[63];
  assign t[51] = t[59] ^ t[64];
  assign t[52] = t[61] ^ t[65];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] & t[17];
  assign y = (t[0]);
endmodule

module R2ind260(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[26] ^ t[27];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[28] & t[29];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[30] ^ t[15];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[54] ^ t[28];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[31] ^ t[32];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[55] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[56] ^ t[38];
  assign t[26] = t[57] ^ t[58];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[58]);
  assign t[29] = ~(t[54] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = t[54] & t[42];
  assign t[31] = t[59] ^ t[60];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[60]);
  assign t[34] = ~(t[55] ^ t[33]);
  assign t[35] = t[55] & t[44];
  assign t[36] = t[61] ^ t[62];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[62]);
  assign t[39] = ~(t[56] ^ t[38]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[56] & t[46];
  assign t[41] = t[54] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[55] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[56] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[58] ^ t[63];
  assign t[48] = t[54] ^ t[26];
  assign t[49] = t[60] ^ t[64];
  assign t[4] = ~t[7];
  assign t[50] = t[55] ^ t[31];
  assign t[51] = t[62] ^ t[65];
  assign t[52] = t[56] ^ t[36];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind261(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[26] ^ t[27];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[28] & t[29];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[30] ^ t[15];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[54] ^ t[28];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[31] ^ t[32];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[55] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[56] ^ t[38];
  assign t[26] = t[57] ^ t[58];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[58]);
  assign t[29] = ~(t[54] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = t[54] & t[42];
  assign t[31] = t[59] ^ t[60];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[60]);
  assign t[34] = ~(t[55] ^ t[33]);
  assign t[35] = t[55] & t[44];
  assign t[36] = t[61] ^ t[62];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[62]);
  assign t[39] = ~(t[56] ^ t[38]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[56] & t[46];
  assign t[41] = t[54] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[55] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[56] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[58] ^ t[63];
  assign t[48] = t[54] ^ t[26];
  assign t[49] = t[60] ^ t[64];
  assign t[4] = ~t[7];
  assign t[50] = t[55] ^ t[31];
  assign t[51] = t[62] ^ t[65];
  assign t[52] = t[56] ^ t[36];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind262(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[26] ^ t[27];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[28] & t[29];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[30] ^ t[15];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[54] ^ t[28];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[31] ^ t[32];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[55] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[56] ^ t[38];
  assign t[26] = t[57] ^ t[58];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[58]);
  assign t[29] = ~(t[54] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = t[54] & t[42];
  assign t[31] = t[59] ^ t[60];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[60]);
  assign t[34] = ~(t[55] ^ t[33]);
  assign t[35] = t[55] & t[44];
  assign t[36] = t[61] ^ t[62];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[62]);
  assign t[39] = ~(t[56] ^ t[38]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[56] & t[46];
  assign t[41] = t[54] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[55] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[56] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[58] ^ t[63];
  assign t[48] = t[54] ^ t[26];
  assign t[49] = t[60] ^ t[64];
  assign t[4] = ~t[7];
  assign t[50] = t[55] ^ t[31];
  assign t[51] = t[62] ^ t[65];
  assign t[52] = t[56] ^ t[36];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind263(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[16];
  assign t[101] = t[153] ^ x[13];
  assign t[102] = t[154] ^ x[14];
  assign t[103] = t[155] ^ x[15];
  assign t[104] = t[156] ^ x[21];
  assign t[105] = t[157] ^ x[18];
  assign t[106] = t[158] ^ x[19];
  assign t[107] = t[159] ^ x[20];
  assign t[108] = t[160] ^ x[26];
  assign t[109] = t[161] ^ x[23];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[162] ^ x[24];
  assign t[111] = t[163] ^ x[25];
  assign t[112] = t[164] ^ x[31];
  assign t[113] = t[165] ^ x[28];
  assign t[114] = t[166] ^ x[29];
  assign t[115] = t[167] ^ x[30];
  assign t[116] = t[168] ^ x[36];
  assign t[117] = t[169] ^ x[33];
  assign t[118] = t[170] ^ x[34];
  assign t[119] = t[171] ^ x[35];
  assign t[11] = t[20] ^ t[21];
  assign t[120] = t[172] ^ x[41];
  assign t[121] = t[173] ^ x[38];
  assign t[122] = t[174] ^ x[39];
  assign t[123] = t[175] ^ x[40];
  assign t[124] = t[176] ^ x[46];
  assign t[125] = t[177] ^ x[43];
  assign t[126] = t[178] ^ x[44];
  assign t[127] = t[179] ^ x[45];
  assign t[128] = t[180] ^ x[51];
  assign t[129] = t[181] ^ x[48];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[182] ^ x[49];
  assign t[131] = t[183] ^ x[50];
  assign t[132] = t[184] ^ x[56];
  assign t[133] = t[185] ^ x[53];
  assign t[134] = t[186] ^ x[54];
  assign t[135] = t[187] ^ x[55];
  assign t[136] = t[188] ^ x[61];
  assign t[137] = t[189] ^ x[58];
  assign t[138] = t[190] ^ x[59];
  assign t[139] = t[191] ^ x[60];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[192] ^ x[66];
  assign t[141] = t[193] ^ x[63];
  assign t[142] = t[194] ^ x[64];
  assign t[143] = t[195] ^ x[65];
  assign t[144] = (x[2]);
  assign t[145] = (x[2]);
  assign t[146] = (x[2]);
  assign t[147] = (x[2]);
  assign t[148] = (x[7]);
  assign t[149] = (x[7]);
  assign t[14] = t[26] ^ t[27];
  assign t[150] = (x[7]);
  assign t[151] = (x[7]);
  assign t[152] = (x[12]);
  assign t[153] = (x[12]);
  assign t[154] = (x[12]);
  assign t[155] = (x[12]);
  assign t[156] = (x[17]);
  assign t[157] = (x[17]);
  assign t[158] = (x[17]);
  assign t[159] = (x[17]);
  assign t[15] = t[28] & t[29];
  assign t[160] = (x[22]);
  assign t[161] = (x[22]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[27]);
  assign t[165] = (x[27]);
  assign t[166] = (x[27]);
  assign t[167] = (x[27]);
  assign t[168] = (x[32]);
  assign t[169] = (x[32]);
  assign t[16] = t[30] ^ t[15];
  assign t[170] = (x[32]);
  assign t[171] = (x[32]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[42]);
  assign t[177] = (x[42]);
  assign t[178] = (x[42]);
  assign t[179] = (x[42]);
  assign t[17] = t[54] ^ t[28];
  assign t[180] = (x[47]);
  assign t[181] = (x[47]);
  assign t[182] = (x[47]);
  assign t[183] = (x[47]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[52]);
  assign t[187] = (x[52]);
  assign t[188] = (x[57]);
  assign t[189] = (x[57]);
  assign t[18] = t[31] ^ t[32];
  assign t[190] = (x[57]);
  assign t[191] = (x[57]);
  assign t[192] = (x[62]);
  assign t[193] = (x[62]);
  assign t[194] = (x[62]);
  assign t[195] = (x[62]);
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[55] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[56] ^ t[38];
  assign t[26] = t[57] ^ t[58];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[58]);
  assign t[29] = ~(t[54] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[53]);
  assign t[30] = t[54] & t[42];
  assign t[31] = t[59] ^ t[60];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[60]);
  assign t[34] = ~(t[55] ^ t[33]);
  assign t[35] = t[55] & t[44];
  assign t[36] = t[61] ^ t[62];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[62]);
  assign t[39] = ~(t[56] ^ t[38]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[56] & t[46];
  assign t[41] = t[54] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[55] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[56] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[58] ^ t[63];
  assign t[48] = t[54] ^ t[26];
  assign t[49] = t[60] ^ t[64];
  assign t[4] = ~t[7];
  assign t[50] = t[55] ^ t[31];
  assign t[51] = t[62] ^ t[65];
  assign t[52] = t[56] ^ t[36];
  assign t[53] = (t[66]);
  assign t[54] = (t[67]);
  assign t[55] = (t[68]);
  assign t[56] = (t[69]);
  assign t[57] = (t[70]);
  assign t[58] = (t[71]);
  assign t[59] = (t[72]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (t[73]);
  assign t[61] = (t[74]);
  assign t[62] = (t[75]);
  assign t[63] = (t[76]);
  assign t[64] = (t[77]);
  assign t[65] = (t[78]);
  assign t[66] = t[79] ^ x[6];
  assign t[67] = t[80] ^ x[11];
  assign t[68] = t[81] ^ x[16];
  assign t[69] = t[82] ^ x[21];
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = t[83] ^ x[26];
  assign t[71] = t[84] ^ x[31];
  assign t[72] = t[85] ^ x[36];
  assign t[73] = t[86] ^ x[41];
  assign t[74] = t[87] ^ x[46];
  assign t[75] = t[88] ^ x[51];
  assign t[76] = t[89] ^ x[56];
  assign t[77] = t[90] ^ x[61];
  assign t[78] = t[91] ^ x[66];
  assign t[79] = (~t[92] & t[93] & t[94] & t[95]) | (t[92] & ~t[94] & ~t[95]) | (t[92] & ~t[93] & ~t[95]) | (t[92] & ~t[93] & ~t[94]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[96] & t[97] & t[98] & t[99]) | (t[96] & ~t[98] & ~t[99]) | (t[96] & ~t[97] & ~t[99]) | (t[96] & ~t[97] & ~t[98]);
  assign t[81] = (~t[100] & t[101] & t[102] & t[103]) | (t[100] & ~t[102] & ~t[103]) | (t[100] & ~t[101] & ~t[103]) | (t[100] & ~t[101] & ~t[102]);
  assign t[82] = (~t[104] & t[105] & t[106] & t[107]) | (t[104] & ~t[106] & ~t[107]) | (t[104] & ~t[105] & ~t[107]) | (t[104] & ~t[105] & ~t[106]);
  assign t[83] = (~t[108] & t[109] & t[110] & t[111]) | (t[108] & ~t[110] & ~t[111]) | (t[108] & ~t[109] & ~t[111]) | (t[108] & ~t[109] & ~t[110]);
  assign t[84] = (~t[112] & t[113] & t[114] & t[115]) | (t[112] & ~t[114] & ~t[115]) | (t[112] & ~t[113] & ~t[115]) | (t[112] & ~t[113] & ~t[114]);
  assign t[85] = (~t[116] & t[117] & t[118] & t[119]) | (t[116] & ~t[118] & ~t[119]) | (t[116] & ~t[117] & ~t[119]) | (t[116] & ~t[117] & ~t[118]);
  assign t[86] = (~t[120] & t[121] & t[122] & t[123]) | (t[120] & ~t[122] & ~t[123]) | (t[120] & ~t[121] & ~t[123]) | (t[120] & ~t[121] & ~t[122]);
  assign t[87] = (~t[124] & t[125] & t[126] & t[127]) | (t[124] & ~t[126] & ~t[127]) | (t[124] & ~t[125] & ~t[127]) | (t[124] & ~t[125] & ~t[126]);
  assign t[88] = (~t[128] & t[129] & t[130] & t[131]) | (t[128] & ~t[130] & ~t[131]) | (t[128] & ~t[129] & ~t[131]) | (t[128] & ~t[129] & ~t[130]);
  assign t[89] = (~t[132] & t[133] & t[134] & t[135]) | (t[132] & ~t[134] & ~t[135]) | (t[132] & ~t[133] & ~t[135]) | (t[132] & ~t[133] & ~t[134]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (~t[136] & t[137] & t[138] & t[139]) | (t[136] & ~t[138] & ~t[139]) | (t[136] & ~t[137] & ~t[139]) | (t[136] & ~t[137] & ~t[138]);
  assign t[91] = (~t[140] & t[141] & t[142] & t[143]) | (t[140] & ~t[142] & ~t[143]) | (t[140] & ~t[141] & ~t[143]) | (t[140] & ~t[141] & ~t[142]);
  assign t[92] = t[144] ^ x[6];
  assign t[93] = t[145] ^ x[3];
  assign t[94] = t[146] ^ x[4];
  assign t[95] = t[147] ^ x[5];
  assign t[96] = t[148] ^ x[11];
  assign t[97] = t[149] ^ x[8];
  assign t[98] = t[150] ^ x[9];
  assign t[99] = t[151] ^ x[10];
  assign t[9] = t[16] ^ t[17];
  assign y = (t[0]);
endmodule

module R2ind264(x, y);
 input [51:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[7]);
  assign t[101] = (x[12]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[17]);
  assign t[106] = (x[17]);
  assign t[107] = (x[17]);
  assign t[108] = (x[17]);
  assign t[109] = (x[22]);
  assign t[10] = t[15] ^ t[16];
  assign t[110] = (x[22]);
  assign t[111] = (x[22]);
  assign t[112] = (x[22]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[32]);
  assign t[118] = (x[32]);
  assign t[119] = (x[32]);
  assign t[11] = t[24] ^ t[25];
  assign t[120] = (x[32]);
  assign t[121] = (x[37]);
  assign t[122] = (x[37]);
  assign t[123] = (x[37]);
  assign t[124] = (x[37]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[127] = (x[42]);
  assign t[128] = (x[42]);
  assign t[129] = (x[47]);
  assign t[12] = t[17] & t[18];
  assign t[130] = (x[47]);
  assign t[131] = (x[47]);
  assign t[132] = (x[47]);
  assign t[13] = t[26] ^ t[27];
  assign t[14] = t[19] & t[20];
  assign t[15] = t[28] ^ t[29];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[30] ^ t[17]);
  assign t[19] = ~(t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] ^ t[19]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[23]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = t[43] ^ x[6];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[21];
  assign t[37] = t[47] ^ x[26];
  assign t[38] = t[48] ^ x[31];
  assign t[39] = t[49] ^ x[36];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[41];
  assign t[41] = t[51] ^ x[46];
  assign t[42] = t[52] ^ x[51];
  assign t[43] = (~t[53] & t[54] & t[55] & t[56]) | (t[53] & ~t[55] & ~t[56]) | (t[53] & ~t[54] & ~t[56]) | (t[53] & ~t[54] & ~t[55]);
  assign t[44] = (~t[57] & t[58] & t[59] & t[60]) | (t[57] & ~t[59] & ~t[60]) | (t[57] & ~t[58] & ~t[60]) | (t[57] & ~t[58] & ~t[59]);
  assign t[45] = (~t[61] & t[62] & t[63] & t[64]) | (t[61] & ~t[63] & ~t[64]) | (t[61] & ~t[62] & ~t[64]) | (t[61] & ~t[62] & ~t[63]);
  assign t[46] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[47] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[48] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[49] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[51] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[52] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[53] = t[93] ^ x[6];
  assign t[54] = t[94] ^ x[3];
  assign t[55] = t[95] ^ x[4];
  assign t[56] = t[96] ^ x[5];
  assign t[57] = t[97] ^ x[11];
  assign t[58] = t[98] ^ x[8];
  assign t[59] = t[99] ^ x[9];
  assign t[5] = ~(t[8]);
  assign t[60] = t[100] ^ x[10];
  assign t[61] = t[101] ^ x[16];
  assign t[62] = t[102] ^ x[13];
  assign t[63] = t[103] ^ x[14];
  assign t[64] = t[104] ^ x[15];
  assign t[65] = t[105] ^ x[21];
  assign t[66] = t[106] ^ x[18];
  assign t[67] = t[107] ^ x[19];
  assign t[68] = t[108] ^ x[20];
  assign t[69] = t[109] ^ x[26];
  assign t[6] = ~(t[9]);
  assign t[70] = t[110] ^ x[23];
  assign t[71] = t[111] ^ x[24];
  assign t[72] = t[112] ^ x[25];
  assign t[73] = t[113] ^ x[31];
  assign t[74] = t[114] ^ x[28];
  assign t[75] = t[115] ^ x[29];
  assign t[76] = t[116] ^ x[30];
  assign t[77] = t[117] ^ x[36];
  assign t[78] = t[118] ^ x[33];
  assign t[79] = t[119] ^ x[34];
  assign t[7] = ~(t[10]);
  assign t[80] = t[120] ^ x[35];
  assign t[81] = t[121] ^ x[41];
  assign t[82] = t[122] ^ x[38];
  assign t[83] = t[123] ^ x[39];
  assign t[84] = t[124] ^ x[40];
  assign t[85] = t[125] ^ x[46];
  assign t[86] = t[126] ^ x[43];
  assign t[87] = t[127] ^ x[44];
  assign t[88] = t[128] ^ x[45];
  assign t[89] = t[129] ^ x[51];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[130] ^ x[48];
  assign t[91] = t[131] ^ x[49];
  assign t[92] = t[132] ^ x[50];
  assign t[93] = (x[2]);
  assign t[94] = (x[2]);
  assign t[95] = (x[2]);
  assign t[96] = (x[2]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[7]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind265(x, y);
 input [51:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[7]);
  assign t[101] = (x[12]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[17]);
  assign t[106] = (x[17]);
  assign t[107] = (x[17]);
  assign t[108] = (x[17]);
  assign t[109] = (x[22]);
  assign t[10] = t[15] ^ t[16];
  assign t[110] = (x[22]);
  assign t[111] = (x[22]);
  assign t[112] = (x[22]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[32]);
  assign t[118] = (x[32]);
  assign t[119] = (x[32]);
  assign t[11] = t[24] ^ t[25];
  assign t[120] = (x[32]);
  assign t[121] = (x[37]);
  assign t[122] = (x[37]);
  assign t[123] = (x[37]);
  assign t[124] = (x[37]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[127] = (x[42]);
  assign t[128] = (x[42]);
  assign t[129] = (x[47]);
  assign t[12] = t[17] & t[18];
  assign t[130] = (x[47]);
  assign t[131] = (x[47]);
  assign t[132] = (x[47]);
  assign t[13] = t[26] ^ t[27];
  assign t[14] = t[19] & t[20];
  assign t[15] = t[28] ^ t[29];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[30] ^ t[17]);
  assign t[19] = ~(t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] ^ t[19]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[23]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = t[43] ^ x[6];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[21];
  assign t[37] = t[47] ^ x[26];
  assign t[38] = t[48] ^ x[31];
  assign t[39] = t[49] ^ x[36];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[41];
  assign t[41] = t[51] ^ x[46];
  assign t[42] = t[52] ^ x[51];
  assign t[43] = (~t[53] & t[54] & t[55] & t[56]) | (t[53] & ~t[55] & ~t[56]) | (t[53] & ~t[54] & ~t[56]) | (t[53] & ~t[54] & ~t[55]);
  assign t[44] = (~t[57] & t[58] & t[59] & t[60]) | (t[57] & ~t[59] & ~t[60]) | (t[57] & ~t[58] & ~t[60]) | (t[57] & ~t[58] & ~t[59]);
  assign t[45] = (~t[61] & t[62] & t[63] & t[64]) | (t[61] & ~t[63] & ~t[64]) | (t[61] & ~t[62] & ~t[64]) | (t[61] & ~t[62] & ~t[63]);
  assign t[46] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[47] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[48] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[49] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[51] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[52] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[53] = t[93] ^ x[6];
  assign t[54] = t[94] ^ x[3];
  assign t[55] = t[95] ^ x[4];
  assign t[56] = t[96] ^ x[5];
  assign t[57] = t[97] ^ x[11];
  assign t[58] = t[98] ^ x[8];
  assign t[59] = t[99] ^ x[9];
  assign t[5] = ~(t[8]);
  assign t[60] = t[100] ^ x[10];
  assign t[61] = t[101] ^ x[16];
  assign t[62] = t[102] ^ x[13];
  assign t[63] = t[103] ^ x[14];
  assign t[64] = t[104] ^ x[15];
  assign t[65] = t[105] ^ x[21];
  assign t[66] = t[106] ^ x[18];
  assign t[67] = t[107] ^ x[19];
  assign t[68] = t[108] ^ x[20];
  assign t[69] = t[109] ^ x[26];
  assign t[6] = ~(t[9]);
  assign t[70] = t[110] ^ x[23];
  assign t[71] = t[111] ^ x[24];
  assign t[72] = t[112] ^ x[25];
  assign t[73] = t[113] ^ x[31];
  assign t[74] = t[114] ^ x[28];
  assign t[75] = t[115] ^ x[29];
  assign t[76] = t[116] ^ x[30];
  assign t[77] = t[117] ^ x[36];
  assign t[78] = t[118] ^ x[33];
  assign t[79] = t[119] ^ x[34];
  assign t[7] = ~(t[10]);
  assign t[80] = t[120] ^ x[35];
  assign t[81] = t[121] ^ x[41];
  assign t[82] = t[122] ^ x[38];
  assign t[83] = t[123] ^ x[39];
  assign t[84] = t[124] ^ x[40];
  assign t[85] = t[125] ^ x[46];
  assign t[86] = t[126] ^ x[43];
  assign t[87] = t[127] ^ x[44];
  assign t[88] = t[128] ^ x[45];
  assign t[89] = t[129] ^ x[51];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[130] ^ x[48];
  assign t[91] = t[131] ^ x[49];
  assign t[92] = t[132] ^ x[50];
  assign t[93] = (x[2]);
  assign t[94] = (x[2]);
  assign t[95] = (x[2]);
  assign t[96] = (x[2]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[7]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind266(x, y);
 input [51:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[7]);
  assign t[101] = (x[12]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[17]);
  assign t[106] = (x[17]);
  assign t[107] = (x[17]);
  assign t[108] = (x[17]);
  assign t[109] = (x[22]);
  assign t[10] = t[15] ^ t[16];
  assign t[110] = (x[22]);
  assign t[111] = (x[22]);
  assign t[112] = (x[22]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[32]);
  assign t[118] = (x[32]);
  assign t[119] = (x[32]);
  assign t[11] = t[24] ^ t[25];
  assign t[120] = (x[32]);
  assign t[121] = (x[37]);
  assign t[122] = (x[37]);
  assign t[123] = (x[37]);
  assign t[124] = (x[37]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[127] = (x[42]);
  assign t[128] = (x[42]);
  assign t[129] = (x[47]);
  assign t[12] = t[17] & t[18];
  assign t[130] = (x[47]);
  assign t[131] = (x[47]);
  assign t[132] = (x[47]);
  assign t[13] = t[26] ^ t[27];
  assign t[14] = t[19] & t[20];
  assign t[15] = t[28] ^ t[29];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[30] ^ t[17]);
  assign t[19] = ~(t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] ^ t[19]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[23]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = t[43] ^ x[6];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[21];
  assign t[37] = t[47] ^ x[26];
  assign t[38] = t[48] ^ x[31];
  assign t[39] = t[49] ^ x[36];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[41];
  assign t[41] = t[51] ^ x[46];
  assign t[42] = t[52] ^ x[51];
  assign t[43] = (~t[53] & t[54] & t[55] & t[56]) | (t[53] & ~t[55] & ~t[56]) | (t[53] & ~t[54] & ~t[56]) | (t[53] & ~t[54] & ~t[55]);
  assign t[44] = (~t[57] & t[58] & t[59] & t[60]) | (t[57] & ~t[59] & ~t[60]) | (t[57] & ~t[58] & ~t[60]) | (t[57] & ~t[58] & ~t[59]);
  assign t[45] = (~t[61] & t[62] & t[63] & t[64]) | (t[61] & ~t[63] & ~t[64]) | (t[61] & ~t[62] & ~t[64]) | (t[61] & ~t[62] & ~t[63]);
  assign t[46] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[47] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[48] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[49] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[51] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[52] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[53] = t[93] ^ x[6];
  assign t[54] = t[94] ^ x[3];
  assign t[55] = t[95] ^ x[4];
  assign t[56] = t[96] ^ x[5];
  assign t[57] = t[97] ^ x[11];
  assign t[58] = t[98] ^ x[8];
  assign t[59] = t[99] ^ x[9];
  assign t[5] = ~(t[8]);
  assign t[60] = t[100] ^ x[10];
  assign t[61] = t[101] ^ x[16];
  assign t[62] = t[102] ^ x[13];
  assign t[63] = t[103] ^ x[14];
  assign t[64] = t[104] ^ x[15];
  assign t[65] = t[105] ^ x[21];
  assign t[66] = t[106] ^ x[18];
  assign t[67] = t[107] ^ x[19];
  assign t[68] = t[108] ^ x[20];
  assign t[69] = t[109] ^ x[26];
  assign t[6] = ~(t[9]);
  assign t[70] = t[110] ^ x[23];
  assign t[71] = t[111] ^ x[24];
  assign t[72] = t[112] ^ x[25];
  assign t[73] = t[113] ^ x[31];
  assign t[74] = t[114] ^ x[28];
  assign t[75] = t[115] ^ x[29];
  assign t[76] = t[116] ^ x[30];
  assign t[77] = t[117] ^ x[36];
  assign t[78] = t[118] ^ x[33];
  assign t[79] = t[119] ^ x[34];
  assign t[7] = ~(t[10]);
  assign t[80] = t[120] ^ x[35];
  assign t[81] = t[121] ^ x[41];
  assign t[82] = t[122] ^ x[38];
  assign t[83] = t[123] ^ x[39];
  assign t[84] = t[124] ^ x[40];
  assign t[85] = t[125] ^ x[46];
  assign t[86] = t[126] ^ x[43];
  assign t[87] = t[127] ^ x[44];
  assign t[88] = t[128] ^ x[45];
  assign t[89] = t[129] ^ x[51];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[130] ^ x[48];
  assign t[91] = t[131] ^ x[49];
  assign t[92] = t[132] ^ x[50];
  assign t[93] = (x[2]);
  assign t[94] = (x[2]);
  assign t[95] = (x[2]);
  assign t[96] = (x[2]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[7]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind267(x, y);
 input [51:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[7]);
  assign t[101] = (x[12]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[17]);
  assign t[106] = (x[17]);
  assign t[107] = (x[17]);
  assign t[108] = (x[17]);
  assign t[109] = (x[22]);
  assign t[10] = t[15] ^ t[16];
  assign t[110] = (x[22]);
  assign t[111] = (x[22]);
  assign t[112] = (x[22]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[32]);
  assign t[118] = (x[32]);
  assign t[119] = (x[32]);
  assign t[11] = t[24] ^ t[25];
  assign t[120] = (x[32]);
  assign t[121] = (x[37]);
  assign t[122] = (x[37]);
  assign t[123] = (x[37]);
  assign t[124] = (x[37]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[127] = (x[42]);
  assign t[128] = (x[42]);
  assign t[129] = (x[47]);
  assign t[12] = t[17] & t[18];
  assign t[130] = (x[47]);
  assign t[131] = (x[47]);
  assign t[132] = (x[47]);
  assign t[13] = t[26] ^ t[27];
  assign t[14] = t[19] & t[20];
  assign t[15] = t[28] ^ t[29];
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[30] ^ t[17]);
  assign t[19] = ~(t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] ^ t[19]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[32] ^ t[21]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[23]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = t[43] ^ x[6];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[21];
  assign t[37] = t[47] ^ x[26];
  assign t[38] = t[48] ^ x[31];
  assign t[39] = t[49] ^ x[36];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[41];
  assign t[41] = t[51] ^ x[46];
  assign t[42] = t[52] ^ x[51];
  assign t[43] = (~t[53] & t[54] & t[55] & t[56]) | (t[53] & ~t[55] & ~t[56]) | (t[53] & ~t[54] & ~t[56]) | (t[53] & ~t[54] & ~t[55]);
  assign t[44] = (~t[57] & t[58] & t[59] & t[60]) | (t[57] & ~t[59] & ~t[60]) | (t[57] & ~t[58] & ~t[60]) | (t[57] & ~t[58] & ~t[59]);
  assign t[45] = (~t[61] & t[62] & t[63] & t[64]) | (t[61] & ~t[63] & ~t[64]) | (t[61] & ~t[62] & ~t[64]) | (t[61] & ~t[62] & ~t[63]);
  assign t[46] = (~t[65] & t[66] & t[67] & t[68]) | (t[65] & ~t[67] & ~t[68]) | (t[65] & ~t[66] & ~t[68]) | (t[65] & ~t[66] & ~t[67]);
  assign t[47] = (~t[69] & t[70] & t[71] & t[72]) | (t[69] & ~t[71] & ~t[72]) | (t[69] & ~t[70] & ~t[72]) | (t[69] & ~t[70] & ~t[71]);
  assign t[48] = (~t[73] & t[74] & t[75] & t[76]) | (t[73] & ~t[75] & ~t[76]) | (t[73] & ~t[74] & ~t[76]) | (t[73] & ~t[74] & ~t[75]);
  assign t[49] = (~t[77] & t[78] & t[79] & t[80]) | (t[77] & ~t[79] & ~t[80]) | (t[77] & ~t[78] & ~t[80]) | (t[77] & ~t[78] & ~t[79]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[81] & t[82] & t[83] & t[84]) | (t[81] & ~t[83] & ~t[84]) | (t[81] & ~t[82] & ~t[84]) | (t[81] & ~t[82] & ~t[83]);
  assign t[51] = (~t[85] & t[86] & t[87] & t[88]) | (t[85] & ~t[87] & ~t[88]) | (t[85] & ~t[86] & ~t[88]) | (t[85] & ~t[86] & ~t[87]);
  assign t[52] = (~t[89] & t[90] & t[91] & t[92]) | (t[89] & ~t[91] & ~t[92]) | (t[89] & ~t[90] & ~t[92]) | (t[89] & ~t[90] & ~t[91]);
  assign t[53] = t[93] ^ x[6];
  assign t[54] = t[94] ^ x[3];
  assign t[55] = t[95] ^ x[4];
  assign t[56] = t[96] ^ x[5];
  assign t[57] = t[97] ^ x[11];
  assign t[58] = t[98] ^ x[8];
  assign t[59] = t[99] ^ x[9];
  assign t[5] = ~(t[8]);
  assign t[60] = t[100] ^ x[10];
  assign t[61] = t[101] ^ x[16];
  assign t[62] = t[102] ^ x[13];
  assign t[63] = t[103] ^ x[14];
  assign t[64] = t[104] ^ x[15];
  assign t[65] = t[105] ^ x[21];
  assign t[66] = t[106] ^ x[18];
  assign t[67] = t[107] ^ x[19];
  assign t[68] = t[108] ^ x[20];
  assign t[69] = t[109] ^ x[26];
  assign t[6] = ~(t[9]);
  assign t[70] = t[110] ^ x[23];
  assign t[71] = t[111] ^ x[24];
  assign t[72] = t[112] ^ x[25];
  assign t[73] = t[113] ^ x[31];
  assign t[74] = t[114] ^ x[28];
  assign t[75] = t[115] ^ x[29];
  assign t[76] = t[116] ^ x[30];
  assign t[77] = t[117] ^ x[36];
  assign t[78] = t[118] ^ x[33];
  assign t[79] = t[119] ^ x[34];
  assign t[7] = ~(t[10]);
  assign t[80] = t[120] ^ x[35];
  assign t[81] = t[121] ^ x[41];
  assign t[82] = t[122] ^ x[38];
  assign t[83] = t[123] ^ x[39];
  assign t[84] = t[124] ^ x[40];
  assign t[85] = t[125] ^ x[46];
  assign t[86] = t[126] ^ x[43];
  assign t[87] = t[127] ^ x[44];
  assign t[88] = t[128] ^ x[45];
  assign t[89] = t[129] ^ x[51];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[130] ^ x[48];
  assign t[91] = t[131] ^ x[49];
  assign t[92] = t[132] ^ x[50];
  assign t[93] = (x[2]);
  assign t[94] = (x[2]);
  assign t[95] = (x[2]);
  assign t[96] = (x[2]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[7]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind268(x, y);
 input [66:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[34];
  assign t[101] = t[153] ^ x[35];
  assign t[102] = t[154] ^ x[41];
  assign t[103] = t[155] ^ x[38];
  assign t[104] = t[156] ^ x[39];
  assign t[105] = t[157] ^ x[40];
  assign t[106] = t[158] ^ x[46];
  assign t[107] = t[159] ^ x[43];
  assign t[108] = t[160] ^ x[44];
  assign t[109] = t[161] ^ x[45];
  assign t[10] = t[15] ^ t[16];
  assign t[110] = t[162] ^ x[51];
  assign t[111] = t[163] ^ x[48];
  assign t[112] = t[164] ^ x[49];
  assign t[113] = t[165] ^ x[50];
  assign t[114] = t[166] ^ x[56];
  assign t[115] = t[167] ^ x[53];
  assign t[116] = t[168] ^ x[54];
  assign t[117] = t[169] ^ x[55];
  assign t[118] = t[170] ^ x[61];
  assign t[119] = t[171] ^ x[58];
  assign t[11] = t[17] ^ t[18];
  assign t[120] = t[172] ^ x[59];
  assign t[121] = t[173] ^ x[60];
  assign t[122] = t[174] ^ x[66];
  assign t[123] = t[175] ^ x[63];
  assign t[124] = t[176] ^ x[64];
  assign t[125] = t[177] ^ x[65];
  assign t[126] = (x[2]);
  assign t[127] = (x[2]);
  assign t[128] = (x[2]);
  assign t[129] = (x[2]);
  assign t[12] = t[19] & t[20];
  assign t[130] = (x[7]);
  assign t[131] = (x[7]);
  assign t[132] = (x[7]);
  assign t[133] = (x[7]);
  assign t[134] = (x[12]);
  assign t[135] = (x[12]);
  assign t[136] = (x[12]);
  assign t[137] = (x[12]);
  assign t[138] = (x[17]);
  assign t[139] = (x[17]);
  assign t[13] = t[21] ^ t[22];
  assign t[140] = (x[17]);
  assign t[141] = (x[17]);
  assign t[142] = (x[22]);
  assign t[143] = (x[22]);
  assign t[144] = (x[22]);
  assign t[145] = (x[22]);
  assign t[146] = (x[27]);
  assign t[147] = (x[27]);
  assign t[148] = (x[27]);
  assign t[149] = (x[27]);
  assign t[14] = t[23] & t[24];
  assign t[150] = (x[32]);
  assign t[151] = (x[32]);
  assign t[152] = (x[32]);
  assign t[153] = (x[32]);
  assign t[154] = (x[37]);
  assign t[155] = (x[37]);
  assign t[156] = (x[37]);
  assign t[157] = (x[37]);
  assign t[158] = (x[42]);
  assign t[159] = (x[42]);
  assign t[15] = t[25] ^ t[26];
  assign t[160] = (x[42]);
  assign t[161] = (x[42]);
  assign t[162] = (x[47]);
  assign t[163] = (x[47]);
  assign t[164] = (x[47]);
  assign t[165] = (x[47]);
  assign t[166] = (x[52]);
  assign t[167] = (x[52]);
  assign t[168] = (x[52]);
  assign t[169] = (x[52]);
  assign t[16] = t[27] & t[28];
  assign t[170] = (x[57]);
  assign t[171] = (x[57]);
  assign t[172] = (x[57]);
  assign t[173] = (x[57]);
  assign t[174] = (x[62]);
  assign t[175] = (x[62]);
  assign t[176] = (x[62]);
  assign t[177] = (x[62]);
  assign t[17] = t[36] ^ t[37];
  assign t[18] = t[19] & t[29];
  assign t[19] = ~(t[37]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[38] ^ t[19]);
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[23] & t[30];
  assign t[23] = ~(t[40]);
  assign t[24] = ~(t[41] ^ t[23]);
  assign t[25] = t[42] ^ t[43];
  assign t[26] = t[27] & t[31];
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[44] ^ t[27]);
  assign t[29] = t[38] ^ t[32];
  assign t[2] = ~(t[4] ^ t[35]);
  assign t[30] = t[41] ^ t[33];
  assign t[31] = t[44] ^ t[34];
  assign t[32] = t[37] ^ t[45];
  assign t[33] = t[40] ^ t[46];
  assign t[34] = t[43] ^ t[47];
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = t[61] ^ x[6];
  assign t[49] = t[62] ^ x[11];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ x[16];
  assign t[51] = t[64] ^ x[21];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[31];
  assign t[54] = t[67] ^ x[36];
  assign t[55] = t[68] ^ x[41];
  assign t[56] = t[69] ^ x[46];
  assign t[57] = t[70] ^ x[51];
  assign t[58] = t[71] ^ x[56];
  assign t[59] = t[72] ^ x[61];
  assign t[5] = ~(t[8]);
  assign t[60] = t[73] ^ x[66];
  assign t[61] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[62] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[63] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[64] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[65] = (~t[90] & t[91] & t[92] & t[93]) | (t[90] & ~t[92] & ~t[93]) | (t[90] & ~t[91] & ~t[93]) | (t[90] & ~t[91] & ~t[92]);
  assign t[66] = (~t[94] & t[95] & t[96] & t[97]) | (t[94] & ~t[96] & ~t[97]) | (t[94] & ~t[95] & ~t[97]) | (t[94] & ~t[95] & ~t[96]);
  assign t[67] = (~t[98] & t[99] & t[100] & t[101]) | (t[98] & ~t[100] & ~t[101]) | (t[98] & ~t[99] & ~t[101]) | (t[98] & ~t[99] & ~t[100]);
  assign t[68] = (~t[102] & t[103] & t[104] & t[105]) | (t[102] & ~t[104] & ~t[105]) | (t[102] & ~t[103] & ~t[105]) | (t[102] & ~t[103] & ~t[104]);
  assign t[69] = (~t[106] & t[107] & t[108] & t[109]) | (t[106] & ~t[108] & ~t[109]) | (t[106] & ~t[107] & ~t[109]) | (t[106] & ~t[107] & ~t[108]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[110] & t[111] & t[112] & t[113]) | (t[110] & ~t[112] & ~t[113]) | (t[110] & ~t[111] & ~t[113]) | (t[110] & ~t[111] & ~t[112]);
  assign t[71] = (~t[114] & t[115] & t[116] & t[117]) | (t[114] & ~t[116] & ~t[117]) | (t[114] & ~t[115] & ~t[117]) | (t[114] & ~t[115] & ~t[116]);
  assign t[72] = (~t[118] & t[119] & t[120] & t[121]) | (t[118] & ~t[120] & ~t[121]) | (t[118] & ~t[119] & ~t[121]) | (t[118] & ~t[119] & ~t[120]);
  assign t[73] = (~t[122] & t[123] & t[124] & t[125]) | (t[122] & ~t[124] & ~t[125]) | (t[122] & ~t[123] & ~t[125]) | (t[122] & ~t[123] & ~t[124]);
  assign t[74] = t[126] ^ x[6];
  assign t[75] = t[127] ^ x[3];
  assign t[76] = t[128] ^ x[4];
  assign t[77] = t[129] ^ x[5];
  assign t[78] = t[130] ^ x[11];
  assign t[79] = t[131] ^ x[8];
  assign t[7] = ~(t[10]);
  assign t[80] = t[132] ^ x[9];
  assign t[81] = t[133] ^ x[10];
  assign t[82] = t[134] ^ x[16];
  assign t[83] = t[135] ^ x[13];
  assign t[84] = t[136] ^ x[14];
  assign t[85] = t[137] ^ x[15];
  assign t[86] = t[138] ^ x[21];
  assign t[87] = t[139] ^ x[18];
  assign t[88] = t[140] ^ x[19];
  assign t[89] = t[141] ^ x[20];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[142] ^ x[26];
  assign t[91] = t[143] ^ x[23];
  assign t[92] = t[144] ^ x[24];
  assign t[93] = t[145] ^ x[25];
  assign t[94] = t[146] ^ x[31];
  assign t[95] = t[147] ^ x[28];
  assign t[96] = t[148] ^ x[29];
  assign t[97] = t[149] ^ x[30];
  assign t[98] = t[150] ^ x[36];
  assign t[99] = t[151] ^ x[33];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind269(x, y);
 input [66:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[34];
  assign t[101] = t[153] ^ x[35];
  assign t[102] = t[154] ^ x[41];
  assign t[103] = t[155] ^ x[38];
  assign t[104] = t[156] ^ x[39];
  assign t[105] = t[157] ^ x[40];
  assign t[106] = t[158] ^ x[46];
  assign t[107] = t[159] ^ x[43];
  assign t[108] = t[160] ^ x[44];
  assign t[109] = t[161] ^ x[45];
  assign t[10] = t[15] ^ t[16];
  assign t[110] = t[162] ^ x[51];
  assign t[111] = t[163] ^ x[48];
  assign t[112] = t[164] ^ x[49];
  assign t[113] = t[165] ^ x[50];
  assign t[114] = t[166] ^ x[56];
  assign t[115] = t[167] ^ x[53];
  assign t[116] = t[168] ^ x[54];
  assign t[117] = t[169] ^ x[55];
  assign t[118] = t[170] ^ x[61];
  assign t[119] = t[171] ^ x[58];
  assign t[11] = t[17] ^ t[18];
  assign t[120] = t[172] ^ x[59];
  assign t[121] = t[173] ^ x[60];
  assign t[122] = t[174] ^ x[66];
  assign t[123] = t[175] ^ x[63];
  assign t[124] = t[176] ^ x[64];
  assign t[125] = t[177] ^ x[65];
  assign t[126] = (x[2]);
  assign t[127] = (x[2]);
  assign t[128] = (x[2]);
  assign t[129] = (x[2]);
  assign t[12] = t[19] & t[20];
  assign t[130] = (x[7]);
  assign t[131] = (x[7]);
  assign t[132] = (x[7]);
  assign t[133] = (x[7]);
  assign t[134] = (x[12]);
  assign t[135] = (x[12]);
  assign t[136] = (x[12]);
  assign t[137] = (x[12]);
  assign t[138] = (x[17]);
  assign t[139] = (x[17]);
  assign t[13] = t[21] ^ t[22];
  assign t[140] = (x[17]);
  assign t[141] = (x[17]);
  assign t[142] = (x[22]);
  assign t[143] = (x[22]);
  assign t[144] = (x[22]);
  assign t[145] = (x[22]);
  assign t[146] = (x[27]);
  assign t[147] = (x[27]);
  assign t[148] = (x[27]);
  assign t[149] = (x[27]);
  assign t[14] = t[23] & t[24];
  assign t[150] = (x[32]);
  assign t[151] = (x[32]);
  assign t[152] = (x[32]);
  assign t[153] = (x[32]);
  assign t[154] = (x[37]);
  assign t[155] = (x[37]);
  assign t[156] = (x[37]);
  assign t[157] = (x[37]);
  assign t[158] = (x[42]);
  assign t[159] = (x[42]);
  assign t[15] = t[25] ^ t[26];
  assign t[160] = (x[42]);
  assign t[161] = (x[42]);
  assign t[162] = (x[47]);
  assign t[163] = (x[47]);
  assign t[164] = (x[47]);
  assign t[165] = (x[47]);
  assign t[166] = (x[52]);
  assign t[167] = (x[52]);
  assign t[168] = (x[52]);
  assign t[169] = (x[52]);
  assign t[16] = t[27] & t[28];
  assign t[170] = (x[57]);
  assign t[171] = (x[57]);
  assign t[172] = (x[57]);
  assign t[173] = (x[57]);
  assign t[174] = (x[62]);
  assign t[175] = (x[62]);
  assign t[176] = (x[62]);
  assign t[177] = (x[62]);
  assign t[17] = t[36] ^ t[37];
  assign t[18] = t[19] & t[29];
  assign t[19] = ~(t[37]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[38] ^ t[19]);
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[23] & t[30];
  assign t[23] = ~(t[40]);
  assign t[24] = ~(t[41] ^ t[23]);
  assign t[25] = t[42] ^ t[43];
  assign t[26] = t[27] & t[31];
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[44] ^ t[27]);
  assign t[29] = t[38] ^ t[32];
  assign t[2] = ~(t[4] ^ t[35]);
  assign t[30] = t[41] ^ t[33];
  assign t[31] = t[44] ^ t[34];
  assign t[32] = t[37] ^ t[45];
  assign t[33] = t[40] ^ t[46];
  assign t[34] = t[43] ^ t[47];
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = t[61] ^ x[6];
  assign t[49] = t[62] ^ x[11];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ x[16];
  assign t[51] = t[64] ^ x[21];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[31];
  assign t[54] = t[67] ^ x[36];
  assign t[55] = t[68] ^ x[41];
  assign t[56] = t[69] ^ x[46];
  assign t[57] = t[70] ^ x[51];
  assign t[58] = t[71] ^ x[56];
  assign t[59] = t[72] ^ x[61];
  assign t[5] = ~(t[8]);
  assign t[60] = t[73] ^ x[66];
  assign t[61] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[62] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[63] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[64] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[65] = (~t[90] & t[91] & t[92] & t[93]) | (t[90] & ~t[92] & ~t[93]) | (t[90] & ~t[91] & ~t[93]) | (t[90] & ~t[91] & ~t[92]);
  assign t[66] = (~t[94] & t[95] & t[96] & t[97]) | (t[94] & ~t[96] & ~t[97]) | (t[94] & ~t[95] & ~t[97]) | (t[94] & ~t[95] & ~t[96]);
  assign t[67] = (~t[98] & t[99] & t[100] & t[101]) | (t[98] & ~t[100] & ~t[101]) | (t[98] & ~t[99] & ~t[101]) | (t[98] & ~t[99] & ~t[100]);
  assign t[68] = (~t[102] & t[103] & t[104] & t[105]) | (t[102] & ~t[104] & ~t[105]) | (t[102] & ~t[103] & ~t[105]) | (t[102] & ~t[103] & ~t[104]);
  assign t[69] = (~t[106] & t[107] & t[108] & t[109]) | (t[106] & ~t[108] & ~t[109]) | (t[106] & ~t[107] & ~t[109]) | (t[106] & ~t[107] & ~t[108]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[110] & t[111] & t[112] & t[113]) | (t[110] & ~t[112] & ~t[113]) | (t[110] & ~t[111] & ~t[113]) | (t[110] & ~t[111] & ~t[112]);
  assign t[71] = (~t[114] & t[115] & t[116] & t[117]) | (t[114] & ~t[116] & ~t[117]) | (t[114] & ~t[115] & ~t[117]) | (t[114] & ~t[115] & ~t[116]);
  assign t[72] = (~t[118] & t[119] & t[120] & t[121]) | (t[118] & ~t[120] & ~t[121]) | (t[118] & ~t[119] & ~t[121]) | (t[118] & ~t[119] & ~t[120]);
  assign t[73] = (~t[122] & t[123] & t[124] & t[125]) | (t[122] & ~t[124] & ~t[125]) | (t[122] & ~t[123] & ~t[125]) | (t[122] & ~t[123] & ~t[124]);
  assign t[74] = t[126] ^ x[6];
  assign t[75] = t[127] ^ x[3];
  assign t[76] = t[128] ^ x[4];
  assign t[77] = t[129] ^ x[5];
  assign t[78] = t[130] ^ x[11];
  assign t[79] = t[131] ^ x[8];
  assign t[7] = ~(t[10]);
  assign t[80] = t[132] ^ x[9];
  assign t[81] = t[133] ^ x[10];
  assign t[82] = t[134] ^ x[16];
  assign t[83] = t[135] ^ x[13];
  assign t[84] = t[136] ^ x[14];
  assign t[85] = t[137] ^ x[15];
  assign t[86] = t[138] ^ x[21];
  assign t[87] = t[139] ^ x[18];
  assign t[88] = t[140] ^ x[19];
  assign t[89] = t[141] ^ x[20];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[142] ^ x[26];
  assign t[91] = t[143] ^ x[23];
  assign t[92] = t[144] ^ x[24];
  assign t[93] = t[145] ^ x[25];
  assign t[94] = t[146] ^ x[31];
  assign t[95] = t[147] ^ x[28];
  assign t[96] = t[148] ^ x[29];
  assign t[97] = t[149] ^ x[30];
  assign t[98] = t[150] ^ x[36];
  assign t[99] = t[151] ^ x[33];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind270(x, y);
 input [66:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[34];
  assign t[101] = t[153] ^ x[35];
  assign t[102] = t[154] ^ x[41];
  assign t[103] = t[155] ^ x[38];
  assign t[104] = t[156] ^ x[39];
  assign t[105] = t[157] ^ x[40];
  assign t[106] = t[158] ^ x[46];
  assign t[107] = t[159] ^ x[43];
  assign t[108] = t[160] ^ x[44];
  assign t[109] = t[161] ^ x[45];
  assign t[10] = t[15] ^ t[16];
  assign t[110] = t[162] ^ x[51];
  assign t[111] = t[163] ^ x[48];
  assign t[112] = t[164] ^ x[49];
  assign t[113] = t[165] ^ x[50];
  assign t[114] = t[166] ^ x[56];
  assign t[115] = t[167] ^ x[53];
  assign t[116] = t[168] ^ x[54];
  assign t[117] = t[169] ^ x[55];
  assign t[118] = t[170] ^ x[61];
  assign t[119] = t[171] ^ x[58];
  assign t[11] = t[17] ^ t[18];
  assign t[120] = t[172] ^ x[59];
  assign t[121] = t[173] ^ x[60];
  assign t[122] = t[174] ^ x[66];
  assign t[123] = t[175] ^ x[63];
  assign t[124] = t[176] ^ x[64];
  assign t[125] = t[177] ^ x[65];
  assign t[126] = (x[2]);
  assign t[127] = (x[2]);
  assign t[128] = (x[2]);
  assign t[129] = (x[2]);
  assign t[12] = t[19] & t[20];
  assign t[130] = (x[7]);
  assign t[131] = (x[7]);
  assign t[132] = (x[7]);
  assign t[133] = (x[7]);
  assign t[134] = (x[12]);
  assign t[135] = (x[12]);
  assign t[136] = (x[12]);
  assign t[137] = (x[12]);
  assign t[138] = (x[17]);
  assign t[139] = (x[17]);
  assign t[13] = t[21] ^ t[22];
  assign t[140] = (x[17]);
  assign t[141] = (x[17]);
  assign t[142] = (x[22]);
  assign t[143] = (x[22]);
  assign t[144] = (x[22]);
  assign t[145] = (x[22]);
  assign t[146] = (x[27]);
  assign t[147] = (x[27]);
  assign t[148] = (x[27]);
  assign t[149] = (x[27]);
  assign t[14] = t[23] & t[24];
  assign t[150] = (x[32]);
  assign t[151] = (x[32]);
  assign t[152] = (x[32]);
  assign t[153] = (x[32]);
  assign t[154] = (x[37]);
  assign t[155] = (x[37]);
  assign t[156] = (x[37]);
  assign t[157] = (x[37]);
  assign t[158] = (x[42]);
  assign t[159] = (x[42]);
  assign t[15] = t[25] ^ t[26];
  assign t[160] = (x[42]);
  assign t[161] = (x[42]);
  assign t[162] = (x[47]);
  assign t[163] = (x[47]);
  assign t[164] = (x[47]);
  assign t[165] = (x[47]);
  assign t[166] = (x[52]);
  assign t[167] = (x[52]);
  assign t[168] = (x[52]);
  assign t[169] = (x[52]);
  assign t[16] = t[27] & t[28];
  assign t[170] = (x[57]);
  assign t[171] = (x[57]);
  assign t[172] = (x[57]);
  assign t[173] = (x[57]);
  assign t[174] = (x[62]);
  assign t[175] = (x[62]);
  assign t[176] = (x[62]);
  assign t[177] = (x[62]);
  assign t[17] = t[36] ^ t[37];
  assign t[18] = t[19] & t[29];
  assign t[19] = ~(t[37]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[38] ^ t[19]);
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[23] & t[30];
  assign t[23] = ~(t[40]);
  assign t[24] = ~(t[41] ^ t[23]);
  assign t[25] = t[42] ^ t[43];
  assign t[26] = t[27] & t[31];
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[44] ^ t[27]);
  assign t[29] = t[38] ^ t[32];
  assign t[2] = ~(t[4] ^ t[35]);
  assign t[30] = t[41] ^ t[33];
  assign t[31] = t[44] ^ t[34];
  assign t[32] = t[37] ^ t[45];
  assign t[33] = t[40] ^ t[46];
  assign t[34] = t[43] ^ t[47];
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = t[61] ^ x[6];
  assign t[49] = t[62] ^ x[11];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ x[16];
  assign t[51] = t[64] ^ x[21];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[31];
  assign t[54] = t[67] ^ x[36];
  assign t[55] = t[68] ^ x[41];
  assign t[56] = t[69] ^ x[46];
  assign t[57] = t[70] ^ x[51];
  assign t[58] = t[71] ^ x[56];
  assign t[59] = t[72] ^ x[61];
  assign t[5] = ~(t[8]);
  assign t[60] = t[73] ^ x[66];
  assign t[61] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[62] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[63] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[64] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[65] = (~t[90] & t[91] & t[92] & t[93]) | (t[90] & ~t[92] & ~t[93]) | (t[90] & ~t[91] & ~t[93]) | (t[90] & ~t[91] & ~t[92]);
  assign t[66] = (~t[94] & t[95] & t[96] & t[97]) | (t[94] & ~t[96] & ~t[97]) | (t[94] & ~t[95] & ~t[97]) | (t[94] & ~t[95] & ~t[96]);
  assign t[67] = (~t[98] & t[99] & t[100] & t[101]) | (t[98] & ~t[100] & ~t[101]) | (t[98] & ~t[99] & ~t[101]) | (t[98] & ~t[99] & ~t[100]);
  assign t[68] = (~t[102] & t[103] & t[104] & t[105]) | (t[102] & ~t[104] & ~t[105]) | (t[102] & ~t[103] & ~t[105]) | (t[102] & ~t[103] & ~t[104]);
  assign t[69] = (~t[106] & t[107] & t[108] & t[109]) | (t[106] & ~t[108] & ~t[109]) | (t[106] & ~t[107] & ~t[109]) | (t[106] & ~t[107] & ~t[108]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[110] & t[111] & t[112] & t[113]) | (t[110] & ~t[112] & ~t[113]) | (t[110] & ~t[111] & ~t[113]) | (t[110] & ~t[111] & ~t[112]);
  assign t[71] = (~t[114] & t[115] & t[116] & t[117]) | (t[114] & ~t[116] & ~t[117]) | (t[114] & ~t[115] & ~t[117]) | (t[114] & ~t[115] & ~t[116]);
  assign t[72] = (~t[118] & t[119] & t[120] & t[121]) | (t[118] & ~t[120] & ~t[121]) | (t[118] & ~t[119] & ~t[121]) | (t[118] & ~t[119] & ~t[120]);
  assign t[73] = (~t[122] & t[123] & t[124] & t[125]) | (t[122] & ~t[124] & ~t[125]) | (t[122] & ~t[123] & ~t[125]) | (t[122] & ~t[123] & ~t[124]);
  assign t[74] = t[126] ^ x[6];
  assign t[75] = t[127] ^ x[3];
  assign t[76] = t[128] ^ x[4];
  assign t[77] = t[129] ^ x[5];
  assign t[78] = t[130] ^ x[11];
  assign t[79] = t[131] ^ x[8];
  assign t[7] = ~(t[10]);
  assign t[80] = t[132] ^ x[9];
  assign t[81] = t[133] ^ x[10];
  assign t[82] = t[134] ^ x[16];
  assign t[83] = t[135] ^ x[13];
  assign t[84] = t[136] ^ x[14];
  assign t[85] = t[137] ^ x[15];
  assign t[86] = t[138] ^ x[21];
  assign t[87] = t[139] ^ x[18];
  assign t[88] = t[140] ^ x[19];
  assign t[89] = t[141] ^ x[20];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[142] ^ x[26];
  assign t[91] = t[143] ^ x[23];
  assign t[92] = t[144] ^ x[24];
  assign t[93] = t[145] ^ x[25];
  assign t[94] = t[146] ^ x[31];
  assign t[95] = t[147] ^ x[28];
  assign t[96] = t[148] ^ x[29];
  assign t[97] = t[149] ^ x[30];
  assign t[98] = t[150] ^ x[36];
  assign t[99] = t[151] ^ x[33];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind271(x, y);
 input [66:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[152] ^ x[34];
  assign t[101] = t[153] ^ x[35];
  assign t[102] = t[154] ^ x[41];
  assign t[103] = t[155] ^ x[38];
  assign t[104] = t[156] ^ x[39];
  assign t[105] = t[157] ^ x[40];
  assign t[106] = t[158] ^ x[46];
  assign t[107] = t[159] ^ x[43];
  assign t[108] = t[160] ^ x[44];
  assign t[109] = t[161] ^ x[45];
  assign t[10] = t[15] ^ t[16];
  assign t[110] = t[162] ^ x[51];
  assign t[111] = t[163] ^ x[48];
  assign t[112] = t[164] ^ x[49];
  assign t[113] = t[165] ^ x[50];
  assign t[114] = t[166] ^ x[56];
  assign t[115] = t[167] ^ x[53];
  assign t[116] = t[168] ^ x[54];
  assign t[117] = t[169] ^ x[55];
  assign t[118] = t[170] ^ x[61];
  assign t[119] = t[171] ^ x[58];
  assign t[11] = t[17] ^ t[18];
  assign t[120] = t[172] ^ x[59];
  assign t[121] = t[173] ^ x[60];
  assign t[122] = t[174] ^ x[66];
  assign t[123] = t[175] ^ x[63];
  assign t[124] = t[176] ^ x[64];
  assign t[125] = t[177] ^ x[65];
  assign t[126] = (x[2]);
  assign t[127] = (x[2]);
  assign t[128] = (x[2]);
  assign t[129] = (x[2]);
  assign t[12] = t[19] & t[20];
  assign t[130] = (x[7]);
  assign t[131] = (x[7]);
  assign t[132] = (x[7]);
  assign t[133] = (x[7]);
  assign t[134] = (x[12]);
  assign t[135] = (x[12]);
  assign t[136] = (x[12]);
  assign t[137] = (x[12]);
  assign t[138] = (x[17]);
  assign t[139] = (x[17]);
  assign t[13] = t[21] ^ t[22];
  assign t[140] = (x[17]);
  assign t[141] = (x[17]);
  assign t[142] = (x[22]);
  assign t[143] = (x[22]);
  assign t[144] = (x[22]);
  assign t[145] = (x[22]);
  assign t[146] = (x[27]);
  assign t[147] = (x[27]);
  assign t[148] = (x[27]);
  assign t[149] = (x[27]);
  assign t[14] = t[23] & t[24];
  assign t[150] = (x[32]);
  assign t[151] = (x[32]);
  assign t[152] = (x[32]);
  assign t[153] = (x[32]);
  assign t[154] = (x[37]);
  assign t[155] = (x[37]);
  assign t[156] = (x[37]);
  assign t[157] = (x[37]);
  assign t[158] = (x[42]);
  assign t[159] = (x[42]);
  assign t[15] = t[25] ^ t[26];
  assign t[160] = (x[42]);
  assign t[161] = (x[42]);
  assign t[162] = (x[47]);
  assign t[163] = (x[47]);
  assign t[164] = (x[47]);
  assign t[165] = (x[47]);
  assign t[166] = (x[52]);
  assign t[167] = (x[52]);
  assign t[168] = (x[52]);
  assign t[169] = (x[52]);
  assign t[16] = t[27] & t[28];
  assign t[170] = (x[57]);
  assign t[171] = (x[57]);
  assign t[172] = (x[57]);
  assign t[173] = (x[57]);
  assign t[174] = (x[62]);
  assign t[175] = (x[62]);
  assign t[176] = (x[62]);
  assign t[177] = (x[62]);
  assign t[17] = t[36] ^ t[37];
  assign t[18] = t[19] & t[29];
  assign t[19] = ~(t[37]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[38] ^ t[19]);
  assign t[21] = t[39] ^ t[40];
  assign t[22] = t[23] & t[30];
  assign t[23] = ~(t[40]);
  assign t[24] = ~(t[41] ^ t[23]);
  assign t[25] = t[42] ^ t[43];
  assign t[26] = t[27] & t[31];
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[44] ^ t[27]);
  assign t[29] = t[38] ^ t[32];
  assign t[2] = ~(t[4] ^ t[35]);
  assign t[30] = t[41] ^ t[33];
  assign t[31] = t[44] ^ t[34];
  assign t[32] = t[37] ^ t[45];
  assign t[33] = t[40] ^ t[46];
  assign t[34] = t[43] ^ t[47];
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = t[61] ^ x[6];
  assign t[49] = t[62] ^ x[11];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ x[16];
  assign t[51] = t[64] ^ x[21];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[31];
  assign t[54] = t[67] ^ x[36];
  assign t[55] = t[68] ^ x[41];
  assign t[56] = t[69] ^ x[46];
  assign t[57] = t[70] ^ x[51];
  assign t[58] = t[71] ^ x[56];
  assign t[59] = t[72] ^ x[61];
  assign t[5] = ~(t[8]);
  assign t[60] = t[73] ^ x[66];
  assign t[61] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[62] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[63] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[64] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[65] = (~t[90] & t[91] & t[92] & t[93]) | (t[90] & ~t[92] & ~t[93]) | (t[90] & ~t[91] & ~t[93]) | (t[90] & ~t[91] & ~t[92]);
  assign t[66] = (~t[94] & t[95] & t[96] & t[97]) | (t[94] & ~t[96] & ~t[97]) | (t[94] & ~t[95] & ~t[97]) | (t[94] & ~t[95] & ~t[96]);
  assign t[67] = (~t[98] & t[99] & t[100] & t[101]) | (t[98] & ~t[100] & ~t[101]) | (t[98] & ~t[99] & ~t[101]) | (t[98] & ~t[99] & ~t[100]);
  assign t[68] = (~t[102] & t[103] & t[104] & t[105]) | (t[102] & ~t[104] & ~t[105]) | (t[102] & ~t[103] & ~t[105]) | (t[102] & ~t[103] & ~t[104]);
  assign t[69] = (~t[106] & t[107] & t[108] & t[109]) | (t[106] & ~t[108] & ~t[109]) | (t[106] & ~t[107] & ~t[109]) | (t[106] & ~t[107] & ~t[108]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[110] & t[111] & t[112] & t[113]) | (t[110] & ~t[112] & ~t[113]) | (t[110] & ~t[111] & ~t[113]) | (t[110] & ~t[111] & ~t[112]);
  assign t[71] = (~t[114] & t[115] & t[116] & t[117]) | (t[114] & ~t[116] & ~t[117]) | (t[114] & ~t[115] & ~t[117]) | (t[114] & ~t[115] & ~t[116]);
  assign t[72] = (~t[118] & t[119] & t[120] & t[121]) | (t[118] & ~t[120] & ~t[121]) | (t[118] & ~t[119] & ~t[121]) | (t[118] & ~t[119] & ~t[120]);
  assign t[73] = (~t[122] & t[123] & t[124] & t[125]) | (t[122] & ~t[124] & ~t[125]) | (t[122] & ~t[123] & ~t[125]) | (t[122] & ~t[123] & ~t[124]);
  assign t[74] = t[126] ^ x[6];
  assign t[75] = t[127] ^ x[3];
  assign t[76] = t[128] ^ x[4];
  assign t[77] = t[129] ^ x[5];
  assign t[78] = t[130] ^ x[11];
  assign t[79] = t[131] ^ x[8];
  assign t[7] = ~(t[10]);
  assign t[80] = t[132] ^ x[9];
  assign t[81] = t[133] ^ x[10];
  assign t[82] = t[134] ^ x[16];
  assign t[83] = t[135] ^ x[13];
  assign t[84] = t[136] ^ x[14];
  assign t[85] = t[137] ^ x[15];
  assign t[86] = t[138] ^ x[21];
  assign t[87] = t[139] ^ x[18];
  assign t[88] = t[140] ^ x[19];
  assign t[89] = t[141] ^ x[20];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[142] ^ x[26];
  assign t[91] = t[143] ^ x[23];
  assign t[92] = t[144] ^ x[24];
  assign t[93] = t[145] ^ x[25];
  assign t[94] = t[146] ^ x[31];
  assign t[95] = t[147] ^ x[28];
  assign t[96] = t[148] ^ x[29];
  assign t[97] = t[149] ^ x[30];
  assign t[98] = t[150] ^ x[36];
  assign t[99] = t[151] ^ x[33];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind272(x, y);
 input [71:0] x;
 output y;

 wire [208:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[156] ^ x[5];
  assign t[101] = t[157] ^ x[11];
  assign t[102] = t[158] ^ x[8];
  assign t[103] = t[159] ^ x[9];
  assign t[104] = t[160] ^ x[10];
  assign t[105] = t[161] ^ x[16];
  assign t[106] = t[162] ^ x[13];
  assign t[107] = t[163] ^ x[14];
  assign t[108] = t[164] ^ x[15];
  assign t[109] = t[165] ^ x[21];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[166] ^ x[18];
  assign t[111] = t[167] ^ x[19];
  assign t[112] = t[168] ^ x[20];
  assign t[113] = t[169] ^ x[26];
  assign t[114] = t[170] ^ x[23];
  assign t[115] = t[171] ^ x[24];
  assign t[116] = t[172] ^ x[25];
  assign t[117] = t[173] ^ x[31];
  assign t[118] = t[174] ^ x[28];
  assign t[119] = t[175] ^ x[29];
  assign t[11] = t[19] & t[20];
  assign t[120] = t[176] ^ x[30];
  assign t[121] = t[177] ^ x[36];
  assign t[122] = t[178] ^ x[33];
  assign t[123] = t[179] ^ x[34];
  assign t[124] = t[180] ^ x[35];
  assign t[125] = t[181] ^ x[41];
  assign t[126] = t[182] ^ x[38];
  assign t[127] = t[183] ^ x[39];
  assign t[128] = t[184] ^ x[40];
  assign t[129] = t[185] ^ x[46];
  assign t[12] = ~t[21];
  assign t[130] = t[186] ^ x[43];
  assign t[131] = t[187] ^ x[44];
  assign t[132] = t[188] ^ x[45];
  assign t[133] = t[189] ^ x[51];
  assign t[134] = t[190] ^ x[48];
  assign t[135] = t[191] ^ x[49];
  assign t[136] = t[192] ^ x[50];
  assign t[137] = t[193] ^ x[56];
  assign t[138] = t[194] ^ x[53];
  assign t[139] = t[195] ^ x[54];
  assign t[13] = t[57] & t[22];
  assign t[140] = t[196] ^ x[55];
  assign t[141] = t[197] ^ x[61];
  assign t[142] = t[198] ^ x[58];
  assign t[143] = t[199] ^ x[59];
  assign t[144] = t[200] ^ x[60];
  assign t[145] = t[201] ^ x[66];
  assign t[146] = t[202] ^ x[63];
  assign t[147] = t[203] ^ x[64];
  assign t[148] = t[204] ^ x[65];
  assign t[149] = t[205] ^ x[71];
  assign t[14] = t[23] & t[24];
  assign t[150] = t[206] ^ x[68];
  assign t[151] = t[207] ^ x[69];
  assign t[152] = t[208] ^ x[70];
  assign t[153] = (x[2]);
  assign t[154] = (x[2]);
  assign t[155] = (x[2]);
  assign t[156] = (x[2]);
  assign t[157] = (x[7]);
  assign t[158] = (x[7]);
  assign t[159] = (x[7]);
  assign t[15] = t[25] ^ t[23];
  assign t[160] = (x[7]);
  assign t[161] = (x[12]);
  assign t[162] = (x[12]);
  assign t[163] = (x[12]);
  assign t[164] = (x[12]);
  assign t[165] = (x[17]);
  assign t[166] = (x[17]);
  assign t[167] = (x[17]);
  assign t[168] = (x[17]);
  assign t[169] = (x[22]);
  assign t[16] = t[26] ^ t[14];
  assign t[170] = (x[22]);
  assign t[171] = (x[22]);
  assign t[172] = (x[22]);
  assign t[173] = (x[27]);
  assign t[174] = (x[27]);
  assign t[175] = (x[27]);
  assign t[176] = (x[27]);
  assign t[177] = (x[32]);
  assign t[178] = (x[32]);
  assign t[179] = (x[32]);
  assign t[17] = t[58] & t[27];
  assign t[180] = (x[32]);
  assign t[181] = (x[37]);
  assign t[182] = (x[37]);
  assign t[183] = (x[37]);
  assign t[184] = (x[37]);
  assign t[185] = (x[42]);
  assign t[186] = (x[42]);
  assign t[187] = (x[42]);
  assign t[188] = (x[42]);
  assign t[189] = (x[47]);
  assign t[18] = t[28] & t[29];
  assign t[190] = (x[47]);
  assign t[191] = (x[47]);
  assign t[192] = (x[47]);
  assign t[193] = (x[52]);
  assign t[194] = (x[52]);
  assign t[195] = (x[52]);
  assign t[196] = (x[52]);
  assign t[197] = (x[57]);
  assign t[198] = (x[57]);
  assign t[199] = (x[57]);
  assign t[19] = t[30] ^ t[28];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[57]);
  assign t[201] = (x[62]);
  assign t[202] = (x[62]);
  assign t[203] = (x[62]);
  assign t[204] = (x[62]);
  assign t[205] = (x[67]);
  assign t[206] = (x[67]);
  assign t[207] = (x[67]);
  assign t[208] = (x[67]);
  assign t[20] = t[31] ^ t[18];
  assign t[21] = t[32] ^ t[33];
  assign t[22] = t[34] ^ t[35];
  assign t[23] = ~(t[59]);
  assign t[24] = ~(t[57] ^ t[23]);
  assign t[25] = t[60] ^ t[59];
  assign t[26] = ~(t[36] ^ t[15]);
  assign t[27] = t[37] ^ t[38];
  assign t[28] = ~(t[61]);
  assign t[29] = ~(t[58] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[55]);
  assign t[30] = t[62] ^ t[61];
  assign t[31] = ~(t[39] ^ t[19]);
  assign t[32] = t[40] ^ t[41];
  assign t[33] = t[42] & t[43];
  assign t[34] = t[57] ^ t[25];
  assign t[35] = t[23] & t[36];
  assign t[36] = t[57] ^ t[44];
  assign t[37] = t[58] ^ t[30];
  assign t[38] = t[28] & t[39];
  assign t[39] = t[58] ^ t[45];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[63] & t[46];
  assign t[41] = t[47] & t[48];
  assign t[42] = t[49] ^ t[47];
  assign t[43] = t[50] ^ t[41];
  assign t[44] = t[59] ^ t[64];
  assign t[45] = t[61] ^ t[65];
  assign t[46] = t[51] ^ t[52];
  assign t[47] = ~(t[66]);
  assign t[48] = ~(t[63] ^ t[47]);
  assign t[49] = t[67] ^ t[66];
  assign t[4] = ~t[7];
  assign t[50] = ~(t[53] ^ t[42]);
  assign t[51] = t[63] ^ t[49];
  assign t[52] = t[47] & t[53];
  assign t[53] = t[63] ^ t[54];
  assign t[54] = t[66] ^ t[68];
  assign t[55] = (t[69]);
  assign t[56] = (t[70]);
  assign t[57] = (t[71]);
  assign t[58] = (t[72]);
  assign t[59] = (t[73]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[74]);
  assign t[61] = (t[75]);
  assign t[62] = (t[76]);
  assign t[63] = (t[77]);
  assign t[64] = (t[78]);
  assign t[65] = (t[79]);
  assign t[66] = (t[80]);
  assign t[67] = (t[81]);
  assign t[68] = (t[82]);
  assign t[69] = t[83] ^ x[6];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[84] ^ x[11];
  assign t[71] = t[85] ^ x[16];
  assign t[72] = t[86] ^ x[21];
  assign t[73] = t[87] ^ x[26];
  assign t[74] = t[88] ^ x[31];
  assign t[75] = t[89] ^ x[36];
  assign t[76] = t[90] ^ x[41];
  assign t[77] = t[91] ^ x[46];
  assign t[78] = t[92] ^ x[51];
  assign t[79] = t[93] ^ x[56];
  assign t[7] = ~(t[12] ^ t[56]);
  assign t[80] = t[94] ^ x[61];
  assign t[81] = t[95] ^ x[66];
  assign t[82] = t[96] ^ x[71];
  assign t[83] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[84] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[85] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[86] = (~t[109] & t[110] & t[111] & t[112]) | (t[109] & ~t[111] & ~t[112]) | (t[109] & ~t[110] & ~t[112]) | (t[109] & ~t[110] & ~t[111]);
  assign t[87] = (~t[113] & t[114] & t[115] & t[116]) | (t[113] & ~t[115] & ~t[116]) | (t[113] & ~t[114] & ~t[116]) | (t[113] & ~t[114] & ~t[115]);
  assign t[88] = (~t[117] & t[118] & t[119] & t[120]) | (t[117] & ~t[119] & ~t[120]) | (t[117] & ~t[118] & ~t[120]) | (t[117] & ~t[118] & ~t[119]);
  assign t[89] = (~t[121] & t[122] & t[123] & t[124]) | (t[121] & ~t[123] & ~t[124]) | (t[121] & ~t[122] & ~t[124]) | (t[121] & ~t[122] & ~t[123]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (~t[125] & t[126] & t[127] & t[128]) | (t[125] & ~t[127] & ~t[128]) | (t[125] & ~t[126] & ~t[128]) | (t[125] & ~t[126] & ~t[127]);
  assign t[91] = (~t[129] & t[130] & t[131] & t[132]) | (t[129] & ~t[131] & ~t[132]) | (t[129] & ~t[130] & ~t[132]) | (t[129] & ~t[130] & ~t[131]);
  assign t[92] = (~t[133] & t[134] & t[135] & t[136]) | (t[133] & ~t[135] & ~t[136]) | (t[133] & ~t[134] & ~t[136]) | (t[133] & ~t[134] & ~t[135]);
  assign t[93] = (~t[137] & t[138] & t[139] & t[140]) | (t[137] & ~t[139] & ~t[140]) | (t[137] & ~t[138] & ~t[140]) | (t[137] & ~t[138] & ~t[139]);
  assign t[94] = (~t[141] & t[142] & t[143] & t[144]) | (t[141] & ~t[143] & ~t[144]) | (t[141] & ~t[142] & ~t[144]) | (t[141] & ~t[142] & ~t[143]);
  assign t[95] = (~t[145] & t[146] & t[147] & t[148]) | (t[145] & ~t[147] & ~t[148]) | (t[145] & ~t[146] & ~t[148]) | (t[145] & ~t[146] & ~t[147]);
  assign t[96] = (~t[149] & t[150] & t[151] & t[152]) | (t[149] & ~t[151] & ~t[152]) | (t[149] & ~t[150] & ~t[152]) | (t[149] & ~t[150] & ~t[151]);
  assign t[97] = t[153] ^ x[6];
  assign t[98] = t[154] ^ x[3];
  assign t[99] = t[155] ^ x[4];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind273(x, y);
 input [71:0] x;
 output y;

 wire [208:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[156] ^ x[5];
  assign t[101] = t[157] ^ x[11];
  assign t[102] = t[158] ^ x[8];
  assign t[103] = t[159] ^ x[9];
  assign t[104] = t[160] ^ x[10];
  assign t[105] = t[161] ^ x[16];
  assign t[106] = t[162] ^ x[13];
  assign t[107] = t[163] ^ x[14];
  assign t[108] = t[164] ^ x[15];
  assign t[109] = t[165] ^ x[21];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[166] ^ x[18];
  assign t[111] = t[167] ^ x[19];
  assign t[112] = t[168] ^ x[20];
  assign t[113] = t[169] ^ x[26];
  assign t[114] = t[170] ^ x[23];
  assign t[115] = t[171] ^ x[24];
  assign t[116] = t[172] ^ x[25];
  assign t[117] = t[173] ^ x[31];
  assign t[118] = t[174] ^ x[28];
  assign t[119] = t[175] ^ x[29];
  assign t[11] = t[19] & t[20];
  assign t[120] = t[176] ^ x[30];
  assign t[121] = t[177] ^ x[36];
  assign t[122] = t[178] ^ x[33];
  assign t[123] = t[179] ^ x[34];
  assign t[124] = t[180] ^ x[35];
  assign t[125] = t[181] ^ x[41];
  assign t[126] = t[182] ^ x[38];
  assign t[127] = t[183] ^ x[39];
  assign t[128] = t[184] ^ x[40];
  assign t[129] = t[185] ^ x[46];
  assign t[12] = ~t[21];
  assign t[130] = t[186] ^ x[43];
  assign t[131] = t[187] ^ x[44];
  assign t[132] = t[188] ^ x[45];
  assign t[133] = t[189] ^ x[51];
  assign t[134] = t[190] ^ x[48];
  assign t[135] = t[191] ^ x[49];
  assign t[136] = t[192] ^ x[50];
  assign t[137] = t[193] ^ x[56];
  assign t[138] = t[194] ^ x[53];
  assign t[139] = t[195] ^ x[54];
  assign t[13] = t[57] & t[22];
  assign t[140] = t[196] ^ x[55];
  assign t[141] = t[197] ^ x[61];
  assign t[142] = t[198] ^ x[58];
  assign t[143] = t[199] ^ x[59];
  assign t[144] = t[200] ^ x[60];
  assign t[145] = t[201] ^ x[66];
  assign t[146] = t[202] ^ x[63];
  assign t[147] = t[203] ^ x[64];
  assign t[148] = t[204] ^ x[65];
  assign t[149] = t[205] ^ x[71];
  assign t[14] = t[23] & t[24];
  assign t[150] = t[206] ^ x[68];
  assign t[151] = t[207] ^ x[69];
  assign t[152] = t[208] ^ x[70];
  assign t[153] = (x[2]);
  assign t[154] = (x[2]);
  assign t[155] = (x[2]);
  assign t[156] = (x[2]);
  assign t[157] = (x[7]);
  assign t[158] = (x[7]);
  assign t[159] = (x[7]);
  assign t[15] = t[25] ^ t[23];
  assign t[160] = (x[7]);
  assign t[161] = (x[12]);
  assign t[162] = (x[12]);
  assign t[163] = (x[12]);
  assign t[164] = (x[12]);
  assign t[165] = (x[17]);
  assign t[166] = (x[17]);
  assign t[167] = (x[17]);
  assign t[168] = (x[17]);
  assign t[169] = (x[22]);
  assign t[16] = t[26] ^ t[14];
  assign t[170] = (x[22]);
  assign t[171] = (x[22]);
  assign t[172] = (x[22]);
  assign t[173] = (x[27]);
  assign t[174] = (x[27]);
  assign t[175] = (x[27]);
  assign t[176] = (x[27]);
  assign t[177] = (x[32]);
  assign t[178] = (x[32]);
  assign t[179] = (x[32]);
  assign t[17] = t[58] & t[27];
  assign t[180] = (x[32]);
  assign t[181] = (x[37]);
  assign t[182] = (x[37]);
  assign t[183] = (x[37]);
  assign t[184] = (x[37]);
  assign t[185] = (x[42]);
  assign t[186] = (x[42]);
  assign t[187] = (x[42]);
  assign t[188] = (x[42]);
  assign t[189] = (x[47]);
  assign t[18] = t[28] & t[29];
  assign t[190] = (x[47]);
  assign t[191] = (x[47]);
  assign t[192] = (x[47]);
  assign t[193] = (x[52]);
  assign t[194] = (x[52]);
  assign t[195] = (x[52]);
  assign t[196] = (x[52]);
  assign t[197] = (x[57]);
  assign t[198] = (x[57]);
  assign t[199] = (x[57]);
  assign t[19] = t[30] ^ t[28];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[57]);
  assign t[201] = (x[62]);
  assign t[202] = (x[62]);
  assign t[203] = (x[62]);
  assign t[204] = (x[62]);
  assign t[205] = (x[67]);
  assign t[206] = (x[67]);
  assign t[207] = (x[67]);
  assign t[208] = (x[67]);
  assign t[20] = t[31] ^ t[18];
  assign t[21] = t[32] ^ t[33];
  assign t[22] = t[34] ^ t[35];
  assign t[23] = ~(t[59]);
  assign t[24] = ~(t[57] ^ t[23]);
  assign t[25] = t[60] ^ t[59];
  assign t[26] = ~(t[36] ^ t[15]);
  assign t[27] = t[37] ^ t[38];
  assign t[28] = ~(t[61]);
  assign t[29] = ~(t[58] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[55]);
  assign t[30] = t[62] ^ t[61];
  assign t[31] = ~(t[39] ^ t[19]);
  assign t[32] = t[40] ^ t[41];
  assign t[33] = t[42] & t[43];
  assign t[34] = t[57] ^ t[25];
  assign t[35] = t[23] & t[36];
  assign t[36] = t[57] ^ t[44];
  assign t[37] = t[58] ^ t[30];
  assign t[38] = t[28] & t[39];
  assign t[39] = t[58] ^ t[45];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[63] & t[46];
  assign t[41] = t[47] & t[48];
  assign t[42] = t[49] ^ t[47];
  assign t[43] = t[50] ^ t[41];
  assign t[44] = t[59] ^ t[64];
  assign t[45] = t[61] ^ t[65];
  assign t[46] = t[51] ^ t[52];
  assign t[47] = ~(t[66]);
  assign t[48] = ~(t[63] ^ t[47]);
  assign t[49] = t[67] ^ t[66];
  assign t[4] = ~t[7];
  assign t[50] = ~(t[53] ^ t[42]);
  assign t[51] = t[63] ^ t[49];
  assign t[52] = t[47] & t[53];
  assign t[53] = t[63] ^ t[54];
  assign t[54] = t[66] ^ t[68];
  assign t[55] = (t[69]);
  assign t[56] = (t[70]);
  assign t[57] = (t[71]);
  assign t[58] = (t[72]);
  assign t[59] = (t[73]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[74]);
  assign t[61] = (t[75]);
  assign t[62] = (t[76]);
  assign t[63] = (t[77]);
  assign t[64] = (t[78]);
  assign t[65] = (t[79]);
  assign t[66] = (t[80]);
  assign t[67] = (t[81]);
  assign t[68] = (t[82]);
  assign t[69] = t[83] ^ x[6];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[84] ^ x[11];
  assign t[71] = t[85] ^ x[16];
  assign t[72] = t[86] ^ x[21];
  assign t[73] = t[87] ^ x[26];
  assign t[74] = t[88] ^ x[31];
  assign t[75] = t[89] ^ x[36];
  assign t[76] = t[90] ^ x[41];
  assign t[77] = t[91] ^ x[46];
  assign t[78] = t[92] ^ x[51];
  assign t[79] = t[93] ^ x[56];
  assign t[7] = ~(t[12] ^ t[56]);
  assign t[80] = t[94] ^ x[61];
  assign t[81] = t[95] ^ x[66];
  assign t[82] = t[96] ^ x[71];
  assign t[83] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[84] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[85] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[86] = (~t[109] & t[110] & t[111] & t[112]) | (t[109] & ~t[111] & ~t[112]) | (t[109] & ~t[110] & ~t[112]) | (t[109] & ~t[110] & ~t[111]);
  assign t[87] = (~t[113] & t[114] & t[115] & t[116]) | (t[113] & ~t[115] & ~t[116]) | (t[113] & ~t[114] & ~t[116]) | (t[113] & ~t[114] & ~t[115]);
  assign t[88] = (~t[117] & t[118] & t[119] & t[120]) | (t[117] & ~t[119] & ~t[120]) | (t[117] & ~t[118] & ~t[120]) | (t[117] & ~t[118] & ~t[119]);
  assign t[89] = (~t[121] & t[122] & t[123] & t[124]) | (t[121] & ~t[123] & ~t[124]) | (t[121] & ~t[122] & ~t[124]) | (t[121] & ~t[122] & ~t[123]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (~t[125] & t[126] & t[127] & t[128]) | (t[125] & ~t[127] & ~t[128]) | (t[125] & ~t[126] & ~t[128]) | (t[125] & ~t[126] & ~t[127]);
  assign t[91] = (~t[129] & t[130] & t[131] & t[132]) | (t[129] & ~t[131] & ~t[132]) | (t[129] & ~t[130] & ~t[132]) | (t[129] & ~t[130] & ~t[131]);
  assign t[92] = (~t[133] & t[134] & t[135] & t[136]) | (t[133] & ~t[135] & ~t[136]) | (t[133] & ~t[134] & ~t[136]) | (t[133] & ~t[134] & ~t[135]);
  assign t[93] = (~t[137] & t[138] & t[139] & t[140]) | (t[137] & ~t[139] & ~t[140]) | (t[137] & ~t[138] & ~t[140]) | (t[137] & ~t[138] & ~t[139]);
  assign t[94] = (~t[141] & t[142] & t[143] & t[144]) | (t[141] & ~t[143] & ~t[144]) | (t[141] & ~t[142] & ~t[144]) | (t[141] & ~t[142] & ~t[143]);
  assign t[95] = (~t[145] & t[146] & t[147] & t[148]) | (t[145] & ~t[147] & ~t[148]) | (t[145] & ~t[146] & ~t[148]) | (t[145] & ~t[146] & ~t[147]);
  assign t[96] = (~t[149] & t[150] & t[151] & t[152]) | (t[149] & ~t[151] & ~t[152]) | (t[149] & ~t[150] & ~t[152]) | (t[149] & ~t[150] & ~t[151]);
  assign t[97] = t[153] ^ x[6];
  assign t[98] = t[154] ^ x[3];
  assign t[99] = t[155] ^ x[4];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind274(x, y);
 input [71:0] x;
 output y;

 wire [208:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[156] ^ x[5];
  assign t[101] = t[157] ^ x[11];
  assign t[102] = t[158] ^ x[8];
  assign t[103] = t[159] ^ x[9];
  assign t[104] = t[160] ^ x[10];
  assign t[105] = t[161] ^ x[16];
  assign t[106] = t[162] ^ x[13];
  assign t[107] = t[163] ^ x[14];
  assign t[108] = t[164] ^ x[15];
  assign t[109] = t[165] ^ x[21];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[166] ^ x[18];
  assign t[111] = t[167] ^ x[19];
  assign t[112] = t[168] ^ x[20];
  assign t[113] = t[169] ^ x[26];
  assign t[114] = t[170] ^ x[23];
  assign t[115] = t[171] ^ x[24];
  assign t[116] = t[172] ^ x[25];
  assign t[117] = t[173] ^ x[31];
  assign t[118] = t[174] ^ x[28];
  assign t[119] = t[175] ^ x[29];
  assign t[11] = t[19] & t[20];
  assign t[120] = t[176] ^ x[30];
  assign t[121] = t[177] ^ x[36];
  assign t[122] = t[178] ^ x[33];
  assign t[123] = t[179] ^ x[34];
  assign t[124] = t[180] ^ x[35];
  assign t[125] = t[181] ^ x[41];
  assign t[126] = t[182] ^ x[38];
  assign t[127] = t[183] ^ x[39];
  assign t[128] = t[184] ^ x[40];
  assign t[129] = t[185] ^ x[46];
  assign t[12] = ~t[21];
  assign t[130] = t[186] ^ x[43];
  assign t[131] = t[187] ^ x[44];
  assign t[132] = t[188] ^ x[45];
  assign t[133] = t[189] ^ x[51];
  assign t[134] = t[190] ^ x[48];
  assign t[135] = t[191] ^ x[49];
  assign t[136] = t[192] ^ x[50];
  assign t[137] = t[193] ^ x[56];
  assign t[138] = t[194] ^ x[53];
  assign t[139] = t[195] ^ x[54];
  assign t[13] = t[57] & t[22];
  assign t[140] = t[196] ^ x[55];
  assign t[141] = t[197] ^ x[61];
  assign t[142] = t[198] ^ x[58];
  assign t[143] = t[199] ^ x[59];
  assign t[144] = t[200] ^ x[60];
  assign t[145] = t[201] ^ x[66];
  assign t[146] = t[202] ^ x[63];
  assign t[147] = t[203] ^ x[64];
  assign t[148] = t[204] ^ x[65];
  assign t[149] = t[205] ^ x[71];
  assign t[14] = t[23] & t[24];
  assign t[150] = t[206] ^ x[68];
  assign t[151] = t[207] ^ x[69];
  assign t[152] = t[208] ^ x[70];
  assign t[153] = (x[2]);
  assign t[154] = (x[2]);
  assign t[155] = (x[2]);
  assign t[156] = (x[2]);
  assign t[157] = (x[7]);
  assign t[158] = (x[7]);
  assign t[159] = (x[7]);
  assign t[15] = t[25] ^ t[23];
  assign t[160] = (x[7]);
  assign t[161] = (x[12]);
  assign t[162] = (x[12]);
  assign t[163] = (x[12]);
  assign t[164] = (x[12]);
  assign t[165] = (x[17]);
  assign t[166] = (x[17]);
  assign t[167] = (x[17]);
  assign t[168] = (x[17]);
  assign t[169] = (x[22]);
  assign t[16] = t[26] ^ t[14];
  assign t[170] = (x[22]);
  assign t[171] = (x[22]);
  assign t[172] = (x[22]);
  assign t[173] = (x[27]);
  assign t[174] = (x[27]);
  assign t[175] = (x[27]);
  assign t[176] = (x[27]);
  assign t[177] = (x[32]);
  assign t[178] = (x[32]);
  assign t[179] = (x[32]);
  assign t[17] = t[58] & t[27];
  assign t[180] = (x[32]);
  assign t[181] = (x[37]);
  assign t[182] = (x[37]);
  assign t[183] = (x[37]);
  assign t[184] = (x[37]);
  assign t[185] = (x[42]);
  assign t[186] = (x[42]);
  assign t[187] = (x[42]);
  assign t[188] = (x[42]);
  assign t[189] = (x[47]);
  assign t[18] = t[28] & t[29];
  assign t[190] = (x[47]);
  assign t[191] = (x[47]);
  assign t[192] = (x[47]);
  assign t[193] = (x[52]);
  assign t[194] = (x[52]);
  assign t[195] = (x[52]);
  assign t[196] = (x[52]);
  assign t[197] = (x[57]);
  assign t[198] = (x[57]);
  assign t[199] = (x[57]);
  assign t[19] = t[30] ^ t[28];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[57]);
  assign t[201] = (x[62]);
  assign t[202] = (x[62]);
  assign t[203] = (x[62]);
  assign t[204] = (x[62]);
  assign t[205] = (x[67]);
  assign t[206] = (x[67]);
  assign t[207] = (x[67]);
  assign t[208] = (x[67]);
  assign t[20] = t[31] ^ t[18];
  assign t[21] = t[32] ^ t[33];
  assign t[22] = t[34] ^ t[35];
  assign t[23] = ~(t[59]);
  assign t[24] = ~(t[57] ^ t[23]);
  assign t[25] = t[60] ^ t[59];
  assign t[26] = ~(t[36] ^ t[15]);
  assign t[27] = t[37] ^ t[38];
  assign t[28] = ~(t[61]);
  assign t[29] = ~(t[58] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[55]);
  assign t[30] = t[62] ^ t[61];
  assign t[31] = ~(t[39] ^ t[19]);
  assign t[32] = t[40] ^ t[41];
  assign t[33] = t[42] & t[43];
  assign t[34] = t[57] ^ t[25];
  assign t[35] = t[23] & t[36];
  assign t[36] = t[57] ^ t[44];
  assign t[37] = t[58] ^ t[30];
  assign t[38] = t[28] & t[39];
  assign t[39] = t[58] ^ t[45];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[63] & t[46];
  assign t[41] = t[47] & t[48];
  assign t[42] = t[49] ^ t[47];
  assign t[43] = t[50] ^ t[41];
  assign t[44] = t[59] ^ t[64];
  assign t[45] = t[61] ^ t[65];
  assign t[46] = t[51] ^ t[52];
  assign t[47] = ~(t[66]);
  assign t[48] = ~(t[63] ^ t[47]);
  assign t[49] = t[67] ^ t[66];
  assign t[4] = ~t[7];
  assign t[50] = ~(t[53] ^ t[42]);
  assign t[51] = t[63] ^ t[49];
  assign t[52] = t[47] & t[53];
  assign t[53] = t[63] ^ t[54];
  assign t[54] = t[66] ^ t[68];
  assign t[55] = (t[69]);
  assign t[56] = (t[70]);
  assign t[57] = (t[71]);
  assign t[58] = (t[72]);
  assign t[59] = (t[73]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[74]);
  assign t[61] = (t[75]);
  assign t[62] = (t[76]);
  assign t[63] = (t[77]);
  assign t[64] = (t[78]);
  assign t[65] = (t[79]);
  assign t[66] = (t[80]);
  assign t[67] = (t[81]);
  assign t[68] = (t[82]);
  assign t[69] = t[83] ^ x[6];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[84] ^ x[11];
  assign t[71] = t[85] ^ x[16];
  assign t[72] = t[86] ^ x[21];
  assign t[73] = t[87] ^ x[26];
  assign t[74] = t[88] ^ x[31];
  assign t[75] = t[89] ^ x[36];
  assign t[76] = t[90] ^ x[41];
  assign t[77] = t[91] ^ x[46];
  assign t[78] = t[92] ^ x[51];
  assign t[79] = t[93] ^ x[56];
  assign t[7] = ~(t[12] ^ t[56]);
  assign t[80] = t[94] ^ x[61];
  assign t[81] = t[95] ^ x[66];
  assign t[82] = t[96] ^ x[71];
  assign t[83] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[84] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[85] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[86] = (~t[109] & t[110] & t[111] & t[112]) | (t[109] & ~t[111] & ~t[112]) | (t[109] & ~t[110] & ~t[112]) | (t[109] & ~t[110] & ~t[111]);
  assign t[87] = (~t[113] & t[114] & t[115] & t[116]) | (t[113] & ~t[115] & ~t[116]) | (t[113] & ~t[114] & ~t[116]) | (t[113] & ~t[114] & ~t[115]);
  assign t[88] = (~t[117] & t[118] & t[119] & t[120]) | (t[117] & ~t[119] & ~t[120]) | (t[117] & ~t[118] & ~t[120]) | (t[117] & ~t[118] & ~t[119]);
  assign t[89] = (~t[121] & t[122] & t[123] & t[124]) | (t[121] & ~t[123] & ~t[124]) | (t[121] & ~t[122] & ~t[124]) | (t[121] & ~t[122] & ~t[123]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (~t[125] & t[126] & t[127] & t[128]) | (t[125] & ~t[127] & ~t[128]) | (t[125] & ~t[126] & ~t[128]) | (t[125] & ~t[126] & ~t[127]);
  assign t[91] = (~t[129] & t[130] & t[131] & t[132]) | (t[129] & ~t[131] & ~t[132]) | (t[129] & ~t[130] & ~t[132]) | (t[129] & ~t[130] & ~t[131]);
  assign t[92] = (~t[133] & t[134] & t[135] & t[136]) | (t[133] & ~t[135] & ~t[136]) | (t[133] & ~t[134] & ~t[136]) | (t[133] & ~t[134] & ~t[135]);
  assign t[93] = (~t[137] & t[138] & t[139] & t[140]) | (t[137] & ~t[139] & ~t[140]) | (t[137] & ~t[138] & ~t[140]) | (t[137] & ~t[138] & ~t[139]);
  assign t[94] = (~t[141] & t[142] & t[143] & t[144]) | (t[141] & ~t[143] & ~t[144]) | (t[141] & ~t[142] & ~t[144]) | (t[141] & ~t[142] & ~t[143]);
  assign t[95] = (~t[145] & t[146] & t[147] & t[148]) | (t[145] & ~t[147] & ~t[148]) | (t[145] & ~t[146] & ~t[148]) | (t[145] & ~t[146] & ~t[147]);
  assign t[96] = (~t[149] & t[150] & t[151] & t[152]) | (t[149] & ~t[151] & ~t[152]) | (t[149] & ~t[150] & ~t[152]) | (t[149] & ~t[150] & ~t[151]);
  assign t[97] = t[153] ^ x[6];
  assign t[98] = t[154] ^ x[3];
  assign t[99] = t[155] ^ x[4];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind275(x, y);
 input [71:0] x;
 output y;

 wire [208:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[156] ^ x[5];
  assign t[101] = t[157] ^ x[11];
  assign t[102] = t[158] ^ x[8];
  assign t[103] = t[159] ^ x[9];
  assign t[104] = t[160] ^ x[10];
  assign t[105] = t[161] ^ x[16];
  assign t[106] = t[162] ^ x[13];
  assign t[107] = t[163] ^ x[14];
  assign t[108] = t[164] ^ x[15];
  assign t[109] = t[165] ^ x[21];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[166] ^ x[18];
  assign t[111] = t[167] ^ x[19];
  assign t[112] = t[168] ^ x[20];
  assign t[113] = t[169] ^ x[26];
  assign t[114] = t[170] ^ x[23];
  assign t[115] = t[171] ^ x[24];
  assign t[116] = t[172] ^ x[25];
  assign t[117] = t[173] ^ x[31];
  assign t[118] = t[174] ^ x[28];
  assign t[119] = t[175] ^ x[29];
  assign t[11] = t[19] & t[20];
  assign t[120] = t[176] ^ x[30];
  assign t[121] = t[177] ^ x[36];
  assign t[122] = t[178] ^ x[33];
  assign t[123] = t[179] ^ x[34];
  assign t[124] = t[180] ^ x[35];
  assign t[125] = t[181] ^ x[41];
  assign t[126] = t[182] ^ x[38];
  assign t[127] = t[183] ^ x[39];
  assign t[128] = t[184] ^ x[40];
  assign t[129] = t[185] ^ x[46];
  assign t[12] = ~t[21];
  assign t[130] = t[186] ^ x[43];
  assign t[131] = t[187] ^ x[44];
  assign t[132] = t[188] ^ x[45];
  assign t[133] = t[189] ^ x[51];
  assign t[134] = t[190] ^ x[48];
  assign t[135] = t[191] ^ x[49];
  assign t[136] = t[192] ^ x[50];
  assign t[137] = t[193] ^ x[56];
  assign t[138] = t[194] ^ x[53];
  assign t[139] = t[195] ^ x[54];
  assign t[13] = t[57] & t[22];
  assign t[140] = t[196] ^ x[55];
  assign t[141] = t[197] ^ x[61];
  assign t[142] = t[198] ^ x[58];
  assign t[143] = t[199] ^ x[59];
  assign t[144] = t[200] ^ x[60];
  assign t[145] = t[201] ^ x[66];
  assign t[146] = t[202] ^ x[63];
  assign t[147] = t[203] ^ x[64];
  assign t[148] = t[204] ^ x[65];
  assign t[149] = t[205] ^ x[71];
  assign t[14] = t[23] & t[24];
  assign t[150] = t[206] ^ x[68];
  assign t[151] = t[207] ^ x[69];
  assign t[152] = t[208] ^ x[70];
  assign t[153] = (x[2]);
  assign t[154] = (x[2]);
  assign t[155] = (x[2]);
  assign t[156] = (x[2]);
  assign t[157] = (x[7]);
  assign t[158] = (x[7]);
  assign t[159] = (x[7]);
  assign t[15] = t[25] ^ t[23];
  assign t[160] = (x[7]);
  assign t[161] = (x[12]);
  assign t[162] = (x[12]);
  assign t[163] = (x[12]);
  assign t[164] = (x[12]);
  assign t[165] = (x[17]);
  assign t[166] = (x[17]);
  assign t[167] = (x[17]);
  assign t[168] = (x[17]);
  assign t[169] = (x[22]);
  assign t[16] = t[26] ^ t[14];
  assign t[170] = (x[22]);
  assign t[171] = (x[22]);
  assign t[172] = (x[22]);
  assign t[173] = (x[27]);
  assign t[174] = (x[27]);
  assign t[175] = (x[27]);
  assign t[176] = (x[27]);
  assign t[177] = (x[32]);
  assign t[178] = (x[32]);
  assign t[179] = (x[32]);
  assign t[17] = t[58] & t[27];
  assign t[180] = (x[32]);
  assign t[181] = (x[37]);
  assign t[182] = (x[37]);
  assign t[183] = (x[37]);
  assign t[184] = (x[37]);
  assign t[185] = (x[42]);
  assign t[186] = (x[42]);
  assign t[187] = (x[42]);
  assign t[188] = (x[42]);
  assign t[189] = (x[47]);
  assign t[18] = t[28] & t[29];
  assign t[190] = (x[47]);
  assign t[191] = (x[47]);
  assign t[192] = (x[47]);
  assign t[193] = (x[52]);
  assign t[194] = (x[52]);
  assign t[195] = (x[52]);
  assign t[196] = (x[52]);
  assign t[197] = (x[57]);
  assign t[198] = (x[57]);
  assign t[199] = (x[57]);
  assign t[19] = t[30] ^ t[28];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[57]);
  assign t[201] = (x[62]);
  assign t[202] = (x[62]);
  assign t[203] = (x[62]);
  assign t[204] = (x[62]);
  assign t[205] = (x[67]);
  assign t[206] = (x[67]);
  assign t[207] = (x[67]);
  assign t[208] = (x[67]);
  assign t[20] = t[31] ^ t[18];
  assign t[21] = t[32] ^ t[33];
  assign t[22] = t[34] ^ t[35];
  assign t[23] = ~(t[59]);
  assign t[24] = ~(t[57] ^ t[23]);
  assign t[25] = t[60] ^ t[59];
  assign t[26] = ~(t[36] ^ t[15]);
  assign t[27] = t[37] ^ t[38];
  assign t[28] = ~(t[61]);
  assign t[29] = ~(t[58] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[55]);
  assign t[30] = t[62] ^ t[61];
  assign t[31] = ~(t[39] ^ t[19]);
  assign t[32] = t[40] ^ t[41];
  assign t[33] = t[42] & t[43];
  assign t[34] = t[57] ^ t[25];
  assign t[35] = t[23] & t[36];
  assign t[36] = t[57] ^ t[44];
  assign t[37] = t[58] ^ t[30];
  assign t[38] = t[28] & t[39];
  assign t[39] = t[58] ^ t[45];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[63] & t[46];
  assign t[41] = t[47] & t[48];
  assign t[42] = t[49] ^ t[47];
  assign t[43] = t[50] ^ t[41];
  assign t[44] = t[59] ^ t[64];
  assign t[45] = t[61] ^ t[65];
  assign t[46] = t[51] ^ t[52];
  assign t[47] = ~(t[66]);
  assign t[48] = ~(t[63] ^ t[47]);
  assign t[49] = t[67] ^ t[66];
  assign t[4] = ~t[7];
  assign t[50] = ~(t[53] ^ t[42]);
  assign t[51] = t[63] ^ t[49];
  assign t[52] = t[47] & t[53];
  assign t[53] = t[63] ^ t[54];
  assign t[54] = t[66] ^ t[68];
  assign t[55] = (t[69]);
  assign t[56] = (t[70]);
  assign t[57] = (t[71]);
  assign t[58] = (t[72]);
  assign t[59] = (t[73]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[74]);
  assign t[61] = (t[75]);
  assign t[62] = (t[76]);
  assign t[63] = (t[77]);
  assign t[64] = (t[78]);
  assign t[65] = (t[79]);
  assign t[66] = (t[80]);
  assign t[67] = (t[81]);
  assign t[68] = (t[82]);
  assign t[69] = t[83] ^ x[6];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[84] ^ x[11];
  assign t[71] = t[85] ^ x[16];
  assign t[72] = t[86] ^ x[21];
  assign t[73] = t[87] ^ x[26];
  assign t[74] = t[88] ^ x[31];
  assign t[75] = t[89] ^ x[36];
  assign t[76] = t[90] ^ x[41];
  assign t[77] = t[91] ^ x[46];
  assign t[78] = t[92] ^ x[51];
  assign t[79] = t[93] ^ x[56];
  assign t[7] = ~(t[12] ^ t[56]);
  assign t[80] = t[94] ^ x[61];
  assign t[81] = t[95] ^ x[66];
  assign t[82] = t[96] ^ x[71];
  assign t[83] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[84] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[85] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[86] = (~t[109] & t[110] & t[111] & t[112]) | (t[109] & ~t[111] & ~t[112]) | (t[109] & ~t[110] & ~t[112]) | (t[109] & ~t[110] & ~t[111]);
  assign t[87] = (~t[113] & t[114] & t[115] & t[116]) | (t[113] & ~t[115] & ~t[116]) | (t[113] & ~t[114] & ~t[116]) | (t[113] & ~t[114] & ~t[115]);
  assign t[88] = (~t[117] & t[118] & t[119] & t[120]) | (t[117] & ~t[119] & ~t[120]) | (t[117] & ~t[118] & ~t[120]) | (t[117] & ~t[118] & ~t[119]);
  assign t[89] = (~t[121] & t[122] & t[123] & t[124]) | (t[121] & ~t[123] & ~t[124]) | (t[121] & ~t[122] & ~t[124]) | (t[121] & ~t[122] & ~t[123]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (~t[125] & t[126] & t[127] & t[128]) | (t[125] & ~t[127] & ~t[128]) | (t[125] & ~t[126] & ~t[128]) | (t[125] & ~t[126] & ~t[127]);
  assign t[91] = (~t[129] & t[130] & t[131] & t[132]) | (t[129] & ~t[131] & ~t[132]) | (t[129] & ~t[130] & ~t[132]) | (t[129] & ~t[130] & ~t[131]);
  assign t[92] = (~t[133] & t[134] & t[135] & t[136]) | (t[133] & ~t[135] & ~t[136]) | (t[133] & ~t[134] & ~t[136]) | (t[133] & ~t[134] & ~t[135]);
  assign t[93] = (~t[137] & t[138] & t[139] & t[140]) | (t[137] & ~t[139] & ~t[140]) | (t[137] & ~t[138] & ~t[140]) | (t[137] & ~t[138] & ~t[139]);
  assign t[94] = (~t[141] & t[142] & t[143] & t[144]) | (t[141] & ~t[143] & ~t[144]) | (t[141] & ~t[142] & ~t[144]) | (t[141] & ~t[142] & ~t[143]);
  assign t[95] = (~t[145] & t[146] & t[147] & t[148]) | (t[145] & ~t[147] & ~t[148]) | (t[145] & ~t[146] & ~t[148]) | (t[145] & ~t[146] & ~t[147]);
  assign t[96] = (~t[149] & t[150] & t[151] & t[152]) | (t[149] & ~t[151] & ~t[152]) | (t[149] & ~t[150] & ~t[152]) | (t[149] & ~t[150] & ~t[151]);
  assign t[97] = t[153] ^ x[6];
  assign t[98] = t[154] ^ x[3];
  assign t[99] = t[155] ^ x[4];
  assign t[9] = t[15] & t[16];
  assign y = (t[0]);
endmodule

module R2ind276(x, y);
 input [71:0] x;
 output y;

 wire [208:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[156] ^ x[5];
  assign t[101] = t[157] ^ x[11];
  assign t[102] = t[158] ^ x[8];
  assign t[103] = t[159] ^ x[9];
  assign t[104] = t[160] ^ x[10];
  assign t[105] = t[161] ^ x[16];
  assign t[106] = t[162] ^ x[13];
  assign t[107] = t[163] ^ x[14];
  assign t[108] = t[164] ^ x[15];
  assign t[109] = t[165] ^ x[21];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[166] ^ x[18];
  assign t[111] = t[167] ^ x[19];
  assign t[112] = t[168] ^ x[20];
  assign t[113] = t[169] ^ x[26];
  assign t[114] = t[170] ^ x[23];
  assign t[115] = t[171] ^ x[24];
  assign t[116] = t[172] ^ x[25];
  assign t[117] = t[173] ^ x[31];
  assign t[118] = t[174] ^ x[28];
  assign t[119] = t[175] ^ x[29];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[176] ^ x[30];
  assign t[121] = t[177] ^ x[36];
  assign t[122] = t[178] ^ x[33];
  assign t[123] = t[179] ^ x[34];
  assign t[124] = t[180] ^ x[35];
  assign t[125] = t[181] ^ x[41];
  assign t[126] = t[182] ^ x[38];
  assign t[127] = t[183] ^ x[39];
  assign t[128] = t[184] ^ x[40];
  assign t[129] = t[185] ^ x[46];
  assign t[12] = ~t[21];
  assign t[130] = t[186] ^ x[43];
  assign t[131] = t[187] ^ x[44];
  assign t[132] = t[188] ^ x[45];
  assign t[133] = t[189] ^ x[51];
  assign t[134] = t[190] ^ x[48];
  assign t[135] = t[191] ^ x[49];
  assign t[136] = t[192] ^ x[50];
  assign t[137] = t[193] ^ x[56];
  assign t[138] = t[194] ^ x[53];
  assign t[139] = t[195] ^ x[54];
  assign t[13] = t[22] ^ t[23];
  assign t[140] = t[196] ^ x[55];
  assign t[141] = t[197] ^ x[61];
  assign t[142] = t[198] ^ x[58];
  assign t[143] = t[199] ^ x[59];
  assign t[144] = t[200] ^ x[60];
  assign t[145] = t[201] ^ x[66];
  assign t[146] = t[202] ^ x[63];
  assign t[147] = t[203] ^ x[64];
  assign t[148] = t[204] ^ x[65];
  assign t[149] = t[205] ^ x[71];
  assign t[14] = t[24] & t[25];
  assign t[150] = t[206] ^ x[68];
  assign t[151] = t[207] ^ x[69];
  assign t[152] = t[208] ^ x[70];
  assign t[153] = (x[2]);
  assign t[154] = (x[2]);
  assign t[155] = (x[2]);
  assign t[156] = (x[2]);
  assign t[157] = (x[7]);
  assign t[158] = (x[7]);
  assign t[159] = (x[7]);
  assign t[15] = t[26] ^ t[14];
  assign t[160] = (x[7]);
  assign t[161] = (x[12]);
  assign t[162] = (x[12]);
  assign t[163] = (x[12]);
  assign t[164] = (x[12]);
  assign t[165] = (x[17]);
  assign t[166] = (x[17]);
  assign t[167] = (x[17]);
  assign t[168] = (x[17]);
  assign t[169] = (x[22]);
  assign t[16] = t[57] ^ t[24];
  assign t[170] = (x[22]);
  assign t[171] = (x[22]);
  assign t[172] = (x[22]);
  assign t[173] = (x[27]);
  assign t[174] = (x[27]);
  assign t[175] = (x[27]);
  assign t[176] = (x[27]);
  assign t[177] = (x[32]);
  assign t[178] = (x[32]);
  assign t[179] = (x[32]);
  assign t[17] = t[27] ^ t[28];
  assign t[180] = (x[32]);
  assign t[181] = (x[37]);
  assign t[182] = (x[37]);
  assign t[183] = (x[37]);
  assign t[184] = (x[37]);
  assign t[185] = (x[42]);
  assign t[186] = (x[42]);
  assign t[187] = (x[42]);
  assign t[188] = (x[42]);
  assign t[189] = (x[47]);
  assign t[18] = t[29] & t[30];
  assign t[190] = (x[47]);
  assign t[191] = (x[47]);
  assign t[192] = (x[47]);
  assign t[193] = (x[52]);
  assign t[194] = (x[52]);
  assign t[195] = (x[52]);
  assign t[196] = (x[52]);
  assign t[197] = (x[57]);
  assign t[198] = (x[57]);
  assign t[199] = (x[57]);
  assign t[19] = t[31] ^ t[18];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[57]);
  assign t[201] = (x[62]);
  assign t[202] = (x[62]);
  assign t[203] = (x[62]);
  assign t[204] = (x[62]);
  assign t[205] = (x[67]);
  assign t[206] = (x[67]);
  assign t[207] = (x[67]);
  assign t[208] = (x[67]);
  assign t[20] = t[58] ^ t[29];
  assign t[21] = ~(t[32] ^ t[33]);
  assign t[22] = t[59] ^ t[60];
  assign t[23] = t[24] & t[34];
  assign t[24] = ~(t[60]);
  assign t[25] = ~(t[57] ^ t[24]);
  assign t[26] = t[57] & t[35];
  assign t[27] = t[61] ^ t[62];
  assign t[28] = t[29] & t[36];
  assign t[29] = ~(t[62]);
  assign t[2] = ~(t[4] ^ t[55]);
  assign t[30] = ~(t[58] ^ t[29]);
  assign t[31] = t[58] & t[37];
  assign t[32] = t[38] ^ t[39];
  assign t[33] = t[40] ^ t[41];
  assign t[34] = t[57] ^ t[42];
  assign t[35] = t[43] ^ t[23];
  assign t[36] = t[58] ^ t[44];
  assign t[37] = t[45] ^ t[28];
  assign t[38] = t[46] ^ t[47];
  assign t[39] = t[48] & t[49];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ t[39];
  assign t[41] = t[63] ^ t[48];
  assign t[42] = t[60] ^ t[64];
  assign t[43] = t[57] ^ t[22];
  assign t[44] = t[62] ^ t[65];
  assign t[45] = t[58] ^ t[27];
  assign t[46] = t[66] ^ t[67];
  assign t[47] = t[48] & t[51];
  assign t[48] = ~(t[67]);
  assign t[49] = ~(t[63] ^ t[48]);
  assign t[4] = ~t[7];
  assign t[50] = t[63] & t[52];
  assign t[51] = t[63] ^ t[53];
  assign t[52] = t[54] ^ t[47];
  assign t[53] = t[67] ^ t[68];
  assign t[54] = t[63] ^ t[46];
  assign t[55] = (t[69]);
  assign t[56] = (t[70]);
  assign t[57] = (t[71]);
  assign t[58] = (t[72]);
  assign t[59] = (t[73]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (t[74]);
  assign t[61] = (t[75]);
  assign t[62] = (t[76]);
  assign t[63] = (t[77]);
  assign t[64] = (t[78]);
  assign t[65] = (t[79]);
  assign t[66] = (t[80]);
  assign t[67] = (t[81]);
  assign t[68] = (t[82]);
  assign t[69] = t[83] ^ x[6];
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = t[84] ^ x[11];
  assign t[71] = t[85] ^ x[16];
  assign t[72] = t[86] ^ x[21];
  assign t[73] = t[87] ^ x[26];
  assign t[74] = t[88] ^ x[31];
  assign t[75] = t[89] ^ x[36];
  assign t[76] = t[90] ^ x[41];
  assign t[77] = t[91] ^ x[46];
  assign t[78] = t[92] ^ x[51];
  assign t[79] = t[93] ^ x[56];
  assign t[7] = ~(t[12] ^ t[56]);
  assign t[80] = t[94] ^ x[61];
  assign t[81] = t[95] ^ x[66];
  assign t[82] = t[96] ^ x[71];
  assign t[83] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[84] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[85] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[86] = (~t[109] & t[110] & t[111] & t[112]) | (t[109] & ~t[111] & ~t[112]) | (t[109] & ~t[110] & ~t[112]) | (t[109] & ~t[110] & ~t[111]);
  assign t[87] = (~t[113] & t[114] & t[115] & t[116]) | (t[113] & ~t[115] & ~t[116]) | (t[113] & ~t[114] & ~t[116]) | (t[113] & ~t[114] & ~t[115]);
  assign t[88] = (~t[117] & t[118] & t[119] & t[120]) | (t[117] & ~t[119] & ~t[120]) | (t[117] & ~t[118] & ~t[120]) | (t[117] & ~t[118] & ~t[119]);
  assign t[89] = (~t[121] & t[122] & t[123] & t[124]) | (t[121] & ~t[123] & ~t[124]) | (t[121] & ~t[122] & ~t[124]) | (t[121] & ~t[122] & ~t[123]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (~t[125] & t[126] & t[127] & t[128]) | (t[125] & ~t[127] & ~t[128]) | (t[125] & ~t[126] & ~t[128]) | (t[125] & ~t[126] & ~t[127]);
  assign t[91] = (~t[129] & t[130] & t[131] & t[132]) | (t[129] & ~t[131] & ~t[132]) | (t[129] & ~t[130] & ~t[132]) | (t[129] & ~t[130] & ~t[131]);
  assign t[92] = (~t[133] & t[134] & t[135] & t[136]) | (t[133] & ~t[135] & ~t[136]) | (t[133] & ~t[134] & ~t[136]) | (t[133] & ~t[134] & ~t[135]);
  assign t[93] = (~t[137] & t[138] & t[139] & t[140]) | (t[137] & ~t[139] & ~t[140]) | (t[137] & ~t[138] & ~t[140]) | (t[137] & ~t[138] & ~t[139]);
  assign t[94] = (~t[141] & t[142] & t[143] & t[144]) | (t[141] & ~t[143] & ~t[144]) | (t[141] & ~t[142] & ~t[144]) | (t[141] & ~t[142] & ~t[143]);
  assign t[95] = (~t[145] & t[146] & t[147] & t[148]) | (t[145] & ~t[147] & ~t[148]) | (t[145] & ~t[146] & ~t[148]) | (t[145] & ~t[146] & ~t[147]);
  assign t[96] = (~t[149] & t[150] & t[151] & t[152]) | (t[149] & ~t[151] & ~t[152]) | (t[149] & ~t[150] & ~t[152]) | (t[149] & ~t[150] & ~t[151]);
  assign t[97] = t[153] ^ x[6];
  assign t[98] = t[154] ^ x[3];
  assign t[99] = t[155] ^ x[4];
  assign t[9] = t[15] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind277(x, y);
 input [71:0] x;
 output y;

 wire [208:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[156] ^ x[5];
  assign t[101] = t[157] ^ x[11];
  assign t[102] = t[158] ^ x[8];
  assign t[103] = t[159] ^ x[9];
  assign t[104] = t[160] ^ x[10];
  assign t[105] = t[161] ^ x[16];
  assign t[106] = t[162] ^ x[13];
  assign t[107] = t[163] ^ x[14];
  assign t[108] = t[164] ^ x[15];
  assign t[109] = t[165] ^ x[21];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[166] ^ x[18];
  assign t[111] = t[167] ^ x[19];
  assign t[112] = t[168] ^ x[20];
  assign t[113] = t[169] ^ x[26];
  assign t[114] = t[170] ^ x[23];
  assign t[115] = t[171] ^ x[24];
  assign t[116] = t[172] ^ x[25];
  assign t[117] = t[173] ^ x[31];
  assign t[118] = t[174] ^ x[28];
  assign t[119] = t[175] ^ x[29];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[176] ^ x[30];
  assign t[121] = t[177] ^ x[36];
  assign t[122] = t[178] ^ x[33];
  assign t[123] = t[179] ^ x[34];
  assign t[124] = t[180] ^ x[35];
  assign t[125] = t[181] ^ x[41];
  assign t[126] = t[182] ^ x[38];
  assign t[127] = t[183] ^ x[39];
  assign t[128] = t[184] ^ x[40];
  assign t[129] = t[185] ^ x[46];
  assign t[12] = ~t[21];
  assign t[130] = t[186] ^ x[43];
  assign t[131] = t[187] ^ x[44];
  assign t[132] = t[188] ^ x[45];
  assign t[133] = t[189] ^ x[51];
  assign t[134] = t[190] ^ x[48];
  assign t[135] = t[191] ^ x[49];
  assign t[136] = t[192] ^ x[50];
  assign t[137] = t[193] ^ x[56];
  assign t[138] = t[194] ^ x[53];
  assign t[139] = t[195] ^ x[54];
  assign t[13] = t[22] ^ t[23];
  assign t[140] = t[196] ^ x[55];
  assign t[141] = t[197] ^ x[61];
  assign t[142] = t[198] ^ x[58];
  assign t[143] = t[199] ^ x[59];
  assign t[144] = t[200] ^ x[60];
  assign t[145] = t[201] ^ x[66];
  assign t[146] = t[202] ^ x[63];
  assign t[147] = t[203] ^ x[64];
  assign t[148] = t[204] ^ x[65];
  assign t[149] = t[205] ^ x[71];
  assign t[14] = t[24] & t[25];
  assign t[150] = t[206] ^ x[68];
  assign t[151] = t[207] ^ x[69];
  assign t[152] = t[208] ^ x[70];
  assign t[153] = (x[2]);
  assign t[154] = (x[2]);
  assign t[155] = (x[2]);
  assign t[156] = (x[2]);
  assign t[157] = (x[7]);
  assign t[158] = (x[7]);
  assign t[159] = (x[7]);
  assign t[15] = t[26] ^ t[14];
  assign t[160] = (x[7]);
  assign t[161] = (x[12]);
  assign t[162] = (x[12]);
  assign t[163] = (x[12]);
  assign t[164] = (x[12]);
  assign t[165] = (x[17]);
  assign t[166] = (x[17]);
  assign t[167] = (x[17]);
  assign t[168] = (x[17]);
  assign t[169] = (x[22]);
  assign t[16] = t[57] ^ t[24];
  assign t[170] = (x[22]);
  assign t[171] = (x[22]);
  assign t[172] = (x[22]);
  assign t[173] = (x[27]);
  assign t[174] = (x[27]);
  assign t[175] = (x[27]);
  assign t[176] = (x[27]);
  assign t[177] = (x[32]);
  assign t[178] = (x[32]);
  assign t[179] = (x[32]);
  assign t[17] = t[27] ^ t[28];
  assign t[180] = (x[32]);
  assign t[181] = (x[37]);
  assign t[182] = (x[37]);
  assign t[183] = (x[37]);
  assign t[184] = (x[37]);
  assign t[185] = (x[42]);
  assign t[186] = (x[42]);
  assign t[187] = (x[42]);
  assign t[188] = (x[42]);
  assign t[189] = (x[47]);
  assign t[18] = t[29] & t[30];
  assign t[190] = (x[47]);
  assign t[191] = (x[47]);
  assign t[192] = (x[47]);
  assign t[193] = (x[52]);
  assign t[194] = (x[52]);
  assign t[195] = (x[52]);
  assign t[196] = (x[52]);
  assign t[197] = (x[57]);
  assign t[198] = (x[57]);
  assign t[199] = (x[57]);
  assign t[19] = t[31] ^ t[18];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[57]);
  assign t[201] = (x[62]);
  assign t[202] = (x[62]);
  assign t[203] = (x[62]);
  assign t[204] = (x[62]);
  assign t[205] = (x[67]);
  assign t[206] = (x[67]);
  assign t[207] = (x[67]);
  assign t[208] = (x[67]);
  assign t[20] = t[58] ^ t[29];
  assign t[21] = ~(t[32] ^ t[33]);
  assign t[22] = t[59] ^ t[60];
  assign t[23] = t[24] & t[34];
  assign t[24] = ~(t[60]);
  assign t[25] = ~(t[57] ^ t[24]);
  assign t[26] = t[57] & t[35];
  assign t[27] = t[61] ^ t[62];
  assign t[28] = t[29] & t[36];
  assign t[29] = ~(t[62]);
  assign t[2] = ~(t[4] ^ t[55]);
  assign t[30] = ~(t[58] ^ t[29]);
  assign t[31] = t[58] & t[37];
  assign t[32] = t[38] ^ t[39];
  assign t[33] = t[40] ^ t[41];
  assign t[34] = t[57] ^ t[42];
  assign t[35] = t[43] ^ t[23];
  assign t[36] = t[58] ^ t[44];
  assign t[37] = t[45] ^ t[28];
  assign t[38] = t[46] ^ t[47];
  assign t[39] = t[48] & t[49];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ t[39];
  assign t[41] = t[63] ^ t[48];
  assign t[42] = t[60] ^ t[64];
  assign t[43] = t[57] ^ t[22];
  assign t[44] = t[62] ^ t[65];
  assign t[45] = t[58] ^ t[27];
  assign t[46] = t[66] ^ t[67];
  assign t[47] = t[48] & t[51];
  assign t[48] = ~(t[67]);
  assign t[49] = ~(t[63] ^ t[48]);
  assign t[4] = ~t[7];
  assign t[50] = t[63] & t[52];
  assign t[51] = t[63] ^ t[53];
  assign t[52] = t[54] ^ t[47];
  assign t[53] = t[67] ^ t[68];
  assign t[54] = t[63] ^ t[46];
  assign t[55] = (t[69]);
  assign t[56] = (t[70]);
  assign t[57] = (t[71]);
  assign t[58] = (t[72]);
  assign t[59] = (t[73]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (t[74]);
  assign t[61] = (t[75]);
  assign t[62] = (t[76]);
  assign t[63] = (t[77]);
  assign t[64] = (t[78]);
  assign t[65] = (t[79]);
  assign t[66] = (t[80]);
  assign t[67] = (t[81]);
  assign t[68] = (t[82]);
  assign t[69] = t[83] ^ x[6];
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = t[84] ^ x[11];
  assign t[71] = t[85] ^ x[16];
  assign t[72] = t[86] ^ x[21];
  assign t[73] = t[87] ^ x[26];
  assign t[74] = t[88] ^ x[31];
  assign t[75] = t[89] ^ x[36];
  assign t[76] = t[90] ^ x[41];
  assign t[77] = t[91] ^ x[46];
  assign t[78] = t[92] ^ x[51];
  assign t[79] = t[93] ^ x[56];
  assign t[7] = ~(t[12] ^ t[56]);
  assign t[80] = t[94] ^ x[61];
  assign t[81] = t[95] ^ x[66];
  assign t[82] = t[96] ^ x[71];
  assign t[83] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[84] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[85] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[86] = (~t[109] & t[110] & t[111] & t[112]) | (t[109] & ~t[111] & ~t[112]) | (t[109] & ~t[110] & ~t[112]) | (t[109] & ~t[110] & ~t[111]);
  assign t[87] = (~t[113] & t[114] & t[115] & t[116]) | (t[113] & ~t[115] & ~t[116]) | (t[113] & ~t[114] & ~t[116]) | (t[113] & ~t[114] & ~t[115]);
  assign t[88] = (~t[117] & t[118] & t[119] & t[120]) | (t[117] & ~t[119] & ~t[120]) | (t[117] & ~t[118] & ~t[120]) | (t[117] & ~t[118] & ~t[119]);
  assign t[89] = (~t[121] & t[122] & t[123] & t[124]) | (t[121] & ~t[123] & ~t[124]) | (t[121] & ~t[122] & ~t[124]) | (t[121] & ~t[122] & ~t[123]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (~t[125] & t[126] & t[127] & t[128]) | (t[125] & ~t[127] & ~t[128]) | (t[125] & ~t[126] & ~t[128]) | (t[125] & ~t[126] & ~t[127]);
  assign t[91] = (~t[129] & t[130] & t[131] & t[132]) | (t[129] & ~t[131] & ~t[132]) | (t[129] & ~t[130] & ~t[132]) | (t[129] & ~t[130] & ~t[131]);
  assign t[92] = (~t[133] & t[134] & t[135] & t[136]) | (t[133] & ~t[135] & ~t[136]) | (t[133] & ~t[134] & ~t[136]) | (t[133] & ~t[134] & ~t[135]);
  assign t[93] = (~t[137] & t[138] & t[139] & t[140]) | (t[137] & ~t[139] & ~t[140]) | (t[137] & ~t[138] & ~t[140]) | (t[137] & ~t[138] & ~t[139]);
  assign t[94] = (~t[141] & t[142] & t[143] & t[144]) | (t[141] & ~t[143] & ~t[144]) | (t[141] & ~t[142] & ~t[144]) | (t[141] & ~t[142] & ~t[143]);
  assign t[95] = (~t[145] & t[146] & t[147] & t[148]) | (t[145] & ~t[147] & ~t[148]) | (t[145] & ~t[146] & ~t[148]) | (t[145] & ~t[146] & ~t[147]);
  assign t[96] = (~t[149] & t[150] & t[151] & t[152]) | (t[149] & ~t[151] & ~t[152]) | (t[149] & ~t[150] & ~t[152]) | (t[149] & ~t[150] & ~t[151]);
  assign t[97] = t[153] ^ x[6];
  assign t[98] = t[154] ^ x[3];
  assign t[99] = t[155] ^ x[4];
  assign t[9] = t[15] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind278(x, y);
 input [71:0] x;
 output y;

 wire [208:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[156] ^ x[5];
  assign t[101] = t[157] ^ x[11];
  assign t[102] = t[158] ^ x[8];
  assign t[103] = t[159] ^ x[9];
  assign t[104] = t[160] ^ x[10];
  assign t[105] = t[161] ^ x[16];
  assign t[106] = t[162] ^ x[13];
  assign t[107] = t[163] ^ x[14];
  assign t[108] = t[164] ^ x[15];
  assign t[109] = t[165] ^ x[21];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[166] ^ x[18];
  assign t[111] = t[167] ^ x[19];
  assign t[112] = t[168] ^ x[20];
  assign t[113] = t[169] ^ x[26];
  assign t[114] = t[170] ^ x[23];
  assign t[115] = t[171] ^ x[24];
  assign t[116] = t[172] ^ x[25];
  assign t[117] = t[173] ^ x[31];
  assign t[118] = t[174] ^ x[28];
  assign t[119] = t[175] ^ x[29];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[176] ^ x[30];
  assign t[121] = t[177] ^ x[36];
  assign t[122] = t[178] ^ x[33];
  assign t[123] = t[179] ^ x[34];
  assign t[124] = t[180] ^ x[35];
  assign t[125] = t[181] ^ x[41];
  assign t[126] = t[182] ^ x[38];
  assign t[127] = t[183] ^ x[39];
  assign t[128] = t[184] ^ x[40];
  assign t[129] = t[185] ^ x[46];
  assign t[12] = ~t[21];
  assign t[130] = t[186] ^ x[43];
  assign t[131] = t[187] ^ x[44];
  assign t[132] = t[188] ^ x[45];
  assign t[133] = t[189] ^ x[51];
  assign t[134] = t[190] ^ x[48];
  assign t[135] = t[191] ^ x[49];
  assign t[136] = t[192] ^ x[50];
  assign t[137] = t[193] ^ x[56];
  assign t[138] = t[194] ^ x[53];
  assign t[139] = t[195] ^ x[54];
  assign t[13] = t[22] ^ t[23];
  assign t[140] = t[196] ^ x[55];
  assign t[141] = t[197] ^ x[61];
  assign t[142] = t[198] ^ x[58];
  assign t[143] = t[199] ^ x[59];
  assign t[144] = t[200] ^ x[60];
  assign t[145] = t[201] ^ x[66];
  assign t[146] = t[202] ^ x[63];
  assign t[147] = t[203] ^ x[64];
  assign t[148] = t[204] ^ x[65];
  assign t[149] = t[205] ^ x[71];
  assign t[14] = t[24] & t[25];
  assign t[150] = t[206] ^ x[68];
  assign t[151] = t[207] ^ x[69];
  assign t[152] = t[208] ^ x[70];
  assign t[153] = (x[2]);
  assign t[154] = (x[2]);
  assign t[155] = (x[2]);
  assign t[156] = (x[2]);
  assign t[157] = (x[7]);
  assign t[158] = (x[7]);
  assign t[159] = (x[7]);
  assign t[15] = t[26] ^ t[14];
  assign t[160] = (x[7]);
  assign t[161] = (x[12]);
  assign t[162] = (x[12]);
  assign t[163] = (x[12]);
  assign t[164] = (x[12]);
  assign t[165] = (x[17]);
  assign t[166] = (x[17]);
  assign t[167] = (x[17]);
  assign t[168] = (x[17]);
  assign t[169] = (x[22]);
  assign t[16] = t[57] ^ t[24];
  assign t[170] = (x[22]);
  assign t[171] = (x[22]);
  assign t[172] = (x[22]);
  assign t[173] = (x[27]);
  assign t[174] = (x[27]);
  assign t[175] = (x[27]);
  assign t[176] = (x[27]);
  assign t[177] = (x[32]);
  assign t[178] = (x[32]);
  assign t[179] = (x[32]);
  assign t[17] = t[27] ^ t[28];
  assign t[180] = (x[32]);
  assign t[181] = (x[37]);
  assign t[182] = (x[37]);
  assign t[183] = (x[37]);
  assign t[184] = (x[37]);
  assign t[185] = (x[42]);
  assign t[186] = (x[42]);
  assign t[187] = (x[42]);
  assign t[188] = (x[42]);
  assign t[189] = (x[47]);
  assign t[18] = t[29] & t[30];
  assign t[190] = (x[47]);
  assign t[191] = (x[47]);
  assign t[192] = (x[47]);
  assign t[193] = (x[52]);
  assign t[194] = (x[52]);
  assign t[195] = (x[52]);
  assign t[196] = (x[52]);
  assign t[197] = (x[57]);
  assign t[198] = (x[57]);
  assign t[199] = (x[57]);
  assign t[19] = t[31] ^ t[18];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[57]);
  assign t[201] = (x[62]);
  assign t[202] = (x[62]);
  assign t[203] = (x[62]);
  assign t[204] = (x[62]);
  assign t[205] = (x[67]);
  assign t[206] = (x[67]);
  assign t[207] = (x[67]);
  assign t[208] = (x[67]);
  assign t[20] = t[58] ^ t[29];
  assign t[21] = ~(t[32] ^ t[33]);
  assign t[22] = t[59] ^ t[60];
  assign t[23] = t[24] & t[34];
  assign t[24] = ~(t[60]);
  assign t[25] = ~(t[57] ^ t[24]);
  assign t[26] = t[57] & t[35];
  assign t[27] = t[61] ^ t[62];
  assign t[28] = t[29] & t[36];
  assign t[29] = ~(t[62]);
  assign t[2] = ~(t[4] ^ t[55]);
  assign t[30] = ~(t[58] ^ t[29]);
  assign t[31] = t[58] & t[37];
  assign t[32] = t[38] ^ t[39];
  assign t[33] = t[40] ^ t[41];
  assign t[34] = t[57] ^ t[42];
  assign t[35] = t[43] ^ t[23];
  assign t[36] = t[58] ^ t[44];
  assign t[37] = t[45] ^ t[28];
  assign t[38] = t[46] ^ t[47];
  assign t[39] = t[48] & t[49];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ t[39];
  assign t[41] = t[63] ^ t[48];
  assign t[42] = t[60] ^ t[64];
  assign t[43] = t[57] ^ t[22];
  assign t[44] = t[62] ^ t[65];
  assign t[45] = t[58] ^ t[27];
  assign t[46] = t[66] ^ t[67];
  assign t[47] = t[48] & t[51];
  assign t[48] = ~(t[67]);
  assign t[49] = ~(t[63] ^ t[48]);
  assign t[4] = ~t[7];
  assign t[50] = t[63] & t[52];
  assign t[51] = t[63] ^ t[53];
  assign t[52] = t[54] ^ t[47];
  assign t[53] = t[67] ^ t[68];
  assign t[54] = t[63] ^ t[46];
  assign t[55] = (t[69]);
  assign t[56] = (t[70]);
  assign t[57] = (t[71]);
  assign t[58] = (t[72]);
  assign t[59] = (t[73]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (t[74]);
  assign t[61] = (t[75]);
  assign t[62] = (t[76]);
  assign t[63] = (t[77]);
  assign t[64] = (t[78]);
  assign t[65] = (t[79]);
  assign t[66] = (t[80]);
  assign t[67] = (t[81]);
  assign t[68] = (t[82]);
  assign t[69] = t[83] ^ x[6];
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = t[84] ^ x[11];
  assign t[71] = t[85] ^ x[16];
  assign t[72] = t[86] ^ x[21];
  assign t[73] = t[87] ^ x[26];
  assign t[74] = t[88] ^ x[31];
  assign t[75] = t[89] ^ x[36];
  assign t[76] = t[90] ^ x[41];
  assign t[77] = t[91] ^ x[46];
  assign t[78] = t[92] ^ x[51];
  assign t[79] = t[93] ^ x[56];
  assign t[7] = ~(t[12] ^ t[56]);
  assign t[80] = t[94] ^ x[61];
  assign t[81] = t[95] ^ x[66];
  assign t[82] = t[96] ^ x[71];
  assign t[83] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[84] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[85] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[86] = (~t[109] & t[110] & t[111] & t[112]) | (t[109] & ~t[111] & ~t[112]) | (t[109] & ~t[110] & ~t[112]) | (t[109] & ~t[110] & ~t[111]);
  assign t[87] = (~t[113] & t[114] & t[115] & t[116]) | (t[113] & ~t[115] & ~t[116]) | (t[113] & ~t[114] & ~t[116]) | (t[113] & ~t[114] & ~t[115]);
  assign t[88] = (~t[117] & t[118] & t[119] & t[120]) | (t[117] & ~t[119] & ~t[120]) | (t[117] & ~t[118] & ~t[120]) | (t[117] & ~t[118] & ~t[119]);
  assign t[89] = (~t[121] & t[122] & t[123] & t[124]) | (t[121] & ~t[123] & ~t[124]) | (t[121] & ~t[122] & ~t[124]) | (t[121] & ~t[122] & ~t[123]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (~t[125] & t[126] & t[127] & t[128]) | (t[125] & ~t[127] & ~t[128]) | (t[125] & ~t[126] & ~t[128]) | (t[125] & ~t[126] & ~t[127]);
  assign t[91] = (~t[129] & t[130] & t[131] & t[132]) | (t[129] & ~t[131] & ~t[132]) | (t[129] & ~t[130] & ~t[132]) | (t[129] & ~t[130] & ~t[131]);
  assign t[92] = (~t[133] & t[134] & t[135] & t[136]) | (t[133] & ~t[135] & ~t[136]) | (t[133] & ~t[134] & ~t[136]) | (t[133] & ~t[134] & ~t[135]);
  assign t[93] = (~t[137] & t[138] & t[139] & t[140]) | (t[137] & ~t[139] & ~t[140]) | (t[137] & ~t[138] & ~t[140]) | (t[137] & ~t[138] & ~t[139]);
  assign t[94] = (~t[141] & t[142] & t[143] & t[144]) | (t[141] & ~t[143] & ~t[144]) | (t[141] & ~t[142] & ~t[144]) | (t[141] & ~t[142] & ~t[143]);
  assign t[95] = (~t[145] & t[146] & t[147] & t[148]) | (t[145] & ~t[147] & ~t[148]) | (t[145] & ~t[146] & ~t[148]) | (t[145] & ~t[146] & ~t[147]);
  assign t[96] = (~t[149] & t[150] & t[151] & t[152]) | (t[149] & ~t[151] & ~t[152]) | (t[149] & ~t[150] & ~t[152]) | (t[149] & ~t[150] & ~t[151]);
  assign t[97] = t[153] ^ x[6];
  assign t[98] = t[154] ^ x[3];
  assign t[99] = t[155] ^ x[4];
  assign t[9] = t[15] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind279(x, y);
 input [71:0] x;
 output y;

 wire [208:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[156] ^ x[5];
  assign t[101] = t[157] ^ x[11];
  assign t[102] = t[158] ^ x[8];
  assign t[103] = t[159] ^ x[9];
  assign t[104] = t[160] ^ x[10];
  assign t[105] = t[161] ^ x[16];
  assign t[106] = t[162] ^ x[13];
  assign t[107] = t[163] ^ x[14];
  assign t[108] = t[164] ^ x[15];
  assign t[109] = t[165] ^ x[21];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[166] ^ x[18];
  assign t[111] = t[167] ^ x[19];
  assign t[112] = t[168] ^ x[20];
  assign t[113] = t[169] ^ x[26];
  assign t[114] = t[170] ^ x[23];
  assign t[115] = t[171] ^ x[24];
  assign t[116] = t[172] ^ x[25];
  assign t[117] = t[173] ^ x[31];
  assign t[118] = t[174] ^ x[28];
  assign t[119] = t[175] ^ x[29];
  assign t[11] = t[19] ^ t[20];
  assign t[120] = t[176] ^ x[30];
  assign t[121] = t[177] ^ x[36];
  assign t[122] = t[178] ^ x[33];
  assign t[123] = t[179] ^ x[34];
  assign t[124] = t[180] ^ x[35];
  assign t[125] = t[181] ^ x[41];
  assign t[126] = t[182] ^ x[38];
  assign t[127] = t[183] ^ x[39];
  assign t[128] = t[184] ^ x[40];
  assign t[129] = t[185] ^ x[46];
  assign t[12] = ~t[21];
  assign t[130] = t[186] ^ x[43];
  assign t[131] = t[187] ^ x[44];
  assign t[132] = t[188] ^ x[45];
  assign t[133] = t[189] ^ x[51];
  assign t[134] = t[190] ^ x[48];
  assign t[135] = t[191] ^ x[49];
  assign t[136] = t[192] ^ x[50];
  assign t[137] = t[193] ^ x[56];
  assign t[138] = t[194] ^ x[53];
  assign t[139] = t[195] ^ x[54];
  assign t[13] = t[22] ^ t[23];
  assign t[140] = t[196] ^ x[55];
  assign t[141] = t[197] ^ x[61];
  assign t[142] = t[198] ^ x[58];
  assign t[143] = t[199] ^ x[59];
  assign t[144] = t[200] ^ x[60];
  assign t[145] = t[201] ^ x[66];
  assign t[146] = t[202] ^ x[63];
  assign t[147] = t[203] ^ x[64];
  assign t[148] = t[204] ^ x[65];
  assign t[149] = t[205] ^ x[71];
  assign t[14] = t[24] & t[25];
  assign t[150] = t[206] ^ x[68];
  assign t[151] = t[207] ^ x[69];
  assign t[152] = t[208] ^ x[70];
  assign t[153] = (x[2]);
  assign t[154] = (x[2]);
  assign t[155] = (x[2]);
  assign t[156] = (x[2]);
  assign t[157] = (x[7]);
  assign t[158] = (x[7]);
  assign t[159] = (x[7]);
  assign t[15] = t[26] ^ t[14];
  assign t[160] = (x[7]);
  assign t[161] = (x[12]);
  assign t[162] = (x[12]);
  assign t[163] = (x[12]);
  assign t[164] = (x[12]);
  assign t[165] = (x[17]);
  assign t[166] = (x[17]);
  assign t[167] = (x[17]);
  assign t[168] = (x[17]);
  assign t[169] = (x[22]);
  assign t[16] = t[57] ^ t[24];
  assign t[170] = (x[22]);
  assign t[171] = (x[22]);
  assign t[172] = (x[22]);
  assign t[173] = (x[27]);
  assign t[174] = (x[27]);
  assign t[175] = (x[27]);
  assign t[176] = (x[27]);
  assign t[177] = (x[32]);
  assign t[178] = (x[32]);
  assign t[179] = (x[32]);
  assign t[17] = t[27] ^ t[28];
  assign t[180] = (x[32]);
  assign t[181] = (x[37]);
  assign t[182] = (x[37]);
  assign t[183] = (x[37]);
  assign t[184] = (x[37]);
  assign t[185] = (x[42]);
  assign t[186] = (x[42]);
  assign t[187] = (x[42]);
  assign t[188] = (x[42]);
  assign t[189] = (x[47]);
  assign t[18] = t[29] & t[30];
  assign t[190] = (x[47]);
  assign t[191] = (x[47]);
  assign t[192] = (x[47]);
  assign t[193] = (x[52]);
  assign t[194] = (x[52]);
  assign t[195] = (x[52]);
  assign t[196] = (x[52]);
  assign t[197] = (x[57]);
  assign t[198] = (x[57]);
  assign t[199] = (x[57]);
  assign t[19] = t[31] ^ t[18];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[57]);
  assign t[201] = (x[62]);
  assign t[202] = (x[62]);
  assign t[203] = (x[62]);
  assign t[204] = (x[62]);
  assign t[205] = (x[67]);
  assign t[206] = (x[67]);
  assign t[207] = (x[67]);
  assign t[208] = (x[67]);
  assign t[20] = t[58] ^ t[29];
  assign t[21] = ~(t[32] ^ t[33]);
  assign t[22] = t[59] ^ t[60];
  assign t[23] = t[24] & t[34];
  assign t[24] = ~(t[60]);
  assign t[25] = ~(t[57] ^ t[24]);
  assign t[26] = t[57] & t[35];
  assign t[27] = t[61] ^ t[62];
  assign t[28] = t[29] & t[36];
  assign t[29] = ~(t[62]);
  assign t[2] = ~(t[4] ^ t[55]);
  assign t[30] = ~(t[58] ^ t[29]);
  assign t[31] = t[58] & t[37];
  assign t[32] = t[38] ^ t[39];
  assign t[33] = t[40] ^ t[41];
  assign t[34] = t[57] ^ t[42];
  assign t[35] = t[43] ^ t[23];
  assign t[36] = t[58] ^ t[44];
  assign t[37] = t[45] ^ t[28];
  assign t[38] = t[46] ^ t[47];
  assign t[39] = t[48] & t[49];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ t[39];
  assign t[41] = t[63] ^ t[48];
  assign t[42] = t[60] ^ t[64];
  assign t[43] = t[57] ^ t[22];
  assign t[44] = t[62] ^ t[65];
  assign t[45] = t[58] ^ t[27];
  assign t[46] = t[66] ^ t[67];
  assign t[47] = t[48] & t[51];
  assign t[48] = ~(t[67]);
  assign t[49] = ~(t[63] ^ t[48]);
  assign t[4] = ~t[7];
  assign t[50] = t[63] & t[52];
  assign t[51] = t[63] ^ t[53];
  assign t[52] = t[54] ^ t[47];
  assign t[53] = t[67] ^ t[68];
  assign t[54] = t[63] ^ t[46];
  assign t[55] = (t[69]);
  assign t[56] = (t[70]);
  assign t[57] = (t[71]);
  assign t[58] = (t[72]);
  assign t[59] = (t[73]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (t[74]);
  assign t[61] = (t[75]);
  assign t[62] = (t[76]);
  assign t[63] = (t[77]);
  assign t[64] = (t[78]);
  assign t[65] = (t[79]);
  assign t[66] = (t[80]);
  assign t[67] = (t[81]);
  assign t[68] = (t[82]);
  assign t[69] = t[83] ^ x[6];
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = t[84] ^ x[11];
  assign t[71] = t[85] ^ x[16];
  assign t[72] = t[86] ^ x[21];
  assign t[73] = t[87] ^ x[26];
  assign t[74] = t[88] ^ x[31];
  assign t[75] = t[89] ^ x[36];
  assign t[76] = t[90] ^ x[41];
  assign t[77] = t[91] ^ x[46];
  assign t[78] = t[92] ^ x[51];
  assign t[79] = t[93] ^ x[56];
  assign t[7] = ~(t[12] ^ t[56]);
  assign t[80] = t[94] ^ x[61];
  assign t[81] = t[95] ^ x[66];
  assign t[82] = t[96] ^ x[71];
  assign t[83] = (~t[97] & t[98] & t[99] & t[100]) | (t[97] & ~t[99] & ~t[100]) | (t[97] & ~t[98] & ~t[100]) | (t[97] & ~t[98] & ~t[99]);
  assign t[84] = (~t[101] & t[102] & t[103] & t[104]) | (t[101] & ~t[103] & ~t[104]) | (t[101] & ~t[102] & ~t[104]) | (t[101] & ~t[102] & ~t[103]);
  assign t[85] = (~t[105] & t[106] & t[107] & t[108]) | (t[105] & ~t[107] & ~t[108]) | (t[105] & ~t[106] & ~t[108]) | (t[105] & ~t[106] & ~t[107]);
  assign t[86] = (~t[109] & t[110] & t[111] & t[112]) | (t[109] & ~t[111] & ~t[112]) | (t[109] & ~t[110] & ~t[112]) | (t[109] & ~t[110] & ~t[111]);
  assign t[87] = (~t[113] & t[114] & t[115] & t[116]) | (t[113] & ~t[115] & ~t[116]) | (t[113] & ~t[114] & ~t[116]) | (t[113] & ~t[114] & ~t[115]);
  assign t[88] = (~t[117] & t[118] & t[119] & t[120]) | (t[117] & ~t[119] & ~t[120]) | (t[117] & ~t[118] & ~t[120]) | (t[117] & ~t[118] & ~t[119]);
  assign t[89] = (~t[121] & t[122] & t[123] & t[124]) | (t[121] & ~t[123] & ~t[124]) | (t[121] & ~t[122] & ~t[124]) | (t[121] & ~t[122] & ~t[123]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (~t[125] & t[126] & t[127] & t[128]) | (t[125] & ~t[127] & ~t[128]) | (t[125] & ~t[126] & ~t[128]) | (t[125] & ~t[126] & ~t[127]);
  assign t[91] = (~t[129] & t[130] & t[131] & t[132]) | (t[129] & ~t[131] & ~t[132]) | (t[129] & ~t[130] & ~t[132]) | (t[129] & ~t[130] & ~t[131]);
  assign t[92] = (~t[133] & t[134] & t[135] & t[136]) | (t[133] & ~t[135] & ~t[136]) | (t[133] & ~t[134] & ~t[136]) | (t[133] & ~t[134] & ~t[135]);
  assign t[93] = (~t[137] & t[138] & t[139] & t[140]) | (t[137] & ~t[139] & ~t[140]) | (t[137] & ~t[138] & ~t[140]) | (t[137] & ~t[138] & ~t[139]);
  assign t[94] = (~t[141] & t[142] & t[143] & t[144]) | (t[141] & ~t[143] & ~t[144]) | (t[141] & ~t[142] & ~t[144]) | (t[141] & ~t[142] & ~t[143]);
  assign t[95] = (~t[145] & t[146] & t[147] & t[148]) | (t[145] & ~t[147] & ~t[148]) | (t[145] & ~t[146] & ~t[148]) | (t[145] & ~t[146] & ~t[147]);
  assign t[96] = (~t[149] & t[150] & t[151] & t[152]) | (t[149] & ~t[151] & ~t[152]) | (t[149] & ~t[150] & ~t[152]) | (t[149] & ~t[150] & ~t[151]);
  assign t[97] = t[153] ^ x[6];
  assign t[98] = t[154] ^ x[3];
  assign t[99] = t[155] ^ x[4];
  assign t[9] = t[15] ^ t[16];
  assign y = (t[0]);
endmodule

module R2ind280(x, y);
 input [56:0] x;
 output y;

 wire [145:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[144] ^ x[54];
  assign t[101] = t[145] ^ x[55];
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[2]);
  assign t[105] = (x[2]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[7]);
  assign t[109] = (x[7]);
  assign t[10] = ~t[15];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[12]);
  assign t[113] = (x[12]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[17]);
  assign t[117] = (x[17]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[27] ^ t[28];
  assign t[120] = (x[22]);
  assign t[121] = (x[22]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[27]);
  assign t[125] = (x[27]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[32]);
  assign t[129] = (x[32]);
  assign t[12] = t[16] & t[17];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[136] = (x[42]);
  assign t[137] = (x[42]);
  assign t[138] = (x[47]);
  assign t[139] = (x[47]);
  assign t[13] = t[29] ^ t[30];
  assign t[140] = (x[47]);
  assign t[141] = (x[47]);
  assign t[142] = (x[52]);
  assign t[143] = (x[52]);
  assign t[144] = (x[52]);
  assign t[145] = (x[52]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[20]);
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[31] ^ t[16]);
  assign t[18] = ~(t[29]);
  assign t[19] = ~(t[32] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] ^ t[22];
  assign t[21] = t[33] ^ t[34];
  assign t[22] = t[23] & t[24];
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[35] ^ t[23]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = ~(t[4] ^ t[25]);
  assign t[30] = (t[41]);
  assign t[31] = (t[42]);
  assign t[32] = (t[43]);
  assign t[33] = (t[44]);
  assign t[34] = (t[45]);
  assign t[35] = (t[46]);
  assign t[36] = t[47] ^ x[6];
  assign t[37] = t[48] ^ x[11];
  assign t[38] = t[49] ^ x[16];
  assign t[39] = t[50] ^ x[21];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[51] ^ x[26];
  assign t[41] = t[52] ^ x[31];
  assign t[42] = t[53] ^ x[36];
  assign t[43] = t[54] ^ x[41];
  assign t[44] = t[55] ^ x[46];
  assign t[45] = t[56] ^ x[51];
  assign t[46] = t[57] ^ x[56];
  assign t[47] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[48] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[49] = (~t[66] & t[67] & t[68] & t[69]) | (t[66] & ~t[68] & ~t[69]) | (t[66] & ~t[67] & ~t[69]) | (t[66] & ~t[67] & ~t[68]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[70] & t[71] & t[72] & t[73]) | (t[70] & ~t[72] & ~t[73]) | (t[70] & ~t[71] & ~t[73]) | (t[70] & ~t[71] & ~t[72]);
  assign t[51] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[52] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[53] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[54] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[55] = (~t[90] & t[91] & t[92] & t[93]) | (t[90] & ~t[92] & ~t[93]) | (t[90] & ~t[91] & ~t[93]) | (t[90] & ~t[91] & ~t[92]);
  assign t[56] = (~t[94] & t[95] & t[96] & t[97]) | (t[94] & ~t[96] & ~t[97]) | (t[94] & ~t[95] & ~t[97]) | (t[94] & ~t[95] & ~t[96]);
  assign t[57] = (~t[98] & t[99] & t[100] & t[101]) | (t[98] & ~t[100] & ~t[101]) | (t[98] & ~t[99] & ~t[101]) | (t[98] & ~t[99] & ~t[100]);
  assign t[58] = t[102] ^ x[6];
  assign t[59] = t[103] ^ x[3];
  assign t[5] = ~(t[8]);
  assign t[60] = t[104] ^ x[4];
  assign t[61] = t[105] ^ x[5];
  assign t[62] = t[106] ^ x[11];
  assign t[63] = t[107] ^ x[8];
  assign t[64] = t[108] ^ x[9];
  assign t[65] = t[109] ^ x[10];
  assign t[66] = t[110] ^ x[16];
  assign t[67] = t[111] ^ x[13];
  assign t[68] = t[112] ^ x[14];
  assign t[69] = t[113] ^ x[15];
  assign t[6] = ~(t[9]);
  assign t[70] = t[114] ^ x[21];
  assign t[71] = t[115] ^ x[18];
  assign t[72] = t[116] ^ x[19];
  assign t[73] = t[117] ^ x[20];
  assign t[74] = t[118] ^ x[26];
  assign t[75] = t[119] ^ x[23];
  assign t[76] = t[120] ^ x[24];
  assign t[77] = t[121] ^ x[25];
  assign t[78] = t[122] ^ x[31];
  assign t[79] = t[123] ^ x[28];
  assign t[7] = ~(t[10] ^ t[26]);
  assign t[80] = t[124] ^ x[29];
  assign t[81] = t[125] ^ x[30];
  assign t[82] = t[126] ^ x[36];
  assign t[83] = t[127] ^ x[33];
  assign t[84] = t[128] ^ x[34];
  assign t[85] = t[129] ^ x[35];
  assign t[86] = t[130] ^ x[41];
  assign t[87] = t[131] ^ x[38];
  assign t[88] = t[132] ^ x[39];
  assign t[89] = t[133] ^ x[40];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[134] ^ x[46];
  assign t[91] = t[135] ^ x[43];
  assign t[92] = t[136] ^ x[44];
  assign t[93] = t[137] ^ x[45];
  assign t[94] = t[138] ^ x[51];
  assign t[95] = t[139] ^ x[48];
  assign t[96] = t[140] ^ x[49];
  assign t[97] = t[141] ^ x[50];
  assign t[98] = t[142] ^ x[56];
  assign t[99] = t[143] ^ x[53];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind281(x, y);
 input [56:0] x;
 output y;

 wire [145:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[144] ^ x[54];
  assign t[101] = t[145] ^ x[55];
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[2]);
  assign t[105] = (x[2]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[7]);
  assign t[109] = (x[7]);
  assign t[10] = ~t[15];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[12]);
  assign t[113] = (x[12]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[17]);
  assign t[117] = (x[17]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[27] ^ t[28];
  assign t[120] = (x[22]);
  assign t[121] = (x[22]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[27]);
  assign t[125] = (x[27]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[32]);
  assign t[129] = (x[32]);
  assign t[12] = t[16] & t[17];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[136] = (x[42]);
  assign t[137] = (x[42]);
  assign t[138] = (x[47]);
  assign t[139] = (x[47]);
  assign t[13] = t[29] ^ t[30];
  assign t[140] = (x[47]);
  assign t[141] = (x[47]);
  assign t[142] = (x[52]);
  assign t[143] = (x[52]);
  assign t[144] = (x[52]);
  assign t[145] = (x[52]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[20]);
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[31] ^ t[16]);
  assign t[18] = ~(t[29]);
  assign t[19] = ~(t[32] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] ^ t[22];
  assign t[21] = t[33] ^ t[34];
  assign t[22] = t[23] & t[24];
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[35] ^ t[23]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = ~(t[4] ^ t[25]);
  assign t[30] = (t[41]);
  assign t[31] = (t[42]);
  assign t[32] = (t[43]);
  assign t[33] = (t[44]);
  assign t[34] = (t[45]);
  assign t[35] = (t[46]);
  assign t[36] = t[47] ^ x[6];
  assign t[37] = t[48] ^ x[11];
  assign t[38] = t[49] ^ x[16];
  assign t[39] = t[50] ^ x[21];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[51] ^ x[26];
  assign t[41] = t[52] ^ x[31];
  assign t[42] = t[53] ^ x[36];
  assign t[43] = t[54] ^ x[41];
  assign t[44] = t[55] ^ x[46];
  assign t[45] = t[56] ^ x[51];
  assign t[46] = t[57] ^ x[56];
  assign t[47] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[48] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[49] = (~t[66] & t[67] & t[68] & t[69]) | (t[66] & ~t[68] & ~t[69]) | (t[66] & ~t[67] & ~t[69]) | (t[66] & ~t[67] & ~t[68]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[70] & t[71] & t[72] & t[73]) | (t[70] & ~t[72] & ~t[73]) | (t[70] & ~t[71] & ~t[73]) | (t[70] & ~t[71] & ~t[72]);
  assign t[51] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[52] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[53] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[54] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[55] = (~t[90] & t[91] & t[92] & t[93]) | (t[90] & ~t[92] & ~t[93]) | (t[90] & ~t[91] & ~t[93]) | (t[90] & ~t[91] & ~t[92]);
  assign t[56] = (~t[94] & t[95] & t[96] & t[97]) | (t[94] & ~t[96] & ~t[97]) | (t[94] & ~t[95] & ~t[97]) | (t[94] & ~t[95] & ~t[96]);
  assign t[57] = (~t[98] & t[99] & t[100] & t[101]) | (t[98] & ~t[100] & ~t[101]) | (t[98] & ~t[99] & ~t[101]) | (t[98] & ~t[99] & ~t[100]);
  assign t[58] = t[102] ^ x[6];
  assign t[59] = t[103] ^ x[3];
  assign t[5] = ~(t[8]);
  assign t[60] = t[104] ^ x[4];
  assign t[61] = t[105] ^ x[5];
  assign t[62] = t[106] ^ x[11];
  assign t[63] = t[107] ^ x[8];
  assign t[64] = t[108] ^ x[9];
  assign t[65] = t[109] ^ x[10];
  assign t[66] = t[110] ^ x[16];
  assign t[67] = t[111] ^ x[13];
  assign t[68] = t[112] ^ x[14];
  assign t[69] = t[113] ^ x[15];
  assign t[6] = ~(t[9]);
  assign t[70] = t[114] ^ x[21];
  assign t[71] = t[115] ^ x[18];
  assign t[72] = t[116] ^ x[19];
  assign t[73] = t[117] ^ x[20];
  assign t[74] = t[118] ^ x[26];
  assign t[75] = t[119] ^ x[23];
  assign t[76] = t[120] ^ x[24];
  assign t[77] = t[121] ^ x[25];
  assign t[78] = t[122] ^ x[31];
  assign t[79] = t[123] ^ x[28];
  assign t[7] = ~(t[10] ^ t[26]);
  assign t[80] = t[124] ^ x[29];
  assign t[81] = t[125] ^ x[30];
  assign t[82] = t[126] ^ x[36];
  assign t[83] = t[127] ^ x[33];
  assign t[84] = t[128] ^ x[34];
  assign t[85] = t[129] ^ x[35];
  assign t[86] = t[130] ^ x[41];
  assign t[87] = t[131] ^ x[38];
  assign t[88] = t[132] ^ x[39];
  assign t[89] = t[133] ^ x[40];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[134] ^ x[46];
  assign t[91] = t[135] ^ x[43];
  assign t[92] = t[136] ^ x[44];
  assign t[93] = t[137] ^ x[45];
  assign t[94] = t[138] ^ x[51];
  assign t[95] = t[139] ^ x[48];
  assign t[96] = t[140] ^ x[49];
  assign t[97] = t[141] ^ x[50];
  assign t[98] = t[142] ^ x[56];
  assign t[99] = t[143] ^ x[53];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind282(x, y);
 input [56:0] x;
 output y;

 wire [145:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[144] ^ x[54];
  assign t[101] = t[145] ^ x[55];
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[2]);
  assign t[105] = (x[2]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[7]);
  assign t[109] = (x[7]);
  assign t[10] = ~t[15];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[12]);
  assign t[113] = (x[12]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[17]);
  assign t[117] = (x[17]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[27] ^ t[28];
  assign t[120] = (x[22]);
  assign t[121] = (x[22]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[27]);
  assign t[125] = (x[27]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[32]);
  assign t[129] = (x[32]);
  assign t[12] = t[16] & t[17];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[136] = (x[42]);
  assign t[137] = (x[42]);
  assign t[138] = (x[47]);
  assign t[139] = (x[47]);
  assign t[13] = t[29] ^ t[30];
  assign t[140] = (x[47]);
  assign t[141] = (x[47]);
  assign t[142] = (x[52]);
  assign t[143] = (x[52]);
  assign t[144] = (x[52]);
  assign t[145] = (x[52]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[20]);
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[31] ^ t[16]);
  assign t[18] = ~(t[29]);
  assign t[19] = ~(t[32] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] ^ t[22];
  assign t[21] = t[33] ^ t[34];
  assign t[22] = t[23] & t[24];
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[35] ^ t[23]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = ~(t[4] ^ t[25]);
  assign t[30] = (t[41]);
  assign t[31] = (t[42]);
  assign t[32] = (t[43]);
  assign t[33] = (t[44]);
  assign t[34] = (t[45]);
  assign t[35] = (t[46]);
  assign t[36] = t[47] ^ x[6];
  assign t[37] = t[48] ^ x[11];
  assign t[38] = t[49] ^ x[16];
  assign t[39] = t[50] ^ x[21];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[51] ^ x[26];
  assign t[41] = t[52] ^ x[31];
  assign t[42] = t[53] ^ x[36];
  assign t[43] = t[54] ^ x[41];
  assign t[44] = t[55] ^ x[46];
  assign t[45] = t[56] ^ x[51];
  assign t[46] = t[57] ^ x[56];
  assign t[47] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[48] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[49] = (~t[66] & t[67] & t[68] & t[69]) | (t[66] & ~t[68] & ~t[69]) | (t[66] & ~t[67] & ~t[69]) | (t[66] & ~t[67] & ~t[68]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[70] & t[71] & t[72] & t[73]) | (t[70] & ~t[72] & ~t[73]) | (t[70] & ~t[71] & ~t[73]) | (t[70] & ~t[71] & ~t[72]);
  assign t[51] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[52] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[53] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[54] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[55] = (~t[90] & t[91] & t[92] & t[93]) | (t[90] & ~t[92] & ~t[93]) | (t[90] & ~t[91] & ~t[93]) | (t[90] & ~t[91] & ~t[92]);
  assign t[56] = (~t[94] & t[95] & t[96] & t[97]) | (t[94] & ~t[96] & ~t[97]) | (t[94] & ~t[95] & ~t[97]) | (t[94] & ~t[95] & ~t[96]);
  assign t[57] = (~t[98] & t[99] & t[100] & t[101]) | (t[98] & ~t[100] & ~t[101]) | (t[98] & ~t[99] & ~t[101]) | (t[98] & ~t[99] & ~t[100]);
  assign t[58] = t[102] ^ x[6];
  assign t[59] = t[103] ^ x[3];
  assign t[5] = ~(t[8]);
  assign t[60] = t[104] ^ x[4];
  assign t[61] = t[105] ^ x[5];
  assign t[62] = t[106] ^ x[11];
  assign t[63] = t[107] ^ x[8];
  assign t[64] = t[108] ^ x[9];
  assign t[65] = t[109] ^ x[10];
  assign t[66] = t[110] ^ x[16];
  assign t[67] = t[111] ^ x[13];
  assign t[68] = t[112] ^ x[14];
  assign t[69] = t[113] ^ x[15];
  assign t[6] = ~(t[9]);
  assign t[70] = t[114] ^ x[21];
  assign t[71] = t[115] ^ x[18];
  assign t[72] = t[116] ^ x[19];
  assign t[73] = t[117] ^ x[20];
  assign t[74] = t[118] ^ x[26];
  assign t[75] = t[119] ^ x[23];
  assign t[76] = t[120] ^ x[24];
  assign t[77] = t[121] ^ x[25];
  assign t[78] = t[122] ^ x[31];
  assign t[79] = t[123] ^ x[28];
  assign t[7] = ~(t[10] ^ t[26]);
  assign t[80] = t[124] ^ x[29];
  assign t[81] = t[125] ^ x[30];
  assign t[82] = t[126] ^ x[36];
  assign t[83] = t[127] ^ x[33];
  assign t[84] = t[128] ^ x[34];
  assign t[85] = t[129] ^ x[35];
  assign t[86] = t[130] ^ x[41];
  assign t[87] = t[131] ^ x[38];
  assign t[88] = t[132] ^ x[39];
  assign t[89] = t[133] ^ x[40];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[134] ^ x[46];
  assign t[91] = t[135] ^ x[43];
  assign t[92] = t[136] ^ x[44];
  assign t[93] = t[137] ^ x[45];
  assign t[94] = t[138] ^ x[51];
  assign t[95] = t[139] ^ x[48];
  assign t[96] = t[140] ^ x[49];
  assign t[97] = t[141] ^ x[50];
  assign t[98] = t[142] ^ x[56];
  assign t[99] = t[143] ^ x[53];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind283(x, y);
 input [56:0] x;
 output y;

 wire [145:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[144] ^ x[54];
  assign t[101] = t[145] ^ x[55];
  assign t[102] = (x[2]);
  assign t[103] = (x[2]);
  assign t[104] = (x[2]);
  assign t[105] = (x[2]);
  assign t[106] = (x[7]);
  assign t[107] = (x[7]);
  assign t[108] = (x[7]);
  assign t[109] = (x[7]);
  assign t[10] = ~t[15];
  assign t[110] = (x[12]);
  assign t[111] = (x[12]);
  assign t[112] = (x[12]);
  assign t[113] = (x[12]);
  assign t[114] = (x[17]);
  assign t[115] = (x[17]);
  assign t[116] = (x[17]);
  assign t[117] = (x[17]);
  assign t[118] = (x[22]);
  assign t[119] = (x[22]);
  assign t[11] = t[27] ^ t[28];
  assign t[120] = (x[22]);
  assign t[121] = (x[22]);
  assign t[122] = (x[27]);
  assign t[123] = (x[27]);
  assign t[124] = (x[27]);
  assign t[125] = (x[27]);
  assign t[126] = (x[32]);
  assign t[127] = (x[32]);
  assign t[128] = (x[32]);
  assign t[129] = (x[32]);
  assign t[12] = t[16] & t[17];
  assign t[130] = (x[37]);
  assign t[131] = (x[37]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[42]);
  assign t[135] = (x[42]);
  assign t[136] = (x[42]);
  assign t[137] = (x[42]);
  assign t[138] = (x[47]);
  assign t[139] = (x[47]);
  assign t[13] = t[29] ^ t[30];
  assign t[140] = (x[47]);
  assign t[141] = (x[47]);
  assign t[142] = (x[52]);
  assign t[143] = (x[52]);
  assign t[144] = (x[52]);
  assign t[145] = (x[52]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[20]);
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[31] ^ t[16]);
  assign t[18] = ~(t[29]);
  assign t[19] = ~(t[32] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[21] ^ t[22];
  assign t[21] = t[33] ^ t[34];
  assign t[22] = t[23] & t[24];
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[35] ^ t[23]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = ~(t[4] ^ t[25]);
  assign t[30] = (t[41]);
  assign t[31] = (t[42]);
  assign t[32] = (t[43]);
  assign t[33] = (t[44]);
  assign t[34] = (t[45]);
  assign t[35] = (t[46]);
  assign t[36] = t[47] ^ x[6];
  assign t[37] = t[48] ^ x[11];
  assign t[38] = t[49] ^ x[16];
  assign t[39] = t[50] ^ x[21];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[51] ^ x[26];
  assign t[41] = t[52] ^ x[31];
  assign t[42] = t[53] ^ x[36];
  assign t[43] = t[54] ^ x[41];
  assign t[44] = t[55] ^ x[46];
  assign t[45] = t[56] ^ x[51];
  assign t[46] = t[57] ^ x[56];
  assign t[47] = (~t[58] & t[59] & t[60] & t[61]) | (t[58] & ~t[60] & ~t[61]) | (t[58] & ~t[59] & ~t[61]) | (t[58] & ~t[59] & ~t[60]);
  assign t[48] = (~t[62] & t[63] & t[64] & t[65]) | (t[62] & ~t[64] & ~t[65]) | (t[62] & ~t[63] & ~t[65]) | (t[62] & ~t[63] & ~t[64]);
  assign t[49] = (~t[66] & t[67] & t[68] & t[69]) | (t[66] & ~t[68] & ~t[69]) | (t[66] & ~t[67] & ~t[69]) | (t[66] & ~t[67] & ~t[68]);
  assign t[4] = ~t[7];
  assign t[50] = (~t[70] & t[71] & t[72] & t[73]) | (t[70] & ~t[72] & ~t[73]) | (t[70] & ~t[71] & ~t[73]) | (t[70] & ~t[71] & ~t[72]);
  assign t[51] = (~t[74] & t[75] & t[76] & t[77]) | (t[74] & ~t[76] & ~t[77]) | (t[74] & ~t[75] & ~t[77]) | (t[74] & ~t[75] & ~t[76]);
  assign t[52] = (~t[78] & t[79] & t[80] & t[81]) | (t[78] & ~t[80] & ~t[81]) | (t[78] & ~t[79] & ~t[81]) | (t[78] & ~t[79] & ~t[80]);
  assign t[53] = (~t[82] & t[83] & t[84] & t[85]) | (t[82] & ~t[84] & ~t[85]) | (t[82] & ~t[83] & ~t[85]) | (t[82] & ~t[83] & ~t[84]);
  assign t[54] = (~t[86] & t[87] & t[88] & t[89]) | (t[86] & ~t[88] & ~t[89]) | (t[86] & ~t[87] & ~t[89]) | (t[86] & ~t[87] & ~t[88]);
  assign t[55] = (~t[90] & t[91] & t[92] & t[93]) | (t[90] & ~t[92] & ~t[93]) | (t[90] & ~t[91] & ~t[93]) | (t[90] & ~t[91] & ~t[92]);
  assign t[56] = (~t[94] & t[95] & t[96] & t[97]) | (t[94] & ~t[96] & ~t[97]) | (t[94] & ~t[95] & ~t[97]) | (t[94] & ~t[95] & ~t[96]);
  assign t[57] = (~t[98] & t[99] & t[100] & t[101]) | (t[98] & ~t[100] & ~t[101]) | (t[98] & ~t[99] & ~t[101]) | (t[98] & ~t[99] & ~t[100]);
  assign t[58] = t[102] ^ x[6];
  assign t[59] = t[103] ^ x[3];
  assign t[5] = ~(t[8]);
  assign t[60] = t[104] ^ x[4];
  assign t[61] = t[105] ^ x[5];
  assign t[62] = t[106] ^ x[11];
  assign t[63] = t[107] ^ x[8];
  assign t[64] = t[108] ^ x[9];
  assign t[65] = t[109] ^ x[10];
  assign t[66] = t[110] ^ x[16];
  assign t[67] = t[111] ^ x[13];
  assign t[68] = t[112] ^ x[14];
  assign t[69] = t[113] ^ x[15];
  assign t[6] = ~(t[9]);
  assign t[70] = t[114] ^ x[21];
  assign t[71] = t[115] ^ x[18];
  assign t[72] = t[116] ^ x[19];
  assign t[73] = t[117] ^ x[20];
  assign t[74] = t[118] ^ x[26];
  assign t[75] = t[119] ^ x[23];
  assign t[76] = t[120] ^ x[24];
  assign t[77] = t[121] ^ x[25];
  assign t[78] = t[122] ^ x[31];
  assign t[79] = t[123] ^ x[28];
  assign t[7] = ~(t[10] ^ t[26]);
  assign t[80] = t[124] ^ x[29];
  assign t[81] = t[125] ^ x[30];
  assign t[82] = t[126] ^ x[36];
  assign t[83] = t[127] ^ x[33];
  assign t[84] = t[128] ^ x[34];
  assign t[85] = t[129] ^ x[35];
  assign t[86] = t[130] ^ x[41];
  assign t[87] = t[131] ^ x[38];
  assign t[88] = t[132] ^ x[39];
  assign t[89] = t[133] ^ x[40];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[134] ^ x[46];
  assign t[91] = t[135] ^ x[43];
  assign t[92] = t[136] ^ x[44];
  assign t[93] = t[137] ^ x[45];
  assign t[94] = t[138] ^ x[51];
  assign t[95] = t[139] ^ x[48];
  assign t[96] = t[140] ^ x[49];
  assign t[97] = t[141] ^ x[50];
  assign t[98] = t[142] ^ x[56];
  assign t[99] = t[143] ^ x[53];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind284(x, y);
 input [71:0] x;
 output y;

 wire [190:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[156] ^ x[28];
  assign t[101] = t[157] ^ x[29];
  assign t[102] = t[158] ^ x[30];
  assign t[103] = t[159] ^ x[36];
  assign t[104] = t[160] ^ x[33];
  assign t[105] = t[161] ^ x[34];
  assign t[106] = t[162] ^ x[35];
  assign t[107] = t[163] ^ x[41];
  assign t[108] = t[164] ^ x[38];
  assign t[109] = t[165] ^ x[39];
  assign t[10] = ~t[15];
  assign t[110] = t[166] ^ x[40];
  assign t[111] = t[167] ^ x[46];
  assign t[112] = t[168] ^ x[43];
  assign t[113] = t[169] ^ x[44];
  assign t[114] = t[170] ^ x[45];
  assign t[115] = t[171] ^ x[51];
  assign t[116] = t[172] ^ x[48];
  assign t[117] = t[173] ^ x[49];
  assign t[118] = t[174] ^ x[50];
  assign t[119] = t[175] ^ x[56];
  assign t[11] = t[16] ^ t[17];
  assign t[120] = t[176] ^ x[53];
  assign t[121] = t[177] ^ x[54];
  assign t[122] = t[178] ^ x[55];
  assign t[123] = t[179] ^ x[61];
  assign t[124] = t[180] ^ x[58];
  assign t[125] = t[181] ^ x[59];
  assign t[126] = t[182] ^ x[60];
  assign t[127] = t[183] ^ x[66];
  assign t[128] = t[184] ^ x[63];
  assign t[129] = t[185] ^ x[64];
  assign t[12] = t[18] & t[19];
  assign t[130] = t[186] ^ x[65];
  assign t[131] = t[187] ^ x[71];
  assign t[132] = t[188] ^ x[68];
  assign t[133] = t[189] ^ x[69];
  assign t[134] = t[190] ^ x[70];
  assign t[135] = (x[2]);
  assign t[136] = (x[2]);
  assign t[137] = (x[2]);
  assign t[138] = (x[2]);
  assign t[139] = (x[7]);
  assign t[13] = t[20] ^ t[21];
  assign t[140] = (x[7]);
  assign t[141] = (x[7]);
  assign t[142] = (x[7]);
  assign t[143] = (x[12]);
  assign t[144] = (x[12]);
  assign t[145] = (x[12]);
  assign t[146] = (x[12]);
  assign t[147] = (x[17]);
  assign t[148] = (x[17]);
  assign t[149] = (x[17]);
  assign t[14] = t[22] & t[23];
  assign t[150] = (x[17]);
  assign t[151] = (x[22]);
  assign t[152] = (x[22]);
  assign t[153] = (x[22]);
  assign t[154] = (x[22]);
  assign t[155] = (x[27]);
  assign t[156] = (x[27]);
  assign t[157] = (x[27]);
  assign t[158] = (x[27]);
  assign t[159] = (x[32]);
  assign t[15] = ~(t[24]);
  assign t[160] = (x[32]);
  assign t[161] = (x[32]);
  assign t[162] = (x[32]);
  assign t[163] = (x[37]);
  assign t[164] = (x[37]);
  assign t[165] = (x[37]);
  assign t[166] = (x[37]);
  assign t[167] = (x[42]);
  assign t[168] = (x[42]);
  assign t[169] = (x[42]);
  assign t[16] = t[39] ^ t[40];
  assign t[170] = (x[42]);
  assign t[171] = (x[47]);
  assign t[172] = (x[47]);
  assign t[173] = (x[47]);
  assign t[174] = (x[47]);
  assign t[175] = (x[52]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[52]);
  assign t[179] = (x[57]);
  assign t[17] = t[18] & t[25];
  assign t[180] = (x[57]);
  assign t[181] = (x[57]);
  assign t[182] = (x[57]);
  assign t[183] = (x[62]);
  assign t[184] = (x[62]);
  assign t[185] = (x[62]);
  assign t[186] = (x[62]);
  assign t[187] = (x[67]);
  assign t[188] = (x[67]);
  assign t[189] = (x[67]);
  assign t[18] = ~(t[40]);
  assign t[190] = (x[67]);
  assign t[19] = ~(t[41] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[42] ^ t[43];
  assign t[21] = t[22] & t[26];
  assign t[22] = ~(t[43]);
  assign t[23] = ~(t[44] ^ t[22]);
  assign t[24] = t[27] ^ t[28];
  assign t[25] = t[41] ^ t[29];
  assign t[26] = t[44] ^ t[30];
  assign t[27] = t[31] ^ t[32];
  assign t[28] = t[33] & t[34];
  assign t[29] = t[40] ^ t[45];
  assign t[2] = ~(t[4] ^ t[37]);
  assign t[30] = t[43] ^ t[46];
  assign t[31] = t[47] ^ t[48];
  assign t[32] = t[33] & t[35];
  assign t[33] = ~(t[48]);
  assign t[34] = ~(t[49] ^ t[33]);
  assign t[35] = t[49] ^ t[36];
  assign t[36] = t[48] ^ t[50];
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = (t[57]);
  assign t[44] = (t[58]);
  assign t[45] = (t[59]);
  assign t[46] = (t[60]);
  assign t[47] = (t[61]);
  assign t[48] = (t[62]);
  assign t[49] = (t[63]);
  assign t[4] = ~t[7];
  assign t[50] = (t[64]);
  assign t[51] = t[65] ^ x[6];
  assign t[52] = t[66] ^ x[11];
  assign t[53] = t[67] ^ x[16];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[26];
  assign t[56] = t[70] ^ x[31];
  assign t[57] = t[71] ^ x[36];
  assign t[58] = t[72] ^ x[41];
  assign t[59] = t[73] ^ x[46];
  assign t[5] = ~(t[8]);
  assign t[60] = t[74] ^ x[51];
  assign t[61] = t[75] ^ x[56];
  assign t[62] = t[76] ^ x[61];
  assign t[63] = t[77] ^ x[66];
  assign t[64] = t[78] ^ x[71];
  assign t[65] = (~t[79] & t[80] & t[81] & t[82]) | (t[79] & ~t[81] & ~t[82]) | (t[79] & ~t[80] & ~t[82]) | (t[79] & ~t[80] & ~t[81]);
  assign t[66] = (~t[83] & t[84] & t[85] & t[86]) | (t[83] & ~t[85] & ~t[86]) | (t[83] & ~t[84] & ~t[86]) | (t[83] & ~t[84] & ~t[85]);
  assign t[67] = (~t[87] & t[88] & t[89] & t[90]) | (t[87] & ~t[89] & ~t[90]) | (t[87] & ~t[88] & ~t[90]) | (t[87] & ~t[88] & ~t[89]);
  assign t[68] = (~t[91] & t[92] & t[93] & t[94]) | (t[91] & ~t[93] & ~t[94]) | (t[91] & ~t[92] & ~t[94]) | (t[91] & ~t[92] & ~t[93]);
  assign t[69] = (~t[95] & t[96] & t[97] & t[98]) | (t[95] & ~t[97] & ~t[98]) | (t[95] & ~t[96] & ~t[98]) | (t[95] & ~t[96] & ~t[97]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[99] & t[100] & t[101] & t[102]) | (t[99] & ~t[101] & ~t[102]) | (t[99] & ~t[100] & ~t[102]) | (t[99] & ~t[100] & ~t[101]);
  assign t[71] = (~t[103] & t[104] & t[105] & t[106]) | (t[103] & ~t[105] & ~t[106]) | (t[103] & ~t[104] & ~t[106]) | (t[103] & ~t[104] & ~t[105]);
  assign t[72] = (~t[107] & t[108] & t[109] & t[110]) | (t[107] & ~t[109] & ~t[110]) | (t[107] & ~t[108] & ~t[110]) | (t[107] & ~t[108] & ~t[109]);
  assign t[73] = (~t[111] & t[112] & t[113] & t[114]) | (t[111] & ~t[113] & ~t[114]) | (t[111] & ~t[112] & ~t[114]) | (t[111] & ~t[112] & ~t[113]);
  assign t[74] = (~t[115] & t[116] & t[117] & t[118]) | (t[115] & ~t[117] & ~t[118]) | (t[115] & ~t[116] & ~t[118]) | (t[115] & ~t[116] & ~t[117]);
  assign t[75] = (~t[119] & t[120] & t[121] & t[122]) | (t[119] & ~t[121] & ~t[122]) | (t[119] & ~t[120] & ~t[122]) | (t[119] & ~t[120] & ~t[121]);
  assign t[76] = (~t[123] & t[124] & t[125] & t[126]) | (t[123] & ~t[125] & ~t[126]) | (t[123] & ~t[124] & ~t[126]) | (t[123] & ~t[124] & ~t[125]);
  assign t[77] = (~t[127] & t[128] & t[129] & t[130]) | (t[127] & ~t[129] & ~t[130]) | (t[127] & ~t[128] & ~t[130]) | (t[127] & ~t[128] & ~t[129]);
  assign t[78] = (~t[131] & t[132] & t[133] & t[134]) | (t[131] & ~t[133] & ~t[134]) | (t[131] & ~t[132] & ~t[134]) | (t[131] & ~t[132] & ~t[133]);
  assign t[79] = t[135] ^ x[6];
  assign t[7] = ~(t[10] ^ t[38]);
  assign t[80] = t[136] ^ x[3];
  assign t[81] = t[137] ^ x[4];
  assign t[82] = t[138] ^ x[5];
  assign t[83] = t[139] ^ x[11];
  assign t[84] = t[140] ^ x[8];
  assign t[85] = t[141] ^ x[9];
  assign t[86] = t[142] ^ x[10];
  assign t[87] = t[143] ^ x[16];
  assign t[88] = t[144] ^ x[13];
  assign t[89] = t[145] ^ x[14];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[146] ^ x[15];
  assign t[91] = t[147] ^ x[21];
  assign t[92] = t[148] ^ x[18];
  assign t[93] = t[149] ^ x[19];
  assign t[94] = t[150] ^ x[20];
  assign t[95] = t[151] ^ x[26];
  assign t[96] = t[152] ^ x[23];
  assign t[97] = t[153] ^ x[24];
  assign t[98] = t[154] ^ x[25];
  assign t[99] = t[155] ^ x[31];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind285(x, y);
 input [71:0] x;
 output y;

 wire [190:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[156] ^ x[28];
  assign t[101] = t[157] ^ x[29];
  assign t[102] = t[158] ^ x[30];
  assign t[103] = t[159] ^ x[36];
  assign t[104] = t[160] ^ x[33];
  assign t[105] = t[161] ^ x[34];
  assign t[106] = t[162] ^ x[35];
  assign t[107] = t[163] ^ x[41];
  assign t[108] = t[164] ^ x[38];
  assign t[109] = t[165] ^ x[39];
  assign t[10] = ~t[15];
  assign t[110] = t[166] ^ x[40];
  assign t[111] = t[167] ^ x[46];
  assign t[112] = t[168] ^ x[43];
  assign t[113] = t[169] ^ x[44];
  assign t[114] = t[170] ^ x[45];
  assign t[115] = t[171] ^ x[51];
  assign t[116] = t[172] ^ x[48];
  assign t[117] = t[173] ^ x[49];
  assign t[118] = t[174] ^ x[50];
  assign t[119] = t[175] ^ x[56];
  assign t[11] = t[16] ^ t[17];
  assign t[120] = t[176] ^ x[53];
  assign t[121] = t[177] ^ x[54];
  assign t[122] = t[178] ^ x[55];
  assign t[123] = t[179] ^ x[61];
  assign t[124] = t[180] ^ x[58];
  assign t[125] = t[181] ^ x[59];
  assign t[126] = t[182] ^ x[60];
  assign t[127] = t[183] ^ x[66];
  assign t[128] = t[184] ^ x[63];
  assign t[129] = t[185] ^ x[64];
  assign t[12] = t[18] & t[19];
  assign t[130] = t[186] ^ x[65];
  assign t[131] = t[187] ^ x[71];
  assign t[132] = t[188] ^ x[68];
  assign t[133] = t[189] ^ x[69];
  assign t[134] = t[190] ^ x[70];
  assign t[135] = (x[2]);
  assign t[136] = (x[2]);
  assign t[137] = (x[2]);
  assign t[138] = (x[2]);
  assign t[139] = (x[7]);
  assign t[13] = t[20] ^ t[21];
  assign t[140] = (x[7]);
  assign t[141] = (x[7]);
  assign t[142] = (x[7]);
  assign t[143] = (x[12]);
  assign t[144] = (x[12]);
  assign t[145] = (x[12]);
  assign t[146] = (x[12]);
  assign t[147] = (x[17]);
  assign t[148] = (x[17]);
  assign t[149] = (x[17]);
  assign t[14] = t[22] & t[23];
  assign t[150] = (x[17]);
  assign t[151] = (x[22]);
  assign t[152] = (x[22]);
  assign t[153] = (x[22]);
  assign t[154] = (x[22]);
  assign t[155] = (x[27]);
  assign t[156] = (x[27]);
  assign t[157] = (x[27]);
  assign t[158] = (x[27]);
  assign t[159] = (x[32]);
  assign t[15] = ~(t[24]);
  assign t[160] = (x[32]);
  assign t[161] = (x[32]);
  assign t[162] = (x[32]);
  assign t[163] = (x[37]);
  assign t[164] = (x[37]);
  assign t[165] = (x[37]);
  assign t[166] = (x[37]);
  assign t[167] = (x[42]);
  assign t[168] = (x[42]);
  assign t[169] = (x[42]);
  assign t[16] = t[39] ^ t[40];
  assign t[170] = (x[42]);
  assign t[171] = (x[47]);
  assign t[172] = (x[47]);
  assign t[173] = (x[47]);
  assign t[174] = (x[47]);
  assign t[175] = (x[52]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[52]);
  assign t[179] = (x[57]);
  assign t[17] = t[18] & t[25];
  assign t[180] = (x[57]);
  assign t[181] = (x[57]);
  assign t[182] = (x[57]);
  assign t[183] = (x[62]);
  assign t[184] = (x[62]);
  assign t[185] = (x[62]);
  assign t[186] = (x[62]);
  assign t[187] = (x[67]);
  assign t[188] = (x[67]);
  assign t[189] = (x[67]);
  assign t[18] = ~(t[40]);
  assign t[190] = (x[67]);
  assign t[19] = ~(t[41] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[42] ^ t[43];
  assign t[21] = t[22] & t[26];
  assign t[22] = ~(t[43]);
  assign t[23] = ~(t[44] ^ t[22]);
  assign t[24] = t[27] ^ t[28];
  assign t[25] = t[41] ^ t[29];
  assign t[26] = t[44] ^ t[30];
  assign t[27] = t[31] ^ t[32];
  assign t[28] = t[33] & t[34];
  assign t[29] = t[40] ^ t[45];
  assign t[2] = ~(t[4] ^ t[37]);
  assign t[30] = t[43] ^ t[46];
  assign t[31] = t[47] ^ t[48];
  assign t[32] = t[33] & t[35];
  assign t[33] = ~(t[48]);
  assign t[34] = ~(t[49] ^ t[33]);
  assign t[35] = t[49] ^ t[36];
  assign t[36] = t[48] ^ t[50];
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = (t[57]);
  assign t[44] = (t[58]);
  assign t[45] = (t[59]);
  assign t[46] = (t[60]);
  assign t[47] = (t[61]);
  assign t[48] = (t[62]);
  assign t[49] = (t[63]);
  assign t[4] = ~t[7];
  assign t[50] = (t[64]);
  assign t[51] = t[65] ^ x[6];
  assign t[52] = t[66] ^ x[11];
  assign t[53] = t[67] ^ x[16];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[26];
  assign t[56] = t[70] ^ x[31];
  assign t[57] = t[71] ^ x[36];
  assign t[58] = t[72] ^ x[41];
  assign t[59] = t[73] ^ x[46];
  assign t[5] = ~(t[8]);
  assign t[60] = t[74] ^ x[51];
  assign t[61] = t[75] ^ x[56];
  assign t[62] = t[76] ^ x[61];
  assign t[63] = t[77] ^ x[66];
  assign t[64] = t[78] ^ x[71];
  assign t[65] = (~t[79] & t[80] & t[81] & t[82]) | (t[79] & ~t[81] & ~t[82]) | (t[79] & ~t[80] & ~t[82]) | (t[79] & ~t[80] & ~t[81]);
  assign t[66] = (~t[83] & t[84] & t[85] & t[86]) | (t[83] & ~t[85] & ~t[86]) | (t[83] & ~t[84] & ~t[86]) | (t[83] & ~t[84] & ~t[85]);
  assign t[67] = (~t[87] & t[88] & t[89] & t[90]) | (t[87] & ~t[89] & ~t[90]) | (t[87] & ~t[88] & ~t[90]) | (t[87] & ~t[88] & ~t[89]);
  assign t[68] = (~t[91] & t[92] & t[93] & t[94]) | (t[91] & ~t[93] & ~t[94]) | (t[91] & ~t[92] & ~t[94]) | (t[91] & ~t[92] & ~t[93]);
  assign t[69] = (~t[95] & t[96] & t[97] & t[98]) | (t[95] & ~t[97] & ~t[98]) | (t[95] & ~t[96] & ~t[98]) | (t[95] & ~t[96] & ~t[97]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[99] & t[100] & t[101] & t[102]) | (t[99] & ~t[101] & ~t[102]) | (t[99] & ~t[100] & ~t[102]) | (t[99] & ~t[100] & ~t[101]);
  assign t[71] = (~t[103] & t[104] & t[105] & t[106]) | (t[103] & ~t[105] & ~t[106]) | (t[103] & ~t[104] & ~t[106]) | (t[103] & ~t[104] & ~t[105]);
  assign t[72] = (~t[107] & t[108] & t[109] & t[110]) | (t[107] & ~t[109] & ~t[110]) | (t[107] & ~t[108] & ~t[110]) | (t[107] & ~t[108] & ~t[109]);
  assign t[73] = (~t[111] & t[112] & t[113] & t[114]) | (t[111] & ~t[113] & ~t[114]) | (t[111] & ~t[112] & ~t[114]) | (t[111] & ~t[112] & ~t[113]);
  assign t[74] = (~t[115] & t[116] & t[117] & t[118]) | (t[115] & ~t[117] & ~t[118]) | (t[115] & ~t[116] & ~t[118]) | (t[115] & ~t[116] & ~t[117]);
  assign t[75] = (~t[119] & t[120] & t[121] & t[122]) | (t[119] & ~t[121] & ~t[122]) | (t[119] & ~t[120] & ~t[122]) | (t[119] & ~t[120] & ~t[121]);
  assign t[76] = (~t[123] & t[124] & t[125] & t[126]) | (t[123] & ~t[125] & ~t[126]) | (t[123] & ~t[124] & ~t[126]) | (t[123] & ~t[124] & ~t[125]);
  assign t[77] = (~t[127] & t[128] & t[129] & t[130]) | (t[127] & ~t[129] & ~t[130]) | (t[127] & ~t[128] & ~t[130]) | (t[127] & ~t[128] & ~t[129]);
  assign t[78] = (~t[131] & t[132] & t[133] & t[134]) | (t[131] & ~t[133] & ~t[134]) | (t[131] & ~t[132] & ~t[134]) | (t[131] & ~t[132] & ~t[133]);
  assign t[79] = t[135] ^ x[6];
  assign t[7] = ~(t[10] ^ t[38]);
  assign t[80] = t[136] ^ x[3];
  assign t[81] = t[137] ^ x[4];
  assign t[82] = t[138] ^ x[5];
  assign t[83] = t[139] ^ x[11];
  assign t[84] = t[140] ^ x[8];
  assign t[85] = t[141] ^ x[9];
  assign t[86] = t[142] ^ x[10];
  assign t[87] = t[143] ^ x[16];
  assign t[88] = t[144] ^ x[13];
  assign t[89] = t[145] ^ x[14];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[146] ^ x[15];
  assign t[91] = t[147] ^ x[21];
  assign t[92] = t[148] ^ x[18];
  assign t[93] = t[149] ^ x[19];
  assign t[94] = t[150] ^ x[20];
  assign t[95] = t[151] ^ x[26];
  assign t[96] = t[152] ^ x[23];
  assign t[97] = t[153] ^ x[24];
  assign t[98] = t[154] ^ x[25];
  assign t[99] = t[155] ^ x[31];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind286(x, y);
 input [71:0] x;
 output y;

 wire [190:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[156] ^ x[28];
  assign t[101] = t[157] ^ x[29];
  assign t[102] = t[158] ^ x[30];
  assign t[103] = t[159] ^ x[36];
  assign t[104] = t[160] ^ x[33];
  assign t[105] = t[161] ^ x[34];
  assign t[106] = t[162] ^ x[35];
  assign t[107] = t[163] ^ x[41];
  assign t[108] = t[164] ^ x[38];
  assign t[109] = t[165] ^ x[39];
  assign t[10] = ~t[15];
  assign t[110] = t[166] ^ x[40];
  assign t[111] = t[167] ^ x[46];
  assign t[112] = t[168] ^ x[43];
  assign t[113] = t[169] ^ x[44];
  assign t[114] = t[170] ^ x[45];
  assign t[115] = t[171] ^ x[51];
  assign t[116] = t[172] ^ x[48];
  assign t[117] = t[173] ^ x[49];
  assign t[118] = t[174] ^ x[50];
  assign t[119] = t[175] ^ x[56];
  assign t[11] = t[16] ^ t[17];
  assign t[120] = t[176] ^ x[53];
  assign t[121] = t[177] ^ x[54];
  assign t[122] = t[178] ^ x[55];
  assign t[123] = t[179] ^ x[61];
  assign t[124] = t[180] ^ x[58];
  assign t[125] = t[181] ^ x[59];
  assign t[126] = t[182] ^ x[60];
  assign t[127] = t[183] ^ x[66];
  assign t[128] = t[184] ^ x[63];
  assign t[129] = t[185] ^ x[64];
  assign t[12] = t[18] & t[19];
  assign t[130] = t[186] ^ x[65];
  assign t[131] = t[187] ^ x[71];
  assign t[132] = t[188] ^ x[68];
  assign t[133] = t[189] ^ x[69];
  assign t[134] = t[190] ^ x[70];
  assign t[135] = (x[2]);
  assign t[136] = (x[2]);
  assign t[137] = (x[2]);
  assign t[138] = (x[2]);
  assign t[139] = (x[7]);
  assign t[13] = t[20] ^ t[21];
  assign t[140] = (x[7]);
  assign t[141] = (x[7]);
  assign t[142] = (x[7]);
  assign t[143] = (x[12]);
  assign t[144] = (x[12]);
  assign t[145] = (x[12]);
  assign t[146] = (x[12]);
  assign t[147] = (x[17]);
  assign t[148] = (x[17]);
  assign t[149] = (x[17]);
  assign t[14] = t[22] & t[23];
  assign t[150] = (x[17]);
  assign t[151] = (x[22]);
  assign t[152] = (x[22]);
  assign t[153] = (x[22]);
  assign t[154] = (x[22]);
  assign t[155] = (x[27]);
  assign t[156] = (x[27]);
  assign t[157] = (x[27]);
  assign t[158] = (x[27]);
  assign t[159] = (x[32]);
  assign t[15] = ~(t[24]);
  assign t[160] = (x[32]);
  assign t[161] = (x[32]);
  assign t[162] = (x[32]);
  assign t[163] = (x[37]);
  assign t[164] = (x[37]);
  assign t[165] = (x[37]);
  assign t[166] = (x[37]);
  assign t[167] = (x[42]);
  assign t[168] = (x[42]);
  assign t[169] = (x[42]);
  assign t[16] = t[39] ^ t[40];
  assign t[170] = (x[42]);
  assign t[171] = (x[47]);
  assign t[172] = (x[47]);
  assign t[173] = (x[47]);
  assign t[174] = (x[47]);
  assign t[175] = (x[52]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[52]);
  assign t[179] = (x[57]);
  assign t[17] = t[18] & t[25];
  assign t[180] = (x[57]);
  assign t[181] = (x[57]);
  assign t[182] = (x[57]);
  assign t[183] = (x[62]);
  assign t[184] = (x[62]);
  assign t[185] = (x[62]);
  assign t[186] = (x[62]);
  assign t[187] = (x[67]);
  assign t[188] = (x[67]);
  assign t[189] = (x[67]);
  assign t[18] = ~(t[40]);
  assign t[190] = (x[67]);
  assign t[19] = ~(t[41] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[42] ^ t[43];
  assign t[21] = t[22] & t[26];
  assign t[22] = ~(t[43]);
  assign t[23] = ~(t[44] ^ t[22]);
  assign t[24] = t[27] ^ t[28];
  assign t[25] = t[41] ^ t[29];
  assign t[26] = t[44] ^ t[30];
  assign t[27] = t[31] ^ t[32];
  assign t[28] = t[33] & t[34];
  assign t[29] = t[40] ^ t[45];
  assign t[2] = ~(t[4] ^ t[37]);
  assign t[30] = t[43] ^ t[46];
  assign t[31] = t[47] ^ t[48];
  assign t[32] = t[33] & t[35];
  assign t[33] = ~(t[48]);
  assign t[34] = ~(t[49] ^ t[33]);
  assign t[35] = t[49] ^ t[36];
  assign t[36] = t[48] ^ t[50];
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = (t[57]);
  assign t[44] = (t[58]);
  assign t[45] = (t[59]);
  assign t[46] = (t[60]);
  assign t[47] = (t[61]);
  assign t[48] = (t[62]);
  assign t[49] = (t[63]);
  assign t[4] = ~t[7];
  assign t[50] = (t[64]);
  assign t[51] = t[65] ^ x[6];
  assign t[52] = t[66] ^ x[11];
  assign t[53] = t[67] ^ x[16];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[26];
  assign t[56] = t[70] ^ x[31];
  assign t[57] = t[71] ^ x[36];
  assign t[58] = t[72] ^ x[41];
  assign t[59] = t[73] ^ x[46];
  assign t[5] = ~(t[8]);
  assign t[60] = t[74] ^ x[51];
  assign t[61] = t[75] ^ x[56];
  assign t[62] = t[76] ^ x[61];
  assign t[63] = t[77] ^ x[66];
  assign t[64] = t[78] ^ x[71];
  assign t[65] = (~t[79] & t[80] & t[81] & t[82]) | (t[79] & ~t[81] & ~t[82]) | (t[79] & ~t[80] & ~t[82]) | (t[79] & ~t[80] & ~t[81]);
  assign t[66] = (~t[83] & t[84] & t[85] & t[86]) | (t[83] & ~t[85] & ~t[86]) | (t[83] & ~t[84] & ~t[86]) | (t[83] & ~t[84] & ~t[85]);
  assign t[67] = (~t[87] & t[88] & t[89] & t[90]) | (t[87] & ~t[89] & ~t[90]) | (t[87] & ~t[88] & ~t[90]) | (t[87] & ~t[88] & ~t[89]);
  assign t[68] = (~t[91] & t[92] & t[93] & t[94]) | (t[91] & ~t[93] & ~t[94]) | (t[91] & ~t[92] & ~t[94]) | (t[91] & ~t[92] & ~t[93]);
  assign t[69] = (~t[95] & t[96] & t[97] & t[98]) | (t[95] & ~t[97] & ~t[98]) | (t[95] & ~t[96] & ~t[98]) | (t[95] & ~t[96] & ~t[97]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[99] & t[100] & t[101] & t[102]) | (t[99] & ~t[101] & ~t[102]) | (t[99] & ~t[100] & ~t[102]) | (t[99] & ~t[100] & ~t[101]);
  assign t[71] = (~t[103] & t[104] & t[105] & t[106]) | (t[103] & ~t[105] & ~t[106]) | (t[103] & ~t[104] & ~t[106]) | (t[103] & ~t[104] & ~t[105]);
  assign t[72] = (~t[107] & t[108] & t[109] & t[110]) | (t[107] & ~t[109] & ~t[110]) | (t[107] & ~t[108] & ~t[110]) | (t[107] & ~t[108] & ~t[109]);
  assign t[73] = (~t[111] & t[112] & t[113] & t[114]) | (t[111] & ~t[113] & ~t[114]) | (t[111] & ~t[112] & ~t[114]) | (t[111] & ~t[112] & ~t[113]);
  assign t[74] = (~t[115] & t[116] & t[117] & t[118]) | (t[115] & ~t[117] & ~t[118]) | (t[115] & ~t[116] & ~t[118]) | (t[115] & ~t[116] & ~t[117]);
  assign t[75] = (~t[119] & t[120] & t[121] & t[122]) | (t[119] & ~t[121] & ~t[122]) | (t[119] & ~t[120] & ~t[122]) | (t[119] & ~t[120] & ~t[121]);
  assign t[76] = (~t[123] & t[124] & t[125] & t[126]) | (t[123] & ~t[125] & ~t[126]) | (t[123] & ~t[124] & ~t[126]) | (t[123] & ~t[124] & ~t[125]);
  assign t[77] = (~t[127] & t[128] & t[129] & t[130]) | (t[127] & ~t[129] & ~t[130]) | (t[127] & ~t[128] & ~t[130]) | (t[127] & ~t[128] & ~t[129]);
  assign t[78] = (~t[131] & t[132] & t[133] & t[134]) | (t[131] & ~t[133] & ~t[134]) | (t[131] & ~t[132] & ~t[134]) | (t[131] & ~t[132] & ~t[133]);
  assign t[79] = t[135] ^ x[6];
  assign t[7] = ~(t[10] ^ t[38]);
  assign t[80] = t[136] ^ x[3];
  assign t[81] = t[137] ^ x[4];
  assign t[82] = t[138] ^ x[5];
  assign t[83] = t[139] ^ x[11];
  assign t[84] = t[140] ^ x[8];
  assign t[85] = t[141] ^ x[9];
  assign t[86] = t[142] ^ x[10];
  assign t[87] = t[143] ^ x[16];
  assign t[88] = t[144] ^ x[13];
  assign t[89] = t[145] ^ x[14];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[146] ^ x[15];
  assign t[91] = t[147] ^ x[21];
  assign t[92] = t[148] ^ x[18];
  assign t[93] = t[149] ^ x[19];
  assign t[94] = t[150] ^ x[20];
  assign t[95] = t[151] ^ x[26];
  assign t[96] = t[152] ^ x[23];
  assign t[97] = t[153] ^ x[24];
  assign t[98] = t[154] ^ x[25];
  assign t[99] = t[155] ^ x[31];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind287(x, y);
 input [71:0] x;
 output y;

 wire [190:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[156] ^ x[28];
  assign t[101] = t[157] ^ x[29];
  assign t[102] = t[158] ^ x[30];
  assign t[103] = t[159] ^ x[36];
  assign t[104] = t[160] ^ x[33];
  assign t[105] = t[161] ^ x[34];
  assign t[106] = t[162] ^ x[35];
  assign t[107] = t[163] ^ x[41];
  assign t[108] = t[164] ^ x[38];
  assign t[109] = t[165] ^ x[39];
  assign t[10] = ~t[15];
  assign t[110] = t[166] ^ x[40];
  assign t[111] = t[167] ^ x[46];
  assign t[112] = t[168] ^ x[43];
  assign t[113] = t[169] ^ x[44];
  assign t[114] = t[170] ^ x[45];
  assign t[115] = t[171] ^ x[51];
  assign t[116] = t[172] ^ x[48];
  assign t[117] = t[173] ^ x[49];
  assign t[118] = t[174] ^ x[50];
  assign t[119] = t[175] ^ x[56];
  assign t[11] = t[16] ^ t[17];
  assign t[120] = t[176] ^ x[53];
  assign t[121] = t[177] ^ x[54];
  assign t[122] = t[178] ^ x[55];
  assign t[123] = t[179] ^ x[61];
  assign t[124] = t[180] ^ x[58];
  assign t[125] = t[181] ^ x[59];
  assign t[126] = t[182] ^ x[60];
  assign t[127] = t[183] ^ x[66];
  assign t[128] = t[184] ^ x[63];
  assign t[129] = t[185] ^ x[64];
  assign t[12] = t[18] & t[19];
  assign t[130] = t[186] ^ x[65];
  assign t[131] = t[187] ^ x[71];
  assign t[132] = t[188] ^ x[68];
  assign t[133] = t[189] ^ x[69];
  assign t[134] = t[190] ^ x[70];
  assign t[135] = (x[2]);
  assign t[136] = (x[2]);
  assign t[137] = (x[2]);
  assign t[138] = (x[2]);
  assign t[139] = (x[7]);
  assign t[13] = t[20] ^ t[21];
  assign t[140] = (x[7]);
  assign t[141] = (x[7]);
  assign t[142] = (x[7]);
  assign t[143] = (x[12]);
  assign t[144] = (x[12]);
  assign t[145] = (x[12]);
  assign t[146] = (x[12]);
  assign t[147] = (x[17]);
  assign t[148] = (x[17]);
  assign t[149] = (x[17]);
  assign t[14] = t[22] & t[23];
  assign t[150] = (x[17]);
  assign t[151] = (x[22]);
  assign t[152] = (x[22]);
  assign t[153] = (x[22]);
  assign t[154] = (x[22]);
  assign t[155] = (x[27]);
  assign t[156] = (x[27]);
  assign t[157] = (x[27]);
  assign t[158] = (x[27]);
  assign t[159] = (x[32]);
  assign t[15] = ~(t[24]);
  assign t[160] = (x[32]);
  assign t[161] = (x[32]);
  assign t[162] = (x[32]);
  assign t[163] = (x[37]);
  assign t[164] = (x[37]);
  assign t[165] = (x[37]);
  assign t[166] = (x[37]);
  assign t[167] = (x[42]);
  assign t[168] = (x[42]);
  assign t[169] = (x[42]);
  assign t[16] = t[39] ^ t[40];
  assign t[170] = (x[42]);
  assign t[171] = (x[47]);
  assign t[172] = (x[47]);
  assign t[173] = (x[47]);
  assign t[174] = (x[47]);
  assign t[175] = (x[52]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[52]);
  assign t[179] = (x[57]);
  assign t[17] = t[18] & t[25];
  assign t[180] = (x[57]);
  assign t[181] = (x[57]);
  assign t[182] = (x[57]);
  assign t[183] = (x[62]);
  assign t[184] = (x[62]);
  assign t[185] = (x[62]);
  assign t[186] = (x[62]);
  assign t[187] = (x[67]);
  assign t[188] = (x[67]);
  assign t[189] = (x[67]);
  assign t[18] = ~(t[40]);
  assign t[190] = (x[67]);
  assign t[19] = ~(t[41] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[42] ^ t[43];
  assign t[21] = t[22] & t[26];
  assign t[22] = ~(t[43]);
  assign t[23] = ~(t[44] ^ t[22]);
  assign t[24] = t[27] ^ t[28];
  assign t[25] = t[41] ^ t[29];
  assign t[26] = t[44] ^ t[30];
  assign t[27] = t[31] ^ t[32];
  assign t[28] = t[33] & t[34];
  assign t[29] = t[40] ^ t[45];
  assign t[2] = ~(t[4] ^ t[37]);
  assign t[30] = t[43] ^ t[46];
  assign t[31] = t[47] ^ t[48];
  assign t[32] = t[33] & t[35];
  assign t[33] = ~(t[48]);
  assign t[34] = ~(t[49] ^ t[33]);
  assign t[35] = t[49] ^ t[36];
  assign t[36] = t[48] ^ t[50];
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = (t[57]);
  assign t[44] = (t[58]);
  assign t[45] = (t[59]);
  assign t[46] = (t[60]);
  assign t[47] = (t[61]);
  assign t[48] = (t[62]);
  assign t[49] = (t[63]);
  assign t[4] = ~t[7];
  assign t[50] = (t[64]);
  assign t[51] = t[65] ^ x[6];
  assign t[52] = t[66] ^ x[11];
  assign t[53] = t[67] ^ x[16];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[26];
  assign t[56] = t[70] ^ x[31];
  assign t[57] = t[71] ^ x[36];
  assign t[58] = t[72] ^ x[41];
  assign t[59] = t[73] ^ x[46];
  assign t[5] = ~(t[8]);
  assign t[60] = t[74] ^ x[51];
  assign t[61] = t[75] ^ x[56];
  assign t[62] = t[76] ^ x[61];
  assign t[63] = t[77] ^ x[66];
  assign t[64] = t[78] ^ x[71];
  assign t[65] = (~t[79] & t[80] & t[81] & t[82]) | (t[79] & ~t[81] & ~t[82]) | (t[79] & ~t[80] & ~t[82]) | (t[79] & ~t[80] & ~t[81]);
  assign t[66] = (~t[83] & t[84] & t[85] & t[86]) | (t[83] & ~t[85] & ~t[86]) | (t[83] & ~t[84] & ~t[86]) | (t[83] & ~t[84] & ~t[85]);
  assign t[67] = (~t[87] & t[88] & t[89] & t[90]) | (t[87] & ~t[89] & ~t[90]) | (t[87] & ~t[88] & ~t[90]) | (t[87] & ~t[88] & ~t[89]);
  assign t[68] = (~t[91] & t[92] & t[93] & t[94]) | (t[91] & ~t[93] & ~t[94]) | (t[91] & ~t[92] & ~t[94]) | (t[91] & ~t[92] & ~t[93]);
  assign t[69] = (~t[95] & t[96] & t[97] & t[98]) | (t[95] & ~t[97] & ~t[98]) | (t[95] & ~t[96] & ~t[98]) | (t[95] & ~t[96] & ~t[97]);
  assign t[6] = ~(t[9]);
  assign t[70] = (~t[99] & t[100] & t[101] & t[102]) | (t[99] & ~t[101] & ~t[102]) | (t[99] & ~t[100] & ~t[102]) | (t[99] & ~t[100] & ~t[101]);
  assign t[71] = (~t[103] & t[104] & t[105] & t[106]) | (t[103] & ~t[105] & ~t[106]) | (t[103] & ~t[104] & ~t[106]) | (t[103] & ~t[104] & ~t[105]);
  assign t[72] = (~t[107] & t[108] & t[109] & t[110]) | (t[107] & ~t[109] & ~t[110]) | (t[107] & ~t[108] & ~t[110]) | (t[107] & ~t[108] & ~t[109]);
  assign t[73] = (~t[111] & t[112] & t[113] & t[114]) | (t[111] & ~t[113] & ~t[114]) | (t[111] & ~t[112] & ~t[114]) | (t[111] & ~t[112] & ~t[113]);
  assign t[74] = (~t[115] & t[116] & t[117] & t[118]) | (t[115] & ~t[117] & ~t[118]) | (t[115] & ~t[116] & ~t[118]) | (t[115] & ~t[116] & ~t[117]);
  assign t[75] = (~t[119] & t[120] & t[121] & t[122]) | (t[119] & ~t[121] & ~t[122]) | (t[119] & ~t[120] & ~t[122]) | (t[119] & ~t[120] & ~t[121]);
  assign t[76] = (~t[123] & t[124] & t[125] & t[126]) | (t[123] & ~t[125] & ~t[126]) | (t[123] & ~t[124] & ~t[126]) | (t[123] & ~t[124] & ~t[125]);
  assign t[77] = (~t[127] & t[128] & t[129] & t[130]) | (t[127] & ~t[129] & ~t[130]) | (t[127] & ~t[128] & ~t[130]) | (t[127] & ~t[128] & ~t[129]);
  assign t[78] = (~t[131] & t[132] & t[133] & t[134]) | (t[131] & ~t[133] & ~t[134]) | (t[131] & ~t[132] & ~t[134]) | (t[131] & ~t[132] & ~t[133]);
  assign t[79] = t[135] ^ x[6];
  assign t[7] = ~(t[10] ^ t[38]);
  assign t[80] = t[136] ^ x[3];
  assign t[81] = t[137] ^ x[4];
  assign t[82] = t[138] ^ x[5];
  assign t[83] = t[139] ^ x[11];
  assign t[84] = t[140] ^ x[8];
  assign t[85] = t[141] ^ x[9];
  assign t[86] = t[142] ^ x[10];
  assign t[87] = t[143] ^ x[16];
  assign t[88] = t[144] ^ x[13];
  assign t[89] = t[145] ^ x[14];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[146] ^ x[15];
  assign t[91] = t[147] ^ x[21];
  assign t[92] = t[148] ^ x[18];
  assign t[93] = t[149] ^ x[19];
  assign t[94] = t[150] ^ x[20];
  assign t[95] = t[151] ^ x[26];
  assign t[96] = t[152] ^ x[23];
  assign t[97] = t[153] ^ x[24];
  assign t[98] = t[154] ^ x[25];
  assign t[99] = t[155] ^ x[31];
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0]);
endmodule

module R2ind288(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind289(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind290(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind291(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind292(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind293(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind294(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind295(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind296(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind297(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind298(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind299(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind300(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind301(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind302(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind303(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind304(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind305(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind306(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind307(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind308(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind309(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind310(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind311(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind312(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind313(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind314(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind315(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind316(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind317(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind318(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind319(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind320(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind321(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind322(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind323(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind324(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind325(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind326(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind327(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind328(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind329(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind330(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind331(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind332(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind333(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind334(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind335(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind336(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind337(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind338(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind339(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind340(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind341(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind342(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind343(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind344(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind345(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind346(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind347(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind348(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind349(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind350(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind351(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind352(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind353(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind354(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind355(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind356(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind357(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind358(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind359(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind360(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind361(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind362(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind363(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind364(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind365(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind366(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind367(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind368(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind369(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind370(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind371(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind372(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind373(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind374(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind375(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind376(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind377(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind378(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind379(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind380(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind381(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind382(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind383(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind384(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind385(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind386(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind387(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind388(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind389(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind390(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind391(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind392(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind393(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind394(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind395(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind396(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind397(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind398(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind399(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind400(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind401(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind402(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind403(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind404(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind405(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind406(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind407(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind408(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind409(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind410(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind411(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind412(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind413(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind414(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind415(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind416(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind417(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind418(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind419(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind420(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind421(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind422(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind423(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind424(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind425(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind426(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind427(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind428(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind429(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind430(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind431(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind432(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind433(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind434(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind435(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind436(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind437(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind438(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind439(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind440(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind441(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind442(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind443(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind444(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind445(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind446(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind447(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind448(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind449(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind450(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind451(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind452(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind453(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind454(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind455(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind456(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind457(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind458(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind459(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind460(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind461(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind462(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind463(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind464(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind465(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind466(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind467(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind468(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind469(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind470(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind471(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind472(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind473(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind474(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind475(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind476(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind477(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind478(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind479(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind480(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind481(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind482(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind483(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind484(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind485(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind486(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind487(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind488(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind489(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind490(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind491(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind492(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind493(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind494(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind495(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind496(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind497(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind498(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind499(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind500(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind501(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind502(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind503(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind504(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind505(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind506(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind507(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind508(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind509(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind510(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind511(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind512(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind513(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind514(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind515(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind516(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind517(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind518(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind519(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind520(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind521(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind522(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind523(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind524(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind525(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind526(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind527(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind528(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind529(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind530(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind531(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind532(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind533(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind534(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind535(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind536(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind537(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind538(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind539(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind540(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind541(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind542(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind543(x, y);
 input [6:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = x[0] ? x[6] : t[1];
  assign t[10] = (x[1]);
  assign t[11] = (x[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[5];
  assign t[3] = (~t[4] & t[5] & t[6] & t[7]) | (t[4] & ~t[6] & ~t[7]) | (t[4] & ~t[5] & ~t[7]) | (t[4] & ~t[5] & ~t[6]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = t[9] ^ x[2];
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = (x[1]);
  assign t[9] = (x[1]);
  assign y = (t[0]);
endmodule

module R2_ind(x, y);
 input [803:0] x;
 output [543:0] y;

  R2ind0 R2ind0_inst(.x({x[4], x[3], x[2], x[1], x[0]}), .y(y[0]));
  R2ind1 R2ind1_inst(.x({x[1], x[3], x[2], x[4], x[0]}), .y(y[1]));
  R2ind2 R2ind2_inst(.x({x[2], x[3], x[1], x[4], x[0]}), .y(y[2]));
  R2ind3 R2ind3_inst(.x({x[3], x[2], x[1], x[4], x[0]}), .y(y[3]));
  R2ind4 R2ind4_inst(.x({x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5]}), .y(y[4]));
  R2ind5 R2ind5_inst(.x({x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5]}), .y(y[5]));
  R2ind6 R2ind6_inst(.x({x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5]}), .y(y[6]));
  R2ind7 R2ind7_inst(.x({x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5]}), .y(y[7]));
  R2ind8 R2ind8_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[34], x[33], x[32], x[31], x[30], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[35]}), .y(y[8]));
  R2ind9 R2ind9_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[34], x[33], x[32], x[31], x[30], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[35]}), .y(y[9]));
  R2ind10 R2ind10_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[34], x[33], x[32], x[31], x[30], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[35]}), .y(y[10]));
  R2ind11 R2ind11_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[34], x[33], x[32], x[31], x[30], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[35]}), .y(y[11]));
  R2ind12 R2ind12_inst(.x({x[34], x[33], x[32], x[31], x[30], x[35]}), .y(y[12]));
  R2ind13 R2ind13_inst(.x({x[34], x[33], x[32], x[31], x[30], x[35]}), .y(y[13]));
  R2ind14 R2ind14_inst(.x({x[34], x[33], x[32], x[31], x[30], x[35]}), .y(y[14]));
  R2ind15 R2ind15_inst(.x({x[34], x[33], x[32], x[31], x[30], x[35]}), .y(y[15]));
  R2ind16 R2ind16_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[34], x[33], x[32], x[31], x[30], x[9], x[8], x[7], x[6], x[5], x[14], x[13], x[12], x[11], x[10], x[19], x[18], x[17], x[16], x[15], x[35]}), .y(y[16]));
  R2ind17 R2ind17_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[34], x[33], x[32], x[31], x[30], x[9], x[8], x[7], x[6], x[5], x[14], x[13], x[12], x[11], x[10], x[19], x[18], x[17], x[16], x[15], x[35]}), .y(y[17]));
  R2ind18 R2ind18_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[34], x[33], x[32], x[31], x[30], x[9], x[8], x[7], x[6], x[5], x[14], x[13], x[12], x[11], x[10], x[19], x[18], x[17], x[16], x[15], x[35]}), .y(y[18]));
  R2ind19 R2ind19_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[34], x[33], x[32], x[31], x[30], x[9], x[8], x[7], x[6], x[5], x[14], x[13], x[12], x[11], x[10], x[19], x[18], x[17], x[16], x[15], x[35]}), .y(y[19]));
  R2ind20 R2ind20_inst(.x({x[24], x[23], x[22], x[21], x[20], x[35]}), .y(y[20]));
  R2ind21 R2ind21_inst(.x({x[24], x[23], x[22], x[21], x[20], x[35]}), .y(y[21]));
  R2ind22 R2ind22_inst(.x({x[24], x[23], x[22], x[21], x[20], x[35]}), .y(y[22]));
  R2ind23 R2ind23_inst(.x({x[24], x[23], x[22], x[21], x[20], x[35]}), .y(y[23]));
  R2ind24 R2ind24_inst(.x({x[29], x[28], x[27], x[26], x[25], x[35]}), .y(y[24]));
  R2ind25 R2ind25_inst(.x({x[29], x[28], x[27], x[26], x[25], x[35]}), .y(y[25]));
  R2ind26 R2ind26_inst(.x({x[29], x[28], x[27], x[26], x[25], x[35]}), .y(y[26]));
  R2ind27 R2ind27_inst(.x({x[29], x[28], x[27], x[26], x[25], x[35]}), .y(y[27]));
  R2ind28 R2ind28_inst(.x({x[19], x[18], x[17], x[16], x[15], x[34], x[33], x[32], x[31], x[30], x[24], x[23], x[22], x[21], x[20], x[14], x[13], x[12], x[11], x[10], x[29], x[28], x[27], x[26], x[25], x[9], x[8], x[7], x[6], x[5], x[35]}), .y(y[28]));
  R2ind29 R2ind29_inst(.x({x[19], x[18], x[17], x[16], x[15], x[34], x[33], x[32], x[31], x[30], x[24], x[23], x[22], x[21], x[20], x[14], x[13], x[12], x[11], x[10], x[29], x[28], x[27], x[26], x[25], x[9], x[8], x[7], x[6], x[5], x[35]}), .y(y[29]));
  R2ind30 R2ind30_inst(.x({x[19], x[18], x[17], x[16], x[15], x[34], x[33], x[32], x[31], x[30], x[24], x[23], x[22], x[21], x[20], x[14], x[13], x[12], x[11], x[10], x[29], x[28], x[27], x[26], x[25], x[9], x[8], x[7], x[6], x[5], x[35]}), .y(y[30]));
  R2ind31 R2ind31_inst(.x({x[19], x[18], x[17], x[16], x[15], x[34], x[33], x[32], x[31], x[30], x[24], x[23], x[22], x[21], x[20], x[14], x[13], x[12], x[11], x[10], x[29], x[28], x[27], x[26], x[25], x[9], x[8], x[7], x[6], x[5], x[35]}), .y(y[31]));
  R2ind32 R2ind32_inst(.x({x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35]}), .y(y[32]));
  R2ind33 R2ind33_inst(.x({x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35]}), .y(y[33]));
  R2ind34 R2ind34_inst(.x({x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35]}), .y(y[34]));
  R2ind35 R2ind35_inst(.x({x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35]}), .y(y[35]));
  R2ind36 R2ind36_inst(.x({x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[46], x[45], x[44], x[43], x[42], x[87], x[86], x[85], x[84], x[83], x[82], x[35]}), .y(y[36]));
  R2ind37 R2ind37_inst(.x({x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[46], x[45], x[44], x[43], x[42], x[87], x[86], x[85], x[84], x[83], x[82], x[35]}), .y(y[37]));
  R2ind38 R2ind38_inst(.x({x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[46], x[45], x[44], x[43], x[42], x[87], x[86], x[85], x[84], x[83], x[82], x[35]}), .y(y[38]));
  R2ind39 R2ind39_inst(.x({x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[46], x[45], x[44], x[43], x[42], x[87], x[86], x[85], x[84], x[83], x[82], x[35]}), .y(y[39]));
  R2ind40 R2ind40_inst(.x({x[61], x[60], x[59], x[58], x[57], x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[46], x[45], x[44], x[43], x[42], x[66], x[65], x[64], x[63], x[62], x[51], x[50], x[49], x[48], x[47], x[93], x[92], x[91], x[90], x[89], x[88], x[35]}), .y(y[40]));
  R2ind41 R2ind41_inst(.x({x[61], x[60], x[59], x[58], x[57], x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[46], x[45], x[44], x[43], x[42], x[66], x[65], x[64], x[63], x[62], x[51], x[50], x[49], x[48], x[47], x[93], x[92], x[91], x[90], x[89], x[88], x[35]}), .y(y[41]));
  R2ind42 R2ind42_inst(.x({x[61], x[60], x[59], x[58], x[57], x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[46], x[45], x[44], x[43], x[42], x[66], x[65], x[64], x[63], x[62], x[51], x[50], x[49], x[48], x[47], x[93], x[92], x[91], x[90], x[89], x[88], x[35]}), .y(y[42]));
  R2ind43 R2ind43_inst(.x({x[61], x[60], x[59], x[58], x[57], x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[46], x[45], x[44], x[43], x[42], x[66], x[65], x[64], x[63], x[62], x[51], x[50], x[49], x[48], x[47], x[93], x[92], x[91], x[90], x[89], x[88], x[35]}), .y(y[43]));
  R2ind44 R2ind44_inst(.x({x[81], x[80], x[79], x[78], x[77], x[61], x[60], x[59], x[58], x[57], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[66], x[65], x[64], x[63], x[62], x[46], x[45], x[44], x[43], x[42], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[99], x[98], x[97], x[96], x[95], x[94], x[35]}), .y(y[44]));
  R2ind45 R2ind45_inst(.x({x[81], x[80], x[79], x[78], x[77], x[61], x[60], x[59], x[58], x[57], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[66], x[65], x[64], x[63], x[62], x[46], x[45], x[44], x[43], x[42], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[99], x[98], x[97], x[96], x[95], x[94], x[35]}), .y(y[45]));
  R2ind46 R2ind46_inst(.x({x[81], x[80], x[79], x[78], x[77], x[61], x[60], x[59], x[58], x[57], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[66], x[65], x[64], x[63], x[62], x[46], x[45], x[44], x[43], x[42], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[99], x[98], x[97], x[96], x[95], x[94], x[35]}), .y(y[46]));
  R2ind47 R2ind47_inst(.x({x[81], x[80], x[79], x[78], x[77], x[61], x[60], x[59], x[58], x[57], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[66], x[65], x[64], x[63], x[62], x[46], x[45], x[44], x[43], x[42], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[99], x[98], x[97], x[96], x[95], x[94], x[35]}), .y(y[47]));
  R2ind48 R2ind48_inst(.x({x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[35]}), .y(y[48]));
  R2ind49 R2ind49_inst(.x({x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[35]}), .y(y[49]));
  R2ind50 R2ind50_inst(.x({x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[35]}), .y(y[50]));
  R2ind51 R2ind51_inst(.x({x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[35]}), .y(y[51]));
  R2ind52 R2ind52_inst(.x({x[145], x[144], x[143], x[142], x[141], x[130], x[129], x[128], x[127], x[126], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[125], x[124], x[123], x[122], x[121], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[110], x[109], x[108], x[107], x[106], x[151], x[150], x[149], x[148], x[147], x[146], x[35]}), .y(y[52]));
  R2ind53 R2ind53_inst(.x({x[145], x[144], x[143], x[142], x[141], x[130], x[129], x[128], x[127], x[126], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[125], x[124], x[123], x[122], x[121], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[110], x[109], x[108], x[107], x[106], x[151], x[150], x[149], x[148], x[147], x[146], x[35]}), .y(y[53]));
  R2ind54 R2ind54_inst(.x({x[145], x[144], x[143], x[142], x[141], x[130], x[129], x[128], x[127], x[126], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[125], x[124], x[123], x[122], x[121], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[110], x[109], x[108], x[107], x[106], x[151], x[150], x[149], x[148], x[147], x[146], x[35]}), .y(y[54]));
  R2ind55 R2ind55_inst(.x({x[145], x[144], x[143], x[142], x[141], x[130], x[129], x[128], x[127], x[126], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[125], x[124], x[123], x[122], x[121], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[110], x[109], x[108], x[107], x[106], x[151], x[150], x[149], x[148], x[147], x[146], x[35]}), .y(y[55]));
  R2ind56 R2ind56_inst(.x({x[125], x[124], x[123], x[122], x[121], x[145], x[144], x[143], x[142], x[141], x[135], x[134], x[133], x[132], x[131], x[110], x[109], x[108], x[107], x[106], x[130], x[129], x[128], x[127], x[126], x[115], x[114], x[113], x[112], x[111], x[157], x[156], x[155], x[154], x[153], x[152], x[35]}), .y(y[56]));
  R2ind57 R2ind57_inst(.x({x[125], x[124], x[123], x[122], x[121], x[145], x[144], x[143], x[142], x[141], x[135], x[134], x[133], x[132], x[131], x[110], x[109], x[108], x[107], x[106], x[130], x[129], x[128], x[127], x[126], x[115], x[114], x[113], x[112], x[111], x[157], x[156], x[155], x[154], x[153], x[152], x[35]}), .y(y[57]));
  R2ind58 R2ind58_inst(.x({x[125], x[124], x[123], x[122], x[121], x[145], x[144], x[143], x[142], x[141], x[135], x[134], x[133], x[132], x[131], x[110], x[109], x[108], x[107], x[106], x[130], x[129], x[128], x[127], x[126], x[115], x[114], x[113], x[112], x[111], x[157], x[156], x[155], x[154], x[153], x[152], x[35]}), .y(y[58]));
  R2ind59 R2ind59_inst(.x({x[125], x[124], x[123], x[122], x[121], x[145], x[144], x[143], x[142], x[141], x[135], x[134], x[133], x[132], x[131], x[110], x[109], x[108], x[107], x[106], x[130], x[129], x[128], x[127], x[126], x[115], x[114], x[113], x[112], x[111], x[157], x[156], x[155], x[154], x[153], x[152], x[35]}), .y(y[59]));
  R2ind60 R2ind60_inst(.x({x[145], x[144], x[143], x[142], x[141], x[125], x[124], x[123], x[122], x[121], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[130], x[129], x[128], x[127], x[126], x[110], x[109], x[108], x[107], x[106], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[163], x[162], x[161], x[160], x[159], x[158], x[35]}), .y(y[60]));
  R2ind61 R2ind61_inst(.x({x[145], x[144], x[143], x[142], x[141], x[125], x[124], x[123], x[122], x[121], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[130], x[129], x[128], x[127], x[126], x[110], x[109], x[108], x[107], x[106], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[163], x[162], x[161], x[160], x[159], x[158], x[35]}), .y(y[61]));
  R2ind62 R2ind62_inst(.x({x[145], x[144], x[143], x[142], x[141], x[125], x[124], x[123], x[122], x[121], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[130], x[129], x[128], x[127], x[126], x[110], x[109], x[108], x[107], x[106], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[163], x[162], x[161], x[160], x[159], x[158], x[35]}), .y(y[62]));
  R2ind63 R2ind63_inst(.x({x[145], x[144], x[143], x[142], x[141], x[125], x[124], x[123], x[122], x[121], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[130], x[129], x[128], x[127], x[126], x[110], x[109], x[108], x[107], x[106], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[163], x[162], x[161], x[160], x[159], x[158], x[35]}), .y(y[63]));
  R2ind64 R2ind64_inst(.x({x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[35]}), .y(y[64]));
  R2ind65 R2ind65_inst(.x({x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[35]}), .y(y[65]));
  R2ind66 R2ind66_inst(.x({x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[35]}), .y(y[66]));
  R2ind67 R2ind67_inst(.x({x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[35]}), .y(y[67]));
  R2ind68 R2ind68_inst(.x({x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[174], x[173], x[172], x[171], x[170], x[215], x[214], x[213], x[212], x[211], x[210], x[35]}), .y(y[68]));
  R2ind69 R2ind69_inst(.x({x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[174], x[173], x[172], x[171], x[170], x[215], x[214], x[213], x[212], x[211], x[210], x[35]}), .y(y[69]));
  R2ind70 R2ind70_inst(.x({x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[174], x[173], x[172], x[171], x[170], x[215], x[214], x[213], x[212], x[211], x[210], x[35]}), .y(y[70]));
  R2ind71 R2ind71_inst(.x({x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[174], x[173], x[172], x[171], x[170], x[215], x[214], x[213], x[212], x[211], x[210], x[35]}), .y(y[71]));
  R2ind72 R2ind72_inst(.x({x[189], x[188], x[187], x[186], x[185], x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[174], x[173], x[172], x[171], x[170], x[194], x[193], x[192], x[191], x[190], x[179], x[178], x[177], x[176], x[175], x[221], x[220], x[219], x[218], x[217], x[216], x[35]}), .y(y[72]));
  R2ind73 R2ind73_inst(.x({x[189], x[188], x[187], x[186], x[185], x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[174], x[173], x[172], x[171], x[170], x[194], x[193], x[192], x[191], x[190], x[179], x[178], x[177], x[176], x[175], x[221], x[220], x[219], x[218], x[217], x[216], x[35]}), .y(y[73]));
  R2ind74 R2ind74_inst(.x({x[189], x[188], x[187], x[186], x[185], x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[174], x[173], x[172], x[171], x[170], x[194], x[193], x[192], x[191], x[190], x[179], x[178], x[177], x[176], x[175], x[221], x[220], x[219], x[218], x[217], x[216], x[35]}), .y(y[74]));
  R2ind75 R2ind75_inst(.x({x[189], x[188], x[187], x[186], x[185], x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[174], x[173], x[172], x[171], x[170], x[194], x[193], x[192], x[191], x[190], x[179], x[178], x[177], x[176], x[175], x[221], x[220], x[219], x[218], x[217], x[216], x[35]}), .y(y[75]));
  R2ind76 R2ind76_inst(.x({x[209], x[208], x[207], x[206], x[205], x[189], x[188], x[187], x[186], x[185], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[194], x[193], x[192], x[191], x[190], x[174], x[173], x[172], x[171], x[170], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[227], x[226], x[225], x[224], x[223], x[222], x[35]}), .y(y[76]));
  R2ind77 R2ind77_inst(.x({x[209], x[208], x[207], x[206], x[205], x[189], x[188], x[187], x[186], x[185], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[194], x[193], x[192], x[191], x[190], x[174], x[173], x[172], x[171], x[170], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[227], x[226], x[225], x[224], x[223], x[222], x[35]}), .y(y[77]));
  R2ind78 R2ind78_inst(.x({x[209], x[208], x[207], x[206], x[205], x[189], x[188], x[187], x[186], x[185], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[194], x[193], x[192], x[191], x[190], x[174], x[173], x[172], x[171], x[170], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[227], x[226], x[225], x[224], x[223], x[222], x[35]}), .y(y[78]));
  R2ind79 R2ind79_inst(.x({x[209], x[208], x[207], x[206], x[205], x[189], x[188], x[187], x[186], x[185], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[194], x[193], x[192], x[191], x[190], x[174], x[173], x[172], x[171], x[170], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[227], x[226], x[225], x[224], x[223], x[222], x[35]}), .y(y[79]));
  R2ind80 R2ind80_inst(.x({x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[34], x[33], x[32], x[31], x[30], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[35]}), .y(y[80]));
  R2ind81 R2ind81_inst(.x({x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[34], x[33], x[32], x[31], x[30], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[35]}), .y(y[81]));
  R2ind82 R2ind82_inst(.x({x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[34], x[33], x[32], x[31], x[30], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[35]}), .y(y[82]));
  R2ind83 R2ind83_inst(.x({x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[34], x[33], x[32], x[31], x[30], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[35]}), .y(y[83]));
  R2ind84 R2ind84_inst(.x({x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[258], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[19], x[18], x[17], x[16], x[15], x[238], x[237], x[236], x[235], x[234], x[279], x[278], x[277], x[276], x[275], x[274], x[35]}), .y(y[84]));
  R2ind85 R2ind85_inst(.x({x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[258], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[19], x[18], x[17], x[16], x[15], x[238], x[237], x[236], x[235], x[234], x[279], x[278], x[277], x[276], x[275], x[274], x[35]}), .y(y[85]));
  R2ind86 R2ind86_inst(.x({x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[258], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[19], x[18], x[17], x[16], x[15], x[238], x[237], x[236], x[235], x[234], x[279], x[278], x[277], x[276], x[275], x[274], x[35]}), .y(y[86]));
  R2ind87 R2ind87_inst(.x({x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[258], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[19], x[18], x[17], x[16], x[15], x[238], x[237], x[236], x[235], x[234], x[279], x[278], x[277], x[276], x[275], x[274], x[35]}), .y(y[87]));
  R2ind88 R2ind88_inst(.x({x[258], x[257], x[256], x[255], x[254], x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[238], x[237], x[236], x[235], x[234], x[24], x[23], x[22], x[21], x[20], x[253], x[252], x[251], x[250], x[249], x[243], x[242], x[241], x[240], x[239], x[285], x[284], x[283], x[282], x[281], x[280], x[35]}), .y(y[88]));
  R2ind89 R2ind89_inst(.x({x[258], x[257], x[256], x[255], x[254], x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[238], x[237], x[236], x[235], x[234], x[24], x[23], x[22], x[21], x[20], x[253], x[252], x[251], x[250], x[249], x[243], x[242], x[241], x[240], x[239], x[285], x[284], x[283], x[282], x[281], x[280], x[35]}), .y(y[89]));
  R2ind90 R2ind90_inst(.x({x[258], x[257], x[256], x[255], x[254], x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[238], x[237], x[236], x[235], x[234], x[24], x[23], x[22], x[21], x[20], x[253], x[252], x[251], x[250], x[249], x[243], x[242], x[241], x[240], x[239], x[285], x[284], x[283], x[282], x[281], x[280], x[35]}), .y(y[90]));
  R2ind91 R2ind91_inst(.x({x[258], x[257], x[256], x[255], x[254], x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[238], x[237], x[236], x[235], x[234], x[24], x[23], x[22], x[21], x[20], x[253], x[252], x[251], x[250], x[249], x[243], x[242], x[241], x[240], x[239], x[285], x[284], x[283], x[282], x[281], x[280], x[35]}), .y(y[91]));
  R2ind92 R2ind92_inst(.x({x[273], x[272], x[271], x[270], x[269], x[258], x[257], x[256], x[255], x[254], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[253], x[252], x[251], x[250], x[249], x[238], x[237], x[236], x[235], x[234], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[29], x[28], x[27], x[26], x[25], x[291], x[290], x[289], x[288], x[287], x[286], x[35]}), .y(y[92]));
  R2ind93 R2ind93_inst(.x({x[273], x[272], x[271], x[270], x[269], x[258], x[257], x[256], x[255], x[254], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[253], x[252], x[251], x[250], x[249], x[238], x[237], x[236], x[235], x[234], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[29], x[28], x[27], x[26], x[25], x[291], x[290], x[289], x[288], x[287], x[286], x[35]}), .y(y[93]));
  R2ind94 R2ind94_inst(.x({x[273], x[272], x[271], x[270], x[269], x[258], x[257], x[256], x[255], x[254], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[253], x[252], x[251], x[250], x[249], x[238], x[237], x[236], x[235], x[234], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[29], x[28], x[27], x[26], x[25], x[291], x[290], x[289], x[288], x[287], x[286], x[35]}), .y(y[94]));
  R2ind95 R2ind95_inst(.x({x[273], x[272], x[271], x[270], x[269], x[258], x[257], x[256], x[255], x[254], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[253], x[252], x[251], x[250], x[249], x[238], x[237], x[236], x[235], x[234], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[29], x[28], x[27], x[26], x[25], x[291], x[290], x[289], x[288], x[287], x[286], x[35]}), .y(y[95]));
  R2ind96 R2ind96_inst(.x({x[317], x[316], x[315], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[66], x[65], x[64], x[63], x[62], x[302], x[301], x[300], x[299], x[298], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[297], x[296], x[295], x[294], x[293], x[292], x[35]}), .y(y[96]));
  R2ind97 R2ind97_inst(.x({x[317], x[316], x[315], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[66], x[65], x[64], x[63], x[62], x[302], x[301], x[300], x[299], x[298], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[297], x[296], x[295], x[294], x[293], x[292], x[35]}), .y(y[97]));
  R2ind98 R2ind98_inst(.x({x[317], x[316], x[315], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[66], x[65], x[64], x[63], x[62], x[302], x[301], x[300], x[299], x[298], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[297], x[296], x[295], x[294], x[293], x[292], x[35]}), .y(y[98]));
  R2ind99 R2ind99_inst(.x({x[317], x[316], x[315], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[66], x[65], x[64], x[63], x[62], x[302], x[301], x[300], x[299], x[298], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[297], x[296], x[295], x[294], x[293], x[292], x[35]}), .y(y[99]));
  R2ind100 R2ind100_inst(.x({x[317], x[316], x[315], x[314], x[313], x[307], x[306], x[305], x[304], x[303], x[312], x[311], x[310], x[309], x[308], x[66], x[65], x[64], x[63], x[62], x[302], x[301], x[300], x[299], x[298], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[46], x[45], x[44], x[43], x[42], x[323], x[322], x[321], x[320], x[319], x[318], x[35]}), .y(y[100]));
  R2ind101 R2ind101_inst(.x({x[317], x[316], x[315], x[314], x[313], x[307], x[306], x[305], x[304], x[303], x[312], x[311], x[310], x[309], x[308], x[66], x[65], x[64], x[63], x[62], x[302], x[301], x[300], x[299], x[298], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[46], x[45], x[44], x[43], x[42], x[323], x[322], x[321], x[320], x[319], x[318], x[35]}), .y(y[101]));
  R2ind102 R2ind102_inst(.x({x[317], x[316], x[315], x[314], x[313], x[307], x[306], x[305], x[304], x[303], x[312], x[311], x[310], x[309], x[308], x[66], x[65], x[64], x[63], x[62], x[302], x[301], x[300], x[299], x[298], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[46], x[45], x[44], x[43], x[42], x[323], x[322], x[321], x[320], x[319], x[318], x[35]}), .y(y[102]));
  R2ind103 R2ind103_inst(.x({x[317], x[316], x[315], x[314], x[313], x[307], x[306], x[305], x[304], x[303], x[312], x[311], x[310], x[309], x[308], x[66], x[65], x[64], x[63], x[62], x[302], x[301], x[300], x[299], x[298], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[46], x[45], x[44], x[43], x[42], x[323], x[322], x[321], x[320], x[319], x[318], x[35]}), .y(y[103]));
  R2ind104 R2ind104_inst(.x({x[302], x[301], x[300], x[299], x[298], x[317], x[316], x[315], x[314], x[313], x[307], x[306], x[305], x[304], x[303], x[46], x[45], x[44], x[43], x[42], x[66], x[65], x[64], x[63], x[62], x[51], x[50], x[49], x[48], x[47], x[329], x[328], x[327], x[326], x[325], x[324], x[35]}), .y(y[104]));
  R2ind105 R2ind105_inst(.x({x[302], x[301], x[300], x[299], x[298], x[317], x[316], x[315], x[314], x[313], x[307], x[306], x[305], x[304], x[303], x[46], x[45], x[44], x[43], x[42], x[66], x[65], x[64], x[63], x[62], x[51], x[50], x[49], x[48], x[47], x[329], x[328], x[327], x[326], x[325], x[324], x[35]}), .y(y[105]));
  R2ind106 R2ind106_inst(.x({x[302], x[301], x[300], x[299], x[298], x[317], x[316], x[315], x[314], x[313], x[307], x[306], x[305], x[304], x[303], x[46], x[45], x[44], x[43], x[42], x[66], x[65], x[64], x[63], x[62], x[51], x[50], x[49], x[48], x[47], x[329], x[328], x[327], x[326], x[325], x[324], x[35]}), .y(y[106]));
  R2ind107 R2ind107_inst(.x({x[302], x[301], x[300], x[299], x[298], x[317], x[316], x[315], x[314], x[313], x[307], x[306], x[305], x[304], x[303], x[46], x[45], x[44], x[43], x[42], x[66], x[65], x[64], x[63], x[62], x[51], x[50], x[49], x[48], x[47], x[329], x[328], x[327], x[326], x[325], x[324], x[35]}), .y(y[107]));
  R2ind108 R2ind108_inst(.x({x[317], x[316], x[315], x[314], x[313], x[302], x[301], x[300], x[299], x[298], x[307], x[306], x[305], x[304], x[303], x[312], x[311], x[310], x[309], x[308], x[66], x[65], x[64], x[63], x[62], x[46], x[45], x[44], x[43], x[42], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[335], x[334], x[333], x[332], x[331], x[330], x[35]}), .y(y[108]));
  R2ind109 R2ind109_inst(.x({x[317], x[316], x[315], x[314], x[313], x[302], x[301], x[300], x[299], x[298], x[307], x[306], x[305], x[304], x[303], x[312], x[311], x[310], x[309], x[308], x[66], x[65], x[64], x[63], x[62], x[46], x[45], x[44], x[43], x[42], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[335], x[334], x[333], x[332], x[331], x[330], x[35]}), .y(y[109]));
  R2ind110 R2ind110_inst(.x({x[317], x[316], x[315], x[314], x[313], x[302], x[301], x[300], x[299], x[298], x[307], x[306], x[305], x[304], x[303], x[312], x[311], x[310], x[309], x[308], x[66], x[65], x[64], x[63], x[62], x[46], x[45], x[44], x[43], x[42], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[335], x[334], x[333], x[332], x[331], x[330], x[35]}), .y(y[110]));
  R2ind111 R2ind111_inst(.x({x[317], x[316], x[315], x[314], x[313], x[302], x[301], x[300], x[299], x[298], x[307], x[306], x[305], x[304], x[303], x[312], x[311], x[310], x[309], x[308], x[66], x[65], x[64], x[63], x[62], x[46], x[45], x[44], x[43], x[42], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[335], x[334], x[333], x[332], x[331], x[330], x[35]}), .y(y[111]));
  R2ind112 R2ind112_inst(.x({x[361], x[360], x[359], x[358], x[357], x[356], x[355], x[354], x[353], x[352], x[351], x[350], x[349], x[348], x[347], x[130], x[129], x[128], x[127], x[126], x[346], x[345], x[344], x[343], x[342], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[341], x[340], x[339], x[338], x[337], x[336], x[35]}), .y(y[112]));
  R2ind113 R2ind113_inst(.x({x[361], x[360], x[359], x[358], x[357], x[356], x[355], x[354], x[353], x[352], x[351], x[350], x[349], x[348], x[347], x[130], x[129], x[128], x[127], x[126], x[346], x[345], x[344], x[343], x[342], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[341], x[340], x[339], x[338], x[337], x[336], x[35]}), .y(y[113]));
  R2ind114 R2ind114_inst(.x({x[361], x[360], x[359], x[358], x[357], x[356], x[355], x[354], x[353], x[352], x[351], x[350], x[349], x[348], x[347], x[130], x[129], x[128], x[127], x[126], x[346], x[345], x[344], x[343], x[342], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[341], x[340], x[339], x[338], x[337], x[336], x[35]}), .y(y[114]));
  R2ind115 R2ind115_inst(.x({x[361], x[360], x[359], x[358], x[357], x[356], x[355], x[354], x[353], x[352], x[351], x[350], x[349], x[348], x[347], x[130], x[129], x[128], x[127], x[126], x[346], x[345], x[344], x[343], x[342], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[341], x[340], x[339], x[338], x[337], x[336], x[35]}), .y(y[115]));
  R2ind116 R2ind116_inst(.x({x[361], x[360], x[359], x[358], x[357], x[130], x[129], x[128], x[127], x[126], x[351], x[350], x[349], x[348], x[347], x[356], x[355], x[354], x[353], x[352], x[346], x[345], x[344], x[343], x[342], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[110], x[109], x[108], x[107], x[106], x[367], x[366], x[365], x[364], x[363], x[362], x[35]}), .y(y[116]));
  R2ind117 R2ind117_inst(.x({x[361], x[360], x[359], x[358], x[357], x[130], x[129], x[128], x[127], x[126], x[351], x[350], x[349], x[348], x[347], x[356], x[355], x[354], x[353], x[352], x[346], x[345], x[344], x[343], x[342], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[110], x[109], x[108], x[107], x[106], x[367], x[366], x[365], x[364], x[363], x[362], x[35]}), .y(y[117]));
  R2ind118 R2ind118_inst(.x({x[361], x[360], x[359], x[358], x[357], x[130], x[129], x[128], x[127], x[126], x[351], x[350], x[349], x[348], x[347], x[356], x[355], x[354], x[353], x[352], x[346], x[345], x[344], x[343], x[342], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[110], x[109], x[108], x[107], x[106], x[367], x[366], x[365], x[364], x[363], x[362], x[35]}), .y(y[118]));
  R2ind119 R2ind119_inst(.x({x[361], x[360], x[359], x[358], x[357], x[130], x[129], x[128], x[127], x[126], x[351], x[350], x[349], x[348], x[347], x[356], x[355], x[354], x[353], x[352], x[346], x[345], x[344], x[343], x[342], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[110], x[109], x[108], x[107], x[106], x[367], x[366], x[365], x[364], x[363], x[362], x[35]}), .y(y[119]));
  R2ind120 R2ind120_inst(.x({x[346], x[345], x[344], x[343], x[342], x[361], x[360], x[359], x[358], x[357], x[351], x[350], x[349], x[348], x[347], x[110], x[109], x[108], x[107], x[106], x[130], x[129], x[128], x[127], x[126], x[115], x[114], x[113], x[112], x[111], x[373], x[372], x[371], x[370], x[369], x[368], x[35]}), .y(y[120]));
  R2ind121 R2ind121_inst(.x({x[346], x[345], x[344], x[343], x[342], x[361], x[360], x[359], x[358], x[357], x[351], x[350], x[349], x[348], x[347], x[110], x[109], x[108], x[107], x[106], x[130], x[129], x[128], x[127], x[126], x[115], x[114], x[113], x[112], x[111], x[373], x[372], x[371], x[370], x[369], x[368], x[35]}), .y(y[121]));
  R2ind122 R2ind122_inst(.x({x[346], x[345], x[344], x[343], x[342], x[361], x[360], x[359], x[358], x[357], x[351], x[350], x[349], x[348], x[347], x[110], x[109], x[108], x[107], x[106], x[130], x[129], x[128], x[127], x[126], x[115], x[114], x[113], x[112], x[111], x[373], x[372], x[371], x[370], x[369], x[368], x[35]}), .y(y[122]));
  R2ind123 R2ind123_inst(.x({x[346], x[345], x[344], x[343], x[342], x[361], x[360], x[359], x[358], x[357], x[351], x[350], x[349], x[348], x[347], x[110], x[109], x[108], x[107], x[106], x[130], x[129], x[128], x[127], x[126], x[115], x[114], x[113], x[112], x[111], x[373], x[372], x[371], x[370], x[369], x[368], x[35]}), .y(y[123]));
  R2ind124 R2ind124_inst(.x({x[361], x[360], x[359], x[358], x[357], x[346], x[345], x[344], x[343], x[342], x[351], x[350], x[349], x[348], x[347], x[356], x[355], x[354], x[353], x[352], x[130], x[129], x[128], x[127], x[126], x[110], x[109], x[108], x[107], x[106], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[379], x[378], x[377], x[376], x[375], x[374], x[35]}), .y(y[124]));
  R2ind125 R2ind125_inst(.x({x[361], x[360], x[359], x[358], x[357], x[346], x[345], x[344], x[343], x[342], x[351], x[350], x[349], x[348], x[347], x[356], x[355], x[354], x[353], x[352], x[130], x[129], x[128], x[127], x[126], x[110], x[109], x[108], x[107], x[106], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[379], x[378], x[377], x[376], x[375], x[374], x[35]}), .y(y[125]));
  R2ind126 R2ind126_inst(.x({x[361], x[360], x[359], x[358], x[357], x[346], x[345], x[344], x[343], x[342], x[351], x[350], x[349], x[348], x[347], x[356], x[355], x[354], x[353], x[352], x[130], x[129], x[128], x[127], x[126], x[110], x[109], x[108], x[107], x[106], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[379], x[378], x[377], x[376], x[375], x[374], x[35]}), .y(y[126]));
  R2ind127 R2ind127_inst(.x({x[361], x[360], x[359], x[358], x[357], x[346], x[345], x[344], x[343], x[342], x[351], x[350], x[349], x[348], x[347], x[356], x[355], x[354], x[353], x[352], x[130], x[129], x[128], x[127], x[126], x[110], x[109], x[108], x[107], x[106], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[379], x[378], x[377], x[376], x[375], x[374], x[35]}), .y(y[127]));
  R2ind128 R2ind128_inst(.x({x[405], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[389], x[388], x[387], x[386], x[194], x[193], x[192], x[191], x[190], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[9], x[8], x[7], x[6], x[5], x[174], x[173], x[172], x[171], x[170], x[385], x[384], x[383], x[382], x[381], x[380], x[35]}), .y(y[128]));
  R2ind129 R2ind129_inst(.x({x[405], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[389], x[388], x[387], x[386], x[194], x[193], x[192], x[191], x[190], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[9], x[8], x[7], x[6], x[5], x[174], x[173], x[172], x[171], x[170], x[385], x[384], x[383], x[382], x[381], x[380], x[35]}), .y(y[129]));
  R2ind130 R2ind130_inst(.x({x[405], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[389], x[388], x[387], x[386], x[194], x[193], x[192], x[191], x[190], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[9], x[8], x[7], x[6], x[5], x[174], x[173], x[172], x[171], x[170], x[385], x[384], x[383], x[382], x[381], x[380], x[35]}), .y(y[130]));
  R2ind131 R2ind131_inst(.x({x[405], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[389], x[388], x[387], x[386], x[194], x[193], x[192], x[191], x[190], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[9], x[8], x[7], x[6], x[5], x[174], x[173], x[172], x[171], x[170], x[385], x[384], x[383], x[382], x[381], x[380], x[35]}), .y(y[131]));
  R2ind132 R2ind132_inst(.x({x[405], x[404], x[403], x[402], x[401], x[395], x[394], x[393], x[392], x[391], x[400], x[399], x[398], x[397], x[396], x[390], x[389], x[388], x[387], x[386], x[194], x[193], x[192], x[191], x[190], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[14], x[13], x[12], x[11], x[10], x[174], x[173], x[172], x[171], x[170], x[411], x[410], x[409], x[408], x[407], x[406], x[35]}), .y(y[132]));
  R2ind133 R2ind133_inst(.x({x[405], x[404], x[403], x[402], x[401], x[395], x[394], x[393], x[392], x[391], x[400], x[399], x[398], x[397], x[396], x[390], x[389], x[388], x[387], x[386], x[194], x[193], x[192], x[191], x[190], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[14], x[13], x[12], x[11], x[10], x[174], x[173], x[172], x[171], x[170], x[411], x[410], x[409], x[408], x[407], x[406], x[35]}), .y(y[133]));
  R2ind134 R2ind134_inst(.x({x[405], x[404], x[403], x[402], x[401], x[395], x[394], x[393], x[392], x[391], x[400], x[399], x[398], x[397], x[396], x[390], x[389], x[388], x[387], x[386], x[194], x[193], x[192], x[191], x[190], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[14], x[13], x[12], x[11], x[10], x[174], x[173], x[172], x[171], x[170], x[411], x[410], x[409], x[408], x[407], x[406], x[35]}), .y(y[134]));
  R2ind135 R2ind135_inst(.x({x[405], x[404], x[403], x[402], x[401], x[395], x[394], x[393], x[392], x[391], x[400], x[399], x[398], x[397], x[396], x[390], x[389], x[388], x[387], x[386], x[194], x[193], x[192], x[191], x[190], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[14], x[13], x[12], x[11], x[10], x[174], x[173], x[172], x[171], x[170], x[411], x[410], x[409], x[408], x[407], x[406], x[35]}), .y(y[135]));
  R2ind136 R2ind136_inst(.x({x[390], x[389], x[388], x[387], x[386], x[405], x[404], x[403], x[402], x[401], x[395], x[394], x[393], x[392], x[391], x[174], x[173], x[172], x[171], x[170], x[194], x[193], x[192], x[191], x[190], x[179], x[178], x[177], x[176], x[175], x[417], x[416], x[415], x[414], x[413], x[412], x[35]}), .y(y[136]));
  R2ind137 R2ind137_inst(.x({x[390], x[389], x[388], x[387], x[386], x[405], x[404], x[403], x[402], x[401], x[395], x[394], x[393], x[392], x[391], x[174], x[173], x[172], x[171], x[170], x[194], x[193], x[192], x[191], x[190], x[179], x[178], x[177], x[176], x[175], x[417], x[416], x[415], x[414], x[413], x[412], x[35]}), .y(y[137]));
  R2ind138 R2ind138_inst(.x({x[390], x[389], x[388], x[387], x[386], x[405], x[404], x[403], x[402], x[401], x[395], x[394], x[393], x[392], x[391], x[174], x[173], x[172], x[171], x[170], x[194], x[193], x[192], x[191], x[190], x[179], x[178], x[177], x[176], x[175], x[417], x[416], x[415], x[414], x[413], x[412], x[35]}), .y(y[138]));
  R2ind139 R2ind139_inst(.x({x[390], x[389], x[388], x[387], x[386], x[405], x[404], x[403], x[402], x[401], x[395], x[394], x[393], x[392], x[391], x[174], x[173], x[172], x[171], x[170], x[194], x[193], x[192], x[191], x[190], x[179], x[178], x[177], x[176], x[175], x[417], x[416], x[415], x[414], x[413], x[412], x[35]}), .y(y[139]));
  R2ind140 R2ind140_inst(.x({x[405], x[404], x[403], x[402], x[401], x[390], x[389], x[388], x[387], x[386], x[395], x[394], x[393], x[392], x[391], x[400], x[399], x[398], x[397], x[396], x[194], x[193], x[192], x[191], x[190], x[174], x[173], x[172], x[171], x[170], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[423], x[422], x[421], x[420], x[419], x[418], x[35]}), .y(y[140]));
  R2ind141 R2ind141_inst(.x({x[405], x[404], x[403], x[402], x[401], x[390], x[389], x[388], x[387], x[386], x[395], x[394], x[393], x[392], x[391], x[400], x[399], x[398], x[397], x[396], x[194], x[193], x[192], x[191], x[190], x[174], x[173], x[172], x[171], x[170], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[423], x[422], x[421], x[420], x[419], x[418], x[35]}), .y(y[141]));
  R2ind142 R2ind142_inst(.x({x[405], x[404], x[403], x[402], x[401], x[390], x[389], x[388], x[387], x[386], x[395], x[394], x[393], x[392], x[391], x[400], x[399], x[398], x[397], x[396], x[194], x[193], x[192], x[191], x[190], x[174], x[173], x[172], x[171], x[170], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[423], x[422], x[421], x[420], x[419], x[418], x[35]}), .y(y[142]));
  R2ind143 R2ind143_inst(.x({x[405], x[404], x[403], x[402], x[401], x[390], x[389], x[388], x[387], x[386], x[395], x[394], x[393], x[392], x[391], x[400], x[399], x[398], x[397], x[396], x[194], x[193], x[192], x[191], x[190], x[174], x[173], x[172], x[171], x[170], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[423], x[422], x[421], x[420], x[419], x[418], x[35]}), .y(y[143]));
  R2ind144 R2ind144_inst(.x({x[449], x[448], x[447], x[446], x[445], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[436], x[435], x[253], x[252], x[251], x[250], x[249], x[434], x[433], x[432], x[431], x[430], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[429], x[428], x[427], x[426], x[425], x[424], x[35]}), .y(y[144]));
  R2ind145 R2ind145_inst(.x({x[449], x[448], x[447], x[446], x[445], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[436], x[435], x[253], x[252], x[251], x[250], x[249], x[434], x[433], x[432], x[431], x[430], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[429], x[428], x[427], x[426], x[425], x[424], x[35]}), .y(y[145]));
  R2ind146 R2ind146_inst(.x({x[449], x[448], x[447], x[446], x[445], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[436], x[435], x[253], x[252], x[251], x[250], x[249], x[434], x[433], x[432], x[431], x[430], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[429], x[428], x[427], x[426], x[425], x[424], x[35]}), .y(y[146]));
  R2ind147 R2ind147_inst(.x({x[449], x[448], x[447], x[446], x[445], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[436], x[435], x[253], x[252], x[251], x[250], x[249], x[434], x[433], x[432], x[431], x[430], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[429], x[428], x[427], x[426], x[425], x[424], x[35]}), .y(y[147]));
  R2ind148 R2ind148_inst(.x({x[449], x[448], x[447], x[446], x[445], x[439], x[438], x[437], x[436], x[435], x[444], x[443], x[442], x[441], x[440], x[253], x[252], x[251], x[250], x[249], x[434], x[433], x[432], x[431], x[430], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[238], x[237], x[236], x[235], x[234], x[455], x[454], x[453], x[452], x[451], x[450], x[35]}), .y(y[148]));
  R2ind149 R2ind149_inst(.x({x[449], x[448], x[447], x[446], x[445], x[439], x[438], x[437], x[436], x[435], x[444], x[443], x[442], x[441], x[440], x[253], x[252], x[251], x[250], x[249], x[434], x[433], x[432], x[431], x[430], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[238], x[237], x[236], x[235], x[234], x[455], x[454], x[453], x[452], x[451], x[450], x[35]}), .y(y[149]));
  R2ind150 R2ind150_inst(.x({x[449], x[448], x[447], x[446], x[445], x[439], x[438], x[437], x[436], x[435], x[444], x[443], x[442], x[441], x[440], x[253], x[252], x[251], x[250], x[249], x[434], x[433], x[432], x[431], x[430], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[238], x[237], x[236], x[235], x[234], x[455], x[454], x[453], x[452], x[451], x[450], x[35]}), .y(y[150]));
  R2ind151 R2ind151_inst(.x({x[449], x[448], x[447], x[446], x[445], x[439], x[438], x[437], x[436], x[435], x[444], x[443], x[442], x[441], x[440], x[253], x[252], x[251], x[250], x[249], x[434], x[433], x[432], x[431], x[430], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[238], x[237], x[236], x[235], x[234], x[455], x[454], x[453], x[452], x[451], x[450], x[35]}), .y(y[151]));
  R2ind152 R2ind152_inst(.x({x[434], x[433], x[432], x[431], x[430], x[449], x[448], x[447], x[446], x[445], x[439], x[438], x[437], x[436], x[435], x[238], x[237], x[236], x[235], x[234], x[253], x[252], x[251], x[250], x[249], x[243], x[242], x[241], x[240], x[239], x[461], x[460], x[459], x[458], x[457], x[456], x[35]}), .y(y[152]));
  R2ind153 R2ind153_inst(.x({x[434], x[433], x[432], x[431], x[430], x[449], x[448], x[447], x[446], x[445], x[439], x[438], x[437], x[436], x[435], x[238], x[237], x[236], x[235], x[234], x[253], x[252], x[251], x[250], x[249], x[243], x[242], x[241], x[240], x[239], x[461], x[460], x[459], x[458], x[457], x[456], x[35]}), .y(y[153]));
  R2ind154 R2ind154_inst(.x({x[434], x[433], x[432], x[431], x[430], x[449], x[448], x[447], x[446], x[445], x[439], x[438], x[437], x[436], x[435], x[238], x[237], x[236], x[235], x[234], x[253], x[252], x[251], x[250], x[249], x[243], x[242], x[241], x[240], x[239], x[461], x[460], x[459], x[458], x[457], x[456], x[35]}), .y(y[154]));
  R2ind155 R2ind155_inst(.x({x[434], x[433], x[432], x[431], x[430], x[449], x[448], x[447], x[446], x[445], x[439], x[438], x[437], x[436], x[435], x[238], x[237], x[236], x[235], x[234], x[253], x[252], x[251], x[250], x[249], x[243], x[242], x[241], x[240], x[239], x[461], x[460], x[459], x[458], x[457], x[456], x[35]}), .y(y[155]));
  R2ind156 R2ind156_inst(.x({x[449], x[448], x[447], x[446], x[445], x[434], x[433], x[432], x[431], x[430], x[439], x[438], x[437], x[436], x[435], x[444], x[443], x[442], x[441], x[440], x[253], x[252], x[251], x[250], x[249], x[238], x[237], x[236], x[235], x[234], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[467], x[466], x[465], x[464], x[463], x[462], x[35]}), .y(y[156]));
  R2ind157 R2ind157_inst(.x({x[449], x[448], x[447], x[446], x[445], x[434], x[433], x[432], x[431], x[430], x[439], x[438], x[437], x[436], x[435], x[444], x[443], x[442], x[441], x[440], x[253], x[252], x[251], x[250], x[249], x[238], x[237], x[236], x[235], x[234], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[467], x[466], x[465], x[464], x[463], x[462], x[35]}), .y(y[157]));
  R2ind158 R2ind158_inst(.x({x[449], x[448], x[447], x[446], x[445], x[434], x[433], x[432], x[431], x[430], x[439], x[438], x[437], x[436], x[435], x[444], x[443], x[442], x[441], x[440], x[253], x[252], x[251], x[250], x[249], x[238], x[237], x[236], x[235], x[234], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[467], x[466], x[465], x[464], x[463], x[462], x[35]}), .y(y[158]));
  R2ind159 R2ind159_inst(.x({x[449], x[448], x[447], x[446], x[445], x[434], x[433], x[432], x[431], x[430], x[439], x[438], x[437], x[436], x[435], x[444], x[443], x[442], x[441], x[440], x[253], x[252], x[251], x[250], x[249], x[238], x[237], x[236], x[235], x[234], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[467], x[466], x[465], x[464], x[463], x[462], x[35]}), .y(y[159]));
  R2ind160 R2ind160_inst(.x({x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[61], x[60], x[59], x[58], x[57], x[41], x[40], x[39], x[38], x[37], x[468], x[35]}), .y(y[160]));
  R2ind161 R2ind161_inst(.x({x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[61], x[60], x[59], x[58], x[57], x[41], x[40], x[39], x[38], x[37], x[468], x[35]}), .y(y[161]));
  R2ind162 R2ind162_inst(.x({x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[61], x[60], x[59], x[58], x[57], x[41], x[40], x[39], x[38], x[37], x[468], x[35]}), .y(y[162]));
  R2ind163 R2ind163_inst(.x({x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[61], x[60], x[59], x[58], x[57], x[41], x[40], x[39], x[38], x[37], x[468], x[35]}), .y(y[163]));
  R2ind164 R2ind164_inst(.x({x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[61], x[60], x[59], x[58], x[57], x[87], x[86], x[85], x[84], x[83], x[469], x[35]}), .y(y[164]));
  R2ind165 R2ind165_inst(.x({x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[61], x[60], x[59], x[58], x[57], x[87], x[86], x[85], x[84], x[83], x[469], x[35]}), .y(y[165]));
  R2ind166 R2ind166_inst(.x({x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[61], x[60], x[59], x[58], x[57], x[87], x[86], x[85], x[84], x[83], x[469], x[35]}), .y(y[166]));
  R2ind167 R2ind167_inst(.x({x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[61], x[60], x[59], x[58], x[57], x[87], x[86], x[85], x[84], x[83], x[469], x[35]}), .y(y[167]));
  R2ind168 R2ind168_inst(.x({x[61], x[60], x[59], x[58], x[57], x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[93], x[92], x[91], x[90], x[89], x[470], x[35]}), .y(y[168]));
  R2ind169 R2ind169_inst(.x({x[61], x[60], x[59], x[58], x[57], x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[93], x[92], x[91], x[90], x[89], x[470], x[35]}), .y(y[169]));
  R2ind170 R2ind170_inst(.x({x[61], x[60], x[59], x[58], x[57], x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[93], x[92], x[91], x[90], x[89], x[470], x[35]}), .y(y[170]));
  R2ind171 R2ind171_inst(.x({x[61], x[60], x[59], x[58], x[57], x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[93], x[92], x[91], x[90], x[89], x[470], x[35]}), .y(y[171]));
  R2ind172 R2ind172_inst(.x({x[81], x[80], x[79], x[78], x[77], x[61], x[60], x[59], x[58], x[57], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[99], x[98], x[97], x[96], x[95], x[471], x[35]}), .y(y[172]));
  R2ind173 R2ind173_inst(.x({x[81], x[80], x[79], x[78], x[77], x[61], x[60], x[59], x[58], x[57], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[99], x[98], x[97], x[96], x[95], x[471], x[35]}), .y(y[173]));
  R2ind174 R2ind174_inst(.x({x[81], x[80], x[79], x[78], x[77], x[61], x[60], x[59], x[58], x[57], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[99], x[98], x[97], x[96], x[95], x[471], x[35]}), .y(y[174]));
  R2ind175 R2ind175_inst(.x({x[81], x[80], x[79], x[78], x[77], x[61], x[60], x[59], x[58], x[57], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[99], x[98], x[97], x[96], x[95], x[471], x[35]}), .y(y[175]));
  R2ind176 R2ind176_inst(.x({x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[125], x[124], x[123], x[122], x[121], x[105], x[104], x[103], x[102], x[101], x[472], x[35]}), .y(y[176]));
  R2ind177 R2ind177_inst(.x({x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[125], x[124], x[123], x[122], x[121], x[105], x[104], x[103], x[102], x[101], x[472], x[35]}), .y(y[177]));
  R2ind178 R2ind178_inst(.x({x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[125], x[124], x[123], x[122], x[121], x[105], x[104], x[103], x[102], x[101], x[472], x[35]}), .y(y[178]));
  R2ind179 R2ind179_inst(.x({x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[125], x[124], x[123], x[122], x[121], x[105], x[104], x[103], x[102], x[101], x[472], x[35]}), .y(y[179]));
  R2ind180 R2ind180_inst(.x({x[145], x[144], x[143], x[142], x[141], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[125], x[124], x[123], x[122], x[121], x[151], x[150], x[149], x[148], x[147], x[473], x[35]}), .y(y[180]));
  R2ind181 R2ind181_inst(.x({x[145], x[144], x[143], x[142], x[141], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[125], x[124], x[123], x[122], x[121], x[151], x[150], x[149], x[148], x[147], x[473], x[35]}), .y(y[181]));
  R2ind182 R2ind182_inst(.x({x[145], x[144], x[143], x[142], x[141], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[125], x[124], x[123], x[122], x[121], x[151], x[150], x[149], x[148], x[147], x[473], x[35]}), .y(y[182]));
  R2ind183 R2ind183_inst(.x({x[145], x[144], x[143], x[142], x[141], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[125], x[124], x[123], x[122], x[121], x[151], x[150], x[149], x[148], x[147], x[473], x[35]}), .y(y[183]));
  R2ind184 R2ind184_inst(.x({x[125], x[124], x[123], x[122], x[121], x[145], x[144], x[143], x[142], x[141], x[135], x[134], x[133], x[132], x[131], x[157], x[156], x[155], x[154], x[153], x[474], x[35]}), .y(y[184]));
  R2ind185 R2ind185_inst(.x({x[125], x[124], x[123], x[122], x[121], x[145], x[144], x[143], x[142], x[141], x[135], x[134], x[133], x[132], x[131], x[157], x[156], x[155], x[154], x[153], x[474], x[35]}), .y(y[185]));
  R2ind186 R2ind186_inst(.x({x[125], x[124], x[123], x[122], x[121], x[145], x[144], x[143], x[142], x[141], x[135], x[134], x[133], x[132], x[131], x[157], x[156], x[155], x[154], x[153], x[474], x[35]}), .y(y[186]));
  R2ind187 R2ind187_inst(.x({x[125], x[124], x[123], x[122], x[121], x[145], x[144], x[143], x[142], x[141], x[135], x[134], x[133], x[132], x[131], x[157], x[156], x[155], x[154], x[153], x[474], x[35]}), .y(y[187]));
  R2ind188 R2ind188_inst(.x({x[145], x[144], x[143], x[142], x[141], x[125], x[124], x[123], x[122], x[121], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[163], x[162], x[161], x[160], x[159], x[475], x[35]}), .y(y[188]));
  R2ind189 R2ind189_inst(.x({x[145], x[144], x[143], x[142], x[141], x[125], x[124], x[123], x[122], x[121], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[163], x[162], x[161], x[160], x[159], x[475], x[35]}), .y(y[189]));
  R2ind190 R2ind190_inst(.x({x[145], x[144], x[143], x[142], x[141], x[125], x[124], x[123], x[122], x[121], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[163], x[162], x[161], x[160], x[159], x[475], x[35]}), .y(y[190]));
  R2ind191 R2ind191_inst(.x({x[145], x[144], x[143], x[142], x[141], x[125], x[124], x[123], x[122], x[121], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[163], x[162], x[161], x[160], x[159], x[475], x[35]}), .y(y[191]));
  R2ind192 R2ind192_inst(.x({x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[189], x[188], x[187], x[186], x[185], x[169], x[168], x[167], x[166], x[165], x[476], x[35]}), .y(y[192]));
  R2ind193 R2ind193_inst(.x({x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[189], x[188], x[187], x[186], x[185], x[169], x[168], x[167], x[166], x[165], x[476], x[35]}), .y(y[193]));
  R2ind194 R2ind194_inst(.x({x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[189], x[188], x[187], x[186], x[185], x[169], x[168], x[167], x[166], x[165], x[476], x[35]}), .y(y[194]));
  R2ind195 R2ind195_inst(.x({x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[189], x[188], x[187], x[186], x[185], x[169], x[168], x[167], x[166], x[165], x[476], x[35]}), .y(y[195]));
  R2ind196 R2ind196_inst(.x({x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[189], x[188], x[187], x[186], x[185], x[215], x[214], x[213], x[212], x[211], x[477], x[35]}), .y(y[196]));
  R2ind197 R2ind197_inst(.x({x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[189], x[188], x[187], x[186], x[185], x[215], x[214], x[213], x[212], x[211], x[477], x[35]}), .y(y[197]));
  R2ind198 R2ind198_inst(.x({x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[189], x[188], x[187], x[186], x[185], x[215], x[214], x[213], x[212], x[211], x[477], x[35]}), .y(y[198]));
  R2ind199 R2ind199_inst(.x({x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[189], x[188], x[187], x[186], x[185], x[215], x[214], x[213], x[212], x[211], x[477], x[35]}), .y(y[199]));
  R2ind200 R2ind200_inst(.x({x[189], x[188], x[187], x[186], x[185], x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[221], x[220], x[219], x[218], x[217], x[478], x[35]}), .y(y[200]));
  R2ind201 R2ind201_inst(.x({x[189], x[188], x[187], x[186], x[185], x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[221], x[220], x[219], x[218], x[217], x[478], x[35]}), .y(y[201]));
  R2ind202 R2ind202_inst(.x({x[189], x[188], x[187], x[186], x[185], x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[221], x[220], x[219], x[218], x[217], x[478], x[35]}), .y(y[202]));
  R2ind203 R2ind203_inst(.x({x[189], x[188], x[187], x[186], x[185], x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[221], x[220], x[219], x[218], x[217], x[478], x[35]}), .y(y[203]));
  R2ind204 R2ind204_inst(.x({x[209], x[208], x[207], x[206], x[205], x[189], x[188], x[187], x[186], x[185], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[227], x[226], x[225], x[224], x[223], x[479], x[35]}), .y(y[204]));
  R2ind205 R2ind205_inst(.x({x[209], x[208], x[207], x[206], x[205], x[189], x[188], x[187], x[186], x[185], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[227], x[226], x[225], x[224], x[223], x[479], x[35]}), .y(y[205]));
  R2ind206 R2ind206_inst(.x({x[209], x[208], x[207], x[206], x[205], x[189], x[188], x[187], x[186], x[185], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[227], x[226], x[225], x[224], x[223], x[479], x[35]}), .y(y[206]));
  R2ind207 R2ind207_inst(.x({x[209], x[208], x[207], x[206], x[205], x[189], x[188], x[187], x[186], x[185], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[227], x[226], x[225], x[224], x[223], x[479], x[35]}), .y(y[207]));
  R2ind208 R2ind208_inst(.x({x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[256], x[255], x[254], x[34], x[33], x[32], x[31], x[30], x[233], x[232], x[231], x[230], x[229], x[480], x[35]}), .y(y[208]));
  R2ind209 R2ind209_inst(.x({x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[256], x[255], x[254], x[34], x[33], x[32], x[31], x[30], x[233], x[232], x[231], x[230], x[229], x[480], x[35]}), .y(y[209]));
  R2ind210 R2ind210_inst(.x({x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[256], x[255], x[254], x[34], x[33], x[32], x[31], x[30], x[233], x[232], x[231], x[230], x[229], x[480], x[35]}), .y(y[210]));
  R2ind211 R2ind211_inst(.x({x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[256], x[255], x[254], x[34], x[33], x[32], x[31], x[30], x[233], x[232], x[231], x[230], x[229], x[480], x[35]}), .y(y[211]));
  R2ind212 R2ind212_inst(.x({x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[258], x[257], x[256], x[255], x[254], x[19], x[18], x[17], x[16], x[15], x[279], x[278], x[277], x[276], x[275], x[481], x[35]}), .y(y[212]));
  R2ind213 R2ind213_inst(.x({x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[258], x[257], x[256], x[255], x[254], x[19], x[18], x[17], x[16], x[15], x[279], x[278], x[277], x[276], x[275], x[481], x[35]}), .y(y[213]));
  R2ind214 R2ind214_inst(.x({x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[258], x[257], x[256], x[255], x[254], x[19], x[18], x[17], x[16], x[15], x[279], x[278], x[277], x[276], x[275], x[481], x[35]}), .y(y[214]));
  R2ind215 R2ind215_inst(.x({x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[258], x[257], x[256], x[255], x[254], x[19], x[18], x[17], x[16], x[15], x[279], x[278], x[277], x[276], x[275], x[481], x[35]}), .y(y[215]));
  R2ind216 R2ind216_inst(.x({x[258], x[257], x[256], x[255], x[254], x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[24], x[23], x[22], x[21], x[20], x[285], x[284], x[283], x[282], x[281], x[482], x[35]}), .y(y[216]));
  R2ind217 R2ind217_inst(.x({x[258], x[257], x[256], x[255], x[254], x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[24], x[23], x[22], x[21], x[20], x[285], x[284], x[283], x[282], x[281], x[482], x[35]}), .y(y[217]));
  R2ind218 R2ind218_inst(.x({x[258], x[257], x[256], x[255], x[254], x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[24], x[23], x[22], x[21], x[20], x[285], x[284], x[283], x[282], x[281], x[482], x[35]}), .y(y[218]));
  R2ind219 R2ind219_inst(.x({x[258], x[257], x[256], x[255], x[254], x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[24], x[23], x[22], x[21], x[20], x[285], x[284], x[283], x[282], x[281], x[482], x[35]}), .y(y[219]));
  R2ind220 R2ind220_inst(.x({x[273], x[272], x[271], x[270], x[269], x[258], x[257], x[256], x[255], x[254], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[29], x[28], x[27], x[26], x[25], x[291], x[290], x[289], x[288], x[287], x[483], x[35]}), .y(y[220]));
  R2ind221 R2ind221_inst(.x({x[273], x[272], x[271], x[270], x[269], x[258], x[257], x[256], x[255], x[254], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[29], x[28], x[27], x[26], x[25], x[291], x[290], x[289], x[288], x[287], x[483], x[35]}), .y(y[221]));
  R2ind222 R2ind222_inst(.x({x[273], x[272], x[271], x[270], x[269], x[258], x[257], x[256], x[255], x[254], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[29], x[28], x[27], x[26], x[25], x[291], x[290], x[289], x[288], x[287], x[483], x[35]}), .y(y[222]));
  R2ind223 R2ind223_inst(.x({x[273], x[272], x[271], x[270], x[269], x[258], x[257], x[256], x[255], x[254], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[29], x[28], x[27], x[26], x[25], x[291], x[290], x[289], x[288], x[287], x[483], x[35]}), .y(y[223]));
  R2ind224 R2ind224_inst(.x({x[81], x[80], x[79], x[78], x[77], x[504], x[503], x[502], x[501], x[500], x[66], x[65], x[64], x[63], x[62], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[499], x[498], x[497], x[496], x[495], x[494], x[493], x[492], x[491], x[490], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[61], x[60], x[59], x[58], x[57], x[489], x[488], x[487], x[486], x[485], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[484], x[35]}), .y(y[224]));
  R2ind225 R2ind225_inst(.x({x[81], x[80], x[79], x[78], x[77], x[504], x[503], x[502], x[501], x[500], x[66], x[65], x[64], x[63], x[62], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[499], x[498], x[497], x[496], x[495], x[494], x[493], x[492], x[491], x[490], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[61], x[60], x[59], x[58], x[57], x[489], x[488], x[487], x[486], x[485], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[484], x[35]}), .y(y[225]));
  R2ind226 R2ind226_inst(.x({x[81], x[80], x[79], x[78], x[77], x[504], x[503], x[502], x[501], x[500], x[66], x[65], x[64], x[63], x[62], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[499], x[498], x[497], x[496], x[495], x[494], x[493], x[492], x[491], x[490], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[61], x[60], x[59], x[58], x[57], x[489], x[488], x[487], x[486], x[485], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[484], x[35]}), .y(y[226]));
  R2ind227 R2ind227_inst(.x({x[81], x[80], x[79], x[78], x[77], x[504], x[503], x[502], x[501], x[500], x[66], x[65], x[64], x[63], x[62], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[499], x[498], x[497], x[496], x[495], x[494], x[493], x[492], x[491], x[490], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[61], x[60], x[59], x[58], x[57], x[489], x[488], x[487], x[486], x[485], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[484], x[35]}), .y(y[227]));
  R2ind228 R2ind228_inst(.x({x[81], x[80], x[79], x[78], x[77], x[504], x[503], x[502], x[501], x[500], x[66], x[65], x[64], x[63], x[62], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[494], x[493], x[492], x[491], x[490], x[499], x[498], x[497], x[496], x[495], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[61], x[60], x[59], x[58], x[57], x[489], x[488], x[487], x[486], x[485], x[46], x[45], x[44], x[43], x[42], x[87], x[86], x[85], x[84], x[83], x[505], x[35]}), .y(y[228]));
  R2ind229 R2ind229_inst(.x({x[81], x[80], x[79], x[78], x[77], x[504], x[503], x[502], x[501], x[500], x[66], x[65], x[64], x[63], x[62], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[494], x[493], x[492], x[491], x[490], x[499], x[498], x[497], x[496], x[495], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[61], x[60], x[59], x[58], x[57], x[489], x[488], x[487], x[486], x[485], x[46], x[45], x[44], x[43], x[42], x[87], x[86], x[85], x[84], x[83], x[505], x[35]}), .y(y[229]));
  R2ind230 R2ind230_inst(.x({x[81], x[80], x[79], x[78], x[77], x[504], x[503], x[502], x[501], x[500], x[66], x[65], x[64], x[63], x[62], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[494], x[493], x[492], x[491], x[490], x[499], x[498], x[497], x[496], x[495], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[61], x[60], x[59], x[58], x[57], x[489], x[488], x[487], x[486], x[485], x[46], x[45], x[44], x[43], x[42], x[87], x[86], x[85], x[84], x[83], x[505], x[35]}), .y(y[230]));
  R2ind231 R2ind231_inst(.x({x[81], x[80], x[79], x[78], x[77], x[504], x[503], x[502], x[501], x[500], x[66], x[65], x[64], x[63], x[62], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[494], x[493], x[492], x[491], x[490], x[499], x[498], x[497], x[496], x[495], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[61], x[60], x[59], x[58], x[57], x[489], x[488], x[487], x[486], x[485], x[46], x[45], x[44], x[43], x[42], x[87], x[86], x[85], x[84], x[83], x[505], x[35]}), .y(y[231]));
  R2ind232 R2ind232_inst(.x({x[61], x[60], x[59], x[58], x[57], x[489], x[488], x[487], x[486], x[485], x[46], x[45], x[44], x[43], x[42], x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[504], x[503], x[502], x[501], x[500], x[494], x[493], x[492], x[491], x[490], x[66], x[65], x[64], x[63], x[62], x[51], x[50], x[49], x[48], x[47], x[93], x[92], x[91], x[90], x[89], x[506], x[35]}), .y(y[232]));
  R2ind233 R2ind233_inst(.x({x[61], x[60], x[59], x[58], x[57], x[489], x[488], x[487], x[486], x[485], x[46], x[45], x[44], x[43], x[42], x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[504], x[503], x[502], x[501], x[500], x[494], x[493], x[492], x[491], x[490], x[66], x[65], x[64], x[63], x[62], x[51], x[50], x[49], x[48], x[47], x[93], x[92], x[91], x[90], x[89], x[506], x[35]}), .y(y[233]));
  R2ind234 R2ind234_inst(.x({x[61], x[60], x[59], x[58], x[57], x[489], x[488], x[487], x[486], x[485], x[46], x[45], x[44], x[43], x[42], x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[504], x[503], x[502], x[501], x[500], x[494], x[493], x[492], x[491], x[490], x[66], x[65], x[64], x[63], x[62], x[51], x[50], x[49], x[48], x[47], x[93], x[92], x[91], x[90], x[89], x[506], x[35]}), .y(y[234]));
  R2ind235 R2ind235_inst(.x({x[61], x[60], x[59], x[58], x[57], x[489], x[488], x[487], x[486], x[485], x[46], x[45], x[44], x[43], x[42], x[81], x[80], x[79], x[78], x[77], x[71], x[70], x[69], x[68], x[67], x[504], x[503], x[502], x[501], x[500], x[494], x[493], x[492], x[491], x[490], x[66], x[65], x[64], x[63], x[62], x[51], x[50], x[49], x[48], x[47], x[93], x[92], x[91], x[90], x[89], x[506], x[35]}), .y(y[235]));
  R2ind236 R2ind236_inst(.x({x[81], x[80], x[79], x[78], x[77], x[504], x[503], x[502], x[501], x[500], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[489], x[488], x[487], x[486], x[485], x[494], x[493], x[492], x[491], x[490], x[499], x[498], x[497], x[496], x[495], x[46], x[45], x[44], x[43], x[42], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[99], x[98], x[97], x[96], x[95], x[507], x[35]}), .y(y[236]));
  R2ind237 R2ind237_inst(.x({x[81], x[80], x[79], x[78], x[77], x[504], x[503], x[502], x[501], x[500], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[489], x[488], x[487], x[486], x[485], x[494], x[493], x[492], x[491], x[490], x[499], x[498], x[497], x[496], x[495], x[46], x[45], x[44], x[43], x[42], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[99], x[98], x[97], x[96], x[95], x[507], x[35]}), .y(y[237]));
  R2ind238 R2ind238_inst(.x({x[81], x[80], x[79], x[78], x[77], x[504], x[503], x[502], x[501], x[500], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[489], x[488], x[487], x[486], x[485], x[494], x[493], x[492], x[491], x[490], x[499], x[498], x[497], x[496], x[495], x[46], x[45], x[44], x[43], x[42], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[99], x[98], x[97], x[96], x[95], x[507], x[35]}), .y(y[238]));
  R2ind239 R2ind239_inst(.x({x[81], x[80], x[79], x[78], x[77], x[504], x[503], x[502], x[501], x[500], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[71], x[70], x[69], x[68], x[67], x[76], x[75], x[74], x[73], x[72], x[489], x[488], x[487], x[486], x[485], x[494], x[493], x[492], x[491], x[490], x[499], x[498], x[497], x[496], x[495], x[46], x[45], x[44], x[43], x[42], x[51], x[50], x[49], x[48], x[47], x[56], x[55], x[54], x[53], x[52], x[99], x[98], x[97], x[96], x[95], x[507], x[35]}), .y(y[239]));
  R2ind240 R2ind240_inst(.x({x[145], x[144], x[143], x[142], x[141], x[528], x[527], x[526], x[525], x[524], x[130], x[129], x[128], x[127], x[126], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[514], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[125], x[124], x[123], x[122], x[121], x[513], x[512], x[511], x[510], x[509], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[508], x[35]}), .y(y[240]));
  R2ind241 R2ind241_inst(.x({x[145], x[144], x[143], x[142], x[141], x[528], x[527], x[526], x[525], x[524], x[130], x[129], x[128], x[127], x[126], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[514], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[125], x[124], x[123], x[122], x[121], x[513], x[512], x[511], x[510], x[509], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[508], x[35]}), .y(y[241]));
  R2ind242 R2ind242_inst(.x({x[145], x[144], x[143], x[142], x[141], x[528], x[527], x[526], x[525], x[524], x[130], x[129], x[128], x[127], x[126], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[514], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[125], x[124], x[123], x[122], x[121], x[513], x[512], x[511], x[510], x[509], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[508], x[35]}), .y(y[242]));
  R2ind243 R2ind243_inst(.x({x[145], x[144], x[143], x[142], x[141], x[528], x[527], x[526], x[525], x[524], x[130], x[129], x[128], x[127], x[126], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[523], x[522], x[521], x[520], x[519], x[518], x[517], x[516], x[515], x[514], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[125], x[124], x[123], x[122], x[121], x[513], x[512], x[511], x[510], x[509], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[508], x[35]}), .y(y[243]));
  R2ind244 R2ind244_inst(.x({x[130], x[129], x[128], x[127], x[126], x[145], x[144], x[143], x[142], x[141], x[528], x[527], x[526], x[525], x[524], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[518], x[517], x[516], x[515], x[514], x[523], x[522], x[521], x[520], x[519], x[110], x[109], x[108], x[107], x[106], x[125], x[124], x[123], x[122], x[121], x[513], x[512], x[511], x[510], x[509], x[151], x[150], x[149], x[148], x[147], x[529], x[35]}), .y(y[244]));
  R2ind245 R2ind245_inst(.x({x[130], x[129], x[128], x[127], x[126], x[145], x[144], x[143], x[142], x[141], x[528], x[527], x[526], x[525], x[524], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[518], x[517], x[516], x[515], x[514], x[523], x[522], x[521], x[520], x[519], x[110], x[109], x[108], x[107], x[106], x[125], x[124], x[123], x[122], x[121], x[513], x[512], x[511], x[510], x[509], x[151], x[150], x[149], x[148], x[147], x[529], x[35]}), .y(y[245]));
  R2ind246 R2ind246_inst(.x({x[130], x[129], x[128], x[127], x[126], x[145], x[144], x[143], x[142], x[141], x[528], x[527], x[526], x[525], x[524], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[518], x[517], x[516], x[515], x[514], x[523], x[522], x[521], x[520], x[519], x[110], x[109], x[108], x[107], x[106], x[125], x[124], x[123], x[122], x[121], x[513], x[512], x[511], x[510], x[509], x[151], x[150], x[149], x[148], x[147], x[529], x[35]}), .y(y[246]));
  R2ind247 R2ind247_inst(.x({x[130], x[129], x[128], x[127], x[126], x[145], x[144], x[143], x[142], x[141], x[528], x[527], x[526], x[525], x[524], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[518], x[517], x[516], x[515], x[514], x[523], x[522], x[521], x[520], x[519], x[110], x[109], x[108], x[107], x[106], x[125], x[124], x[123], x[122], x[121], x[513], x[512], x[511], x[510], x[509], x[151], x[150], x[149], x[148], x[147], x[529], x[35]}), .y(y[247]));
  R2ind248 R2ind248_inst(.x({x[125], x[124], x[123], x[122], x[121], x[513], x[512], x[511], x[510], x[509], x[110], x[109], x[108], x[107], x[106], x[145], x[144], x[143], x[142], x[141], x[135], x[134], x[133], x[132], x[131], x[528], x[527], x[526], x[525], x[524], x[518], x[517], x[516], x[515], x[514], x[130], x[129], x[128], x[127], x[126], x[115], x[114], x[113], x[112], x[111], x[157], x[156], x[155], x[154], x[153], x[530], x[35]}), .y(y[248]));
  R2ind249 R2ind249_inst(.x({x[125], x[124], x[123], x[122], x[121], x[513], x[512], x[511], x[510], x[509], x[110], x[109], x[108], x[107], x[106], x[145], x[144], x[143], x[142], x[141], x[135], x[134], x[133], x[132], x[131], x[528], x[527], x[526], x[525], x[524], x[518], x[517], x[516], x[515], x[514], x[130], x[129], x[128], x[127], x[126], x[115], x[114], x[113], x[112], x[111], x[157], x[156], x[155], x[154], x[153], x[530], x[35]}), .y(y[249]));
  R2ind250 R2ind250_inst(.x({x[125], x[124], x[123], x[122], x[121], x[513], x[512], x[511], x[510], x[509], x[110], x[109], x[108], x[107], x[106], x[145], x[144], x[143], x[142], x[141], x[135], x[134], x[133], x[132], x[131], x[528], x[527], x[526], x[525], x[524], x[518], x[517], x[516], x[515], x[514], x[130], x[129], x[128], x[127], x[126], x[115], x[114], x[113], x[112], x[111], x[157], x[156], x[155], x[154], x[153], x[530], x[35]}), .y(y[250]));
  R2ind251 R2ind251_inst(.x({x[125], x[124], x[123], x[122], x[121], x[513], x[512], x[511], x[510], x[509], x[110], x[109], x[108], x[107], x[106], x[145], x[144], x[143], x[142], x[141], x[135], x[134], x[133], x[132], x[131], x[528], x[527], x[526], x[525], x[524], x[518], x[517], x[516], x[515], x[514], x[130], x[129], x[128], x[127], x[126], x[115], x[114], x[113], x[112], x[111], x[157], x[156], x[155], x[154], x[153], x[530], x[35]}), .y(y[251]));
  R2ind252 R2ind252_inst(.x({x[145], x[144], x[143], x[142], x[141], x[528], x[527], x[526], x[525], x[524], x[130], x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[513], x[512], x[511], x[510], x[509], x[518], x[517], x[516], x[515], x[514], x[523], x[522], x[521], x[520], x[519], x[110], x[109], x[108], x[107], x[106], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[163], x[162], x[161], x[160], x[159], x[531], x[35]}), .y(y[252]));
  R2ind253 R2ind253_inst(.x({x[145], x[144], x[143], x[142], x[141], x[528], x[527], x[526], x[525], x[524], x[130], x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[513], x[512], x[511], x[510], x[509], x[518], x[517], x[516], x[515], x[514], x[523], x[522], x[521], x[520], x[519], x[110], x[109], x[108], x[107], x[106], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[163], x[162], x[161], x[160], x[159], x[531], x[35]}), .y(y[253]));
  R2ind254 R2ind254_inst(.x({x[145], x[144], x[143], x[142], x[141], x[528], x[527], x[526], x[525], x[524], x[130], x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[513], x[512], x[511], x[510], x[509], x[518], x[517], x[516], x[515], x[514], x[523], x[522], x[521], x[520], x[519], x[110], x[109], x[108], x[107], x[106], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[163], x[162], x[161], x[160], x[159], x[531], x[35]}), .y(y[254]));
  R2ind255 R2ind255_inst(.x({x[145], x[144], x[143], x[142], x[141], x[528], x[527], x[526], x[525], x[524], x[130], x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121], x[135], x[134], x[133], x[132], x[131], x[140], x[139], x[138], x[137], x[136], x[513], x[512], x[511], x[510], x[509], x[518], x[517], x[516], x[515], x[514], x[523], x[522], x[521], x[520], x[519], x[110], x[109], x[108], x[107], x[106], x[115], x[114], x[113], x[112], x[111], x[120], x[119], x[118], x[117], x[116], x[163], x[162], x[161], x[160], x[159], x[531], x[35]}), .y(y[255]));
  R2ind256 R2ind256_inst(.x({x[209], x[208], x[207], x[206], x[205], x[552], x[551], x[550], x[549], x[548], x[194], x[193], x[192], x[191], x[190], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[547], x[546], x[545], x[544], x[543], x[542], x[541], x[540], x[539], x[538], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[189], x[188], x[187], x[186], x[185], x[537], x[536], x[535], x[534], x[533], x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[532], x[35]}), .y(y[256]));
  R2ind257 R2ind257_inst(.x({x[209], x[208], x[207], x[206], x[205], x[552], x[551], x[550], x[549], x[548], x[194], x[193], x[192], x[191], x[190], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[547], x[546], x[545], x[544], x[543], x[542], x[541], x[540], x[539], x[538], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[189], x[188], x[187], x[186], x[185], x[537], x[536], x[535], x[534], x[533], x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[532], x[35]}), .y(y[257]));
  R2ind258 R2ind258_inst(.x({x[209], x[208], x[207], x[206], x[205], x[552], x[551], x[550], x[549], x[548], x[194], x[193], x[192], x[191], x[190], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[547], x[546], x[545], x[544], x[543], x[542], x[541], x[540], x[539], x[538], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[189], x[188], x[187], x[186], x[185], x[537], x[536], x[535], x[534], x[533], x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[532], x[35]}), .y(y[258]));
  R2ind259 R2ind259_inst(.x({x[209], x[208], x[207], x[206], x[205], x[552], x[551], x[550], x[549], x[548], x[194], x[193], x[192], x[191], x[190], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[547], x[546], x[545], x[544], x[543], x[542], x[541], x[540], x[539], x[538], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[189], x[188], x[187], x[186], x[185], x[537], x[536], x[535], x[534], x[533], x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[532], x[35]}), .y(y[259]));
  R2ind260 R2ind260_inst(.x({x[209], x[208], x[207], x[206], x[205], x[552], x[551], x[550], x[549], x[548], x[194], x[193], x[192], x[191], x[190], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[542], x[541], x[540], x[539], x[538], x[547], x[546], x[545], x[544], x[543], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[189], x[188], x[187], x[186], x[185], x[537], x[536], x[535], x[534], x[533], x[174], x[173], x[172], x[171], x[170], x[215], x[214], x[213], x[212], x[211], x[553], x[35]}), .y(y[260]));
  R2ind261 R2ind261_inst(.x({x[209], x[208], x[207], x[206], x[205], x[552], x[551], x[550], x[549], x[548], x[194], x[193], x[192], x[191], x[190], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[542], x[541], x[540], x[539], x[538], x[547], x[546], x[545], x[544], x[543], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[189], x[188], x[187], x[186], x[185], x[537], x[536], x[535], x[534], x[533], x[174], x[173], x[172], x[171], x[170], x[215], x[214], x[213], x[212], x[211], x[553], x[35]}), .y(y[261]));
  R2ind262 R2ind262_inst(.x({x[209], x[208], x[207], x[206], x[205], x[552], x[551], x[550], x[549], x[548], x[194], x[193], x[192], x[191], x[190], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[542], x[541], x[540], x[539], x[538], x[547], x[546], x[545], x[544], x[543], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[189], x[188], x[187], x[186], x[185], x[537], x[536], x[535], x[534], x[533], x[174], x[173], x[172], x[171], x[170], x[215], x[214], x[213], x[212], x[211], x[553], x[35]}), .y(y[262]));
  R2ind263 R2ind263_inst(.x({x[209], x[208], x[207], x[206], x[205], x[552], x[551], x[550], x[549], x[548], x[194], x[193], x[192], x[191], x[190], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[542], x[541], x[540], x[539], x[538], x[547], x[546], x[545], x[544], x[543], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[189], x[188], x[187], x[186], x[185], x[537], x[536], x[535], x[534], x[533], x[174], x[173], x[172], x[171], x[170], x[215], x[214], x[213], x[212], x[211], x[553], x[35]}), .y(y[263]));
  R2ind264 R2ind264_inst(.x({x[189], x[188], x[187], x[186], x[185], x[537], x[536], x[535], x[534], x[533], x[174], x[173], x[172], x[171], x[170], x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[552], x[551], x[550], x[549], x[548], x[542], x[541], x[540], x[539], x[538], x[194], x[193], x[192], x[191], x[190], x[179], x[178], x[177], x[176], x[175], x[221], x[220], x[219], x[218], x[217], x[554], x[35]}), .y(y[264]));
  R2ind265 R2ind265_inst(.x({x[189], x[188], x[187], x[186], x[185], x[537], x[536], x[535], x[534], x[533], x[174], x[173], x[172], x[171], x[170], x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[552], x[551], x[550], x[549], x[548], x[542], x[541], x[540], x[539], x[538], x[194], x[193], x[192], x[191], x[190], x[179], x[178], x[177], x[176], x[175], x[221], x[220], x[219], x[218], x[217], x[554], x[35]}), .y(y[265]));
  R2ind266 R2ind266_inst(.x({x[189], x[188], x[187], x[186], x[185], x[537], x[536], x[535], x[534], x[533], x[174], x[173], x[172], x[171], x[170], x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[552], x[551], x[550], x[549], x[548], x[542], x[541], x[540], x[539], x[538], x[194], x[193], x[192], x[191], x[190], x[179], x[178], x[177], x[176], x[175], x[221], x[220], x[219], x[218], x[217], x[554], x[35]}), .y(y[266]));
  R2ind267 R2ind267_inst(.x({x[189], x[188], x[187], x[186], x[185], x[537], x[536], x[535], x[534], x[533], x[174], x[173], x[172], x[171], x[170], x[209], x[208], x[207], x[206], x[205], x[199], x[198], x[197], x[196], x[195], x[552], x[551], x[550], x[549], x[548], x[542], x[541], x[540], x[539], x[538], x[194], x[193], x[192], x[191], x[190], x[179], x[178], x[177], x[176], x[175], x[221], x[220], x[219], x[218], x[217], x[554], x[35]}), .y(y[267]));
  R2ind268 R2ind268_inst(.x({x[209], x[208], x[207], x[206], x[205], x[552], x[551], x[550], x[549], x[548], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[537], x[536], x[535], x[534], x[533], x[542], x[541], x[540], x[539], x[538], x[547], x[546], x[545], x[544], x[543], x[174], x[173], x[172], x[171], x[170], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[227], x[226], x[225], x[224], x[223], x[555], x[35]}), .y(y[268]));
  R2ind269 R2ind269_inst(.x({x[209], x[208], x[207], x[206], x[205], x[552], x[551], x[550], x[549], x[548], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[537], x[536], x[535], x[534], x[533], x[542], x[541], x[540], x[539], x[538], x[547], x[546], x[545], x[544], x[543], x[174], x[173], x[172], x[171], x[170], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[227], x[226], x[225], x[224], x[223], x[555], x[35]}), .y(y[269]));
  R2ind270 R2ind270_inst(.x({x[209], x[208], x[207], x[206], x[205], x[552], x[551], x[550], x[549], x[548], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[537], x[536], x[535], x[534], x[533], x[542], x[541], x[540], x[539], x[538], x[547], x[546], x[545], x[544], x[543], x[174], x[173], x[172], x[171], x[170], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[227], x[226], x[225], x[224], x[223], x[555], x[35]}), .y(y[270]));
  R2ind271 R2ind271_inst(.x({x[209], x[208], x[207], x[206], x[205], x[552], x[551], x[550], x[549], x[548], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[199], x[198], x[197], x[196], x[195], x[204], x[203], x[202], x[201], x[200], x[537], x[536], x[535], x[534], x[533], x[542], x[541], x[540], x[539], x[538], x[547], x[546], x[545], x[544], x[543], x[174], x[173], x[172], x[171], x[170], x[179], x[178], x[177], x[176], x[175], x[184], x[183], x[182], x[181], x[180], x[227], x[226], x[225], x[224], x[223], x[555], x[35]}), .y(y[271]));
  R2ind272 R2ind272_inst(.x({x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[576], x[575], x[574], x[573], x[572], x[253], x[252], x[251], x[250], x[249], x[258], x[257], x[256], x[255], x[254], x[571], x[570], x[569], x[568], x[567], x[566], x[565], x[564], x[563], x[562], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[561], x[560], x[559], x[558], x[557], x[238], x[237], x[236], x[235], x[234], x[34], x[33], x[32], x[31], x[30], x[233], x[232], x[231], x[230], x[229], x[556], x[35]}), .y(y[272]));
  R2ind273 R2ind273_inst(.x({x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[576], x[575], x[574], x[573], x[572], x[253], x[252], x[251], x[250], x[249], x[258], x[257], x[256], x[255], x[254], x[571], x[570], x[569], x[568], x[567], x[566], x[565], x[564], x[563], x[562], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[561], x[560], x[559], x[558], x[557], x[238], x[237], x[236], x[235], x[234], x[34], x[33], x[32], x[31], x[30], x[233], x[232], x[231], x[230], x[229], x[556], x[35]}), .y(y[273]));
  R2ind274 R2ind274_inst(.x({x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[576], x[575], x[574], x[573], x[572], x[253], x[252], x[251], x[250], x[249], x[258], x[257], x[256], x[255], x[254], x[571], x[570], x[569], x[568], x[567], x[566], x[565], x[564], x[563], x[562], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[561], x[560], x[559], x[558], x[557], x[238], x[237], x[236], x[235], x[234], x[34], x[33], x[32], x[31], x[30], x[233], x[232], x[231], x[230], x[229], x[556], x[35]}), .y(y[274]));
  R2ind275 R2ind275_inst(.x({x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[576], x[575], x[574], x[573], x[572], x[253], x[252], x[251], x[250], x[249], x[258], x[257], x[256], x[255], x[254], x[571], x[570], x[569], x[568], x[567], x[566], x[565], x[564], x[563], x[562], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[561], x[560], x[559], x[558], x[557], x[238], x[237], x[236], x[235], x[234], x[34], x[33], x[32], x[31], x[30], x[233], x[232], x[231], x[230], x[229], x[556], x[35]}), .y(y[275]));
  R2ind276 R2ind276_inst(.x({x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[576], x[575], x[574], x[573], x[572], x[253], x[252], x[251], x[250], x[249], x[258], x[257], x[256], x[255], x[254], x[566], x[565], x[564], x[563], x[562], x[571], x[570], x[569], x[568], x[567], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[561], x[560], x[559], x[558], x[557], x[238], x[237], x[236], x[235], x[234], x[19], x[18], x[17], x[16], x[15], x[279], x[278], x[277], x[276], x[275], x[577], x[35]}), .y(y[276]));
  R2ind277 R2ind277_inst(.x({x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[576], x[575], x[574], x[573], x[572], x[253], x[252], x[251], x[250], x[249], x[258], x[257], x[256], x[255], x[254], x[566], x[565], x[564], x[563], x[562], x[571], x[570], x[569], x[568], x[567], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[561], x[560], x[559], x[558], x[557], x[238], x[237], x[236], x[235], x[234], x[19], x[18], x[17], x[16], x[15], x[279], x[278], x[277], x[276], x[275], x[577], x[35]}), .y(y[277]));
  R2ind278 R2ind278_inst(.x({x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[576], x[575], x[574], x[573], x[572], x[253], x[252], x[251], x[250], x[249], x[258], x[257], x[256], x[255], x[254], x[566], x[565], x[564], x[563], x[562], x[571], x[570], x[569], x[568], x[567], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[561], x[560], x[559], x[558], x[557], x[238], x[237], x[236], x[235], x[234], x[19], x[18], x[17], x[16], x[15], x[279], x[278], x[277], x[276], x[275], x[577], x[35]}), .y(y[278]));
  R2ind279 R2ind279_inst(.x({x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[576], x[575], x[574], x[573], x[572], x[253], x[252], x[251], x[250], x[249], x[258], x[257], x[256], x[255], x[254], x[566], x[565], x[564], x[563], x[562], x[571], x[570], x[569], x[568], x[567], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[561], x[560], x[559], x[558], x[557], x[238], x[237], x[236], x[235], x[234], x[19], x[18], x[17], x[16], x[15], x[279], x[278], x[277], x[276], x[275], x[577], x[35]}), .y(y[279]));
  R2ind280 R2ind280_inst(.x({x[258], x[257], x[256], x[255], x[254], x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[561], x[560], x[559], x[558], x[557], x[238], x[237], x[236], x[235], x[234], x[576], x[575], x[574], x[573], x[572], x[566], x[565], x[564], x[563], x[562], x[253], x[252], x[251], x[250], x[249], x[243], x[242], x[241], x[240], x[239], x[24], x[23], x[22], x[21], x[20], x[285], x[284], x[283], x[282], x[281], x[578], x[35]}), .y(y[280]));
  R2ind281 R2ind281_inst(.x({x[258], x[257], x[256], x[255], x[254], x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[561], x[560], x[559], x[558], x[557], x[238], x[237], x[236], x[235], x[234], x[576], x[575], x[574], x[573], x[572], x[566], x[565], x[564], x[563], x[562], x[253], x[252], x[251], x[250], x[249], x[243], x[242], x[241], x[240], x[239], x[24], x[23], x[22], x[21], x[20], x[285], x[284], x[283], x[282], x[281], x[578], x[35]}), .y(y[281]));
  R2ind282 R2ind282_inst(.x({x[258], x[257], x[256], x[255], x[254], x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[561], x[560], x[559], x[558], x[557], x[238], x[237], x[236], x[235], x[234], x[576], x[575], x[574], x[573], x[572], x[566], x[565], x[564], x[563], x[562], x[253], x[252], x[251], x[250], x[249], x[243], x[242], x[241], x[240], x[239], x[24], x[23], x[22], x[21], x[20], x[285], x[284], x[283], x[282], x[281], x[578], x[35]}), .y(y[282]));
  R2ind283 R2ind283_inst(.x({x[258], x[257], x[256], x[255], x[254], x[273], x[272], x[271], x[270], x[269], x[263], x[262], x[261], x[260], x[259], x[561], x[560], x[559], x[558], x[557], x[238], x[237], x[236], x[235], x[234], x[576], x[575], x[574], x[573], x[572], x[566], x[565], x[564], x[563], x[562], x[253], x[252], x[251], x[250], x[249], x[243], x[242], x[241], x[240], x[239], x[24], x[23], x[22], x[21], x[20], x[285], x[284], x[283], x[282], x[281], x[578], x[35]}), .y(y[283]));
  R2ind284 R2ind284_inst(.x({x[273], x[272], x[271], x[270], x[269], x[258], x[257], x[256], x[255], x[254], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[576], x[575], x[574], x[573], x[572], x[253], x[252], x[251], x[250], x[249], x[561], x[560], x[559], x[558], x[557], x[566], x[565], x[564], x[563], x[562], x[571], x[570], x[569], x[568], x[567], x[238], x[237], x[236], x[235], x[234], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[29], x[28], x[27], x[26], x[25], x[291], x[290], x[289], x[288], x[287], x[579], x[35]}), .y(y[284]));
  R2ind285 R2ind285_inst(.x({x[273], x[272], x[271], x[270], x[269], x[258], x[257], x[256], x[255], x[254], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[576], x[575], x[574], x[573], x[572], x[253], x[252], x[251], x[250], x[249], x[561], x[560], x[559], x[558], x[557], x[566], x[565], x[564], x[563], x[562], x[571], x[570], x[569], x[568], x[567], x[238], x[237], x[236], x[235], x[234], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[29], x[28], x[27], x[26], x[25], x[291], x[290], x[289], x[288], x[287], x[579], x[35]}), .y(y[285]));
  R2ind286 R2ind286_inst(.x({x[273], x[272], x[271], x[270], x[269], x[258], x[257], x[256], x[255], x[254], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[576], x[575], x[574], x[573], x[572], x[253], x[252], x[251], x[250], x[249], x[561], x[560], x[559], x[558], x[557], x[566], x[565], x[564], x[563], x[562], x[571], x[570], x[569], x[568], x[567], x[238], x[237], x[236], x[235], x[234], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[29], x[28], x[27], x[26], x[25], x[291], x[290], x[289], x[288], x[287], x[579], x[35]}), .y(y[286]));
  R2ind287 R2ind287_inst(.x({x[273], x[272], x[271], x[270], x[269], x[258], x[257], x[256], x[255], x[254], x[263], x[262], x[261], x[260], x[259], x[268], x[267], x[266], x[265], x[264], x[576], x[575], x[574], x[573], x[572], x[253], x[252], x[251], x[250], x[249], x[561], x[560], x[559], x[558], x[557], x[566], x[565], x[564], x[563], x[562], x[571], x[570], x[569], x[568], x[567], x[238], x[237], x[236], x[235], x[234], x[243], x[242], x[241], x[240], x[239], x[248], x[247], x[246], x[245], x[244], x[29], x[28], x[27], x[26], x[25], x[291], x[290], x[289], x[288], x[287], x[579], x[35]}), .y(y[287]));
  R2ind288 R2ind288_inst(.x({x[580], x[429], x[428], x[427], x[426], x[425], x[35]}), .y(y[288]));
  R2ind289 R2ind289_inst(.x({x[580], x[429], x[428], x[427], x[426], x[425], x[35]}), .y(y[289]));
  R2ind290 R2ind290_inst(.x({x[580], x[429], x[428], x[427], x[426], x[425], x[35]}), .y(y[290]));
  R2ind291 R2ind291_inst(.x({x[580], x[429], x[428], x[427], x[426], x[425], x[35]}), .y(y[291]));
  R2ind292 R2ind292_inst(.x({x[581], x[455], x[454], x[453], x[452], x[451], x[35]}), .y(y[292]));
  R2ind293 R2ind293_inst(.x({x[581], x[455], x[454], x[453], x[452], x[451], x[35]}), .y(y[293]));
  R2ind294 R2ind294_inst(.x({x[581], x[455], x[454], x[453], x[452], x[451], x[35]}), .y(y[294]));
  R2ind295 R2ind295_inst(.x({x[581], x[455], x[454], x[453], x[452], x[451], x[35]}), .y(y[295]));
  R2ind296 R2ind296_inst(.x({x[582], x[461], x[460], x[459], x[458], x[457], x[35]}), .y(y[296]));
  R2ind297 R2ind297_inst(.x({x[582], x[461], x[460], x[459], x[458], x[457], x[35]}), .y(y[297]));
  R2ind298 R2ind298_inst(.x({x[582], x[461], x[460], x[459], x[458], x[457], x[35]}), .y(y[298]));
  R2ind299 R2ind299_inst(.x({x[582], x[461], x[460], x[459], x[458], x[457], x[35]}), .y(y[299]));
  R2ind300 R2ind300_inst(.x({x[583], x[467], x[466], x[465], x[464], x[463], x[35]}), .y(y[300]));
  R2ind301 R2ind301_inst(.x({x[583], x[467], x[466], x[465], x[464], x[463], x[35]}), .y(y[301]));
  R2ind302 R2ind302_inst(.x({x[583], x[467], x[466], x[465], x[464], x[463], x[35]}), .y(y[302]));
  R2ind303 R2ind303_inst(.x({x[583], x[467], x[466], x[465], x[464], x[463], x[35]}), .y(y[303]));
  R2ind304 R2ind304_inst(.x({x[584], x[297], x[296], x[295], x[294], x[293], x[35]}), .y(y[304]));
  R2ind305 R2ind305_inst(.x({x[584], x[297], x[296], x[295], x[294], x[293], x[35]}), .y(y[305]));
  R2ind306 R2ind306_inst(.x({x[584], x[297], x[296], x[295], x[294], x[293], x[35]}), .y(y[306]));
  R2ind307 R2ind307_inst(.x({x[584], x[297], x[296], x[295], x[294], x[293], x[35]}), .y(y[307]));
  R2ind308 R2ind308_inst(.x({x[585], x[323], x[322], x[321], x[320], x[319], x[35]}), .y(y[308]));
  R2ind309 R2ind309_inst(.x({x[585], x[323], x[322], x[321], x[320], x[319], x[35]}), .y(y[309]));
  R2ind310 R2ind310_inst(.x({x[585], x[323], x[322], x[321], x[320], x[319], x[35]}), .y(y[310]));
  R2ind311 R2ind311_inst(.x({x[585], x[323], x[322], x[321], x[320], x[319], x[35]}), .y(y[311]));
  R2ind312 R2ind312_inst(.x({x[586], x[329], x[328], x[327], x[326], x[325], x[35]}), .y(y[312]));
  R2ind313 R2ind313_inst(.x({x[586], x[329], x[328], x[327], x[326], x[325], x[35]}), .y(y[313]));
  R2ind314 R2ind314_inst(.x({x[586], x[329], x[328], x[327], x[326], x[325], x[35]}), .y(y[314]));
  R2ind315 R2ind315_inst(.x({x[586], x[329], x[328], x[327], x[326], x[325], x[35]}), .y(y[315]));
  R2ind316 R2ind316_inst(.x({x[587], x[335], x[334], x[333], x[332], x[331], x[35]}), .y(y[316]));
  R2ind317 R2ind317_inst(.x({x[587], x[335], x[334], x[333], x[332], x[331], x[35]}), .y(y[317]));
  R2ind318 R2ind318_inst(.x({x[587], x[335], x[334], x[333], x[332], x[331], x[35]}), .y(y[318]));
  R2ind319 R2ind319_inst(.x({x[587], x[335], x[334], x[333], x[332], x[331], x[35]}), .y(y[319]));
  R2ind320 R2ind320_inst(.x({x[588], x[341], x[340], x[339], x[338], x[337], x[35]}), .y(y[320]));
  R2ind321 R2ind321_inst(.x({x[588], x[341], x[340], x[339], x[338], x[337], x[35]}), .y(y[321]));
  R2ind322 R2ind322_inst(.x({x[588], x[341], x[340], x[339], x[338], x[337], x[35]}), .y(y[322]));
  R2ind323 R2ind323_inst(.x({x[588], x[341], x[340], x[339], x[338], x[337], x[35]}), .y(y[323]));
  R2ind324 R2ind324_inst(.x({x[589], x[367], x[366], x[365], x[364], x[363], x[35]}), .y(y[324]));
  R2ind325 R2ind325_inst(.x({x[589], x[367], x[366], x[365], x[364], x[363], x[35]}), .y(y[325]));
  R2ind326 R2ind326_inst(.x({x[589], x[367], x[366], x[365], x[364], x[363], x[35]}), .y(y[326]));
  R2ind327 R2ind327_inst(.x({x[589], x[367], x[366], x[365], x[364], x[363], x[35]}), .y(y[327]));
  R2ind328 R2ind328_inst(.x({x[590], x[373], x[372], x[371], x[370], x[369], x[35]}), .y(y[328]));
  R2ind329 R2ind329_inst(.x({x[590], x[373], x[372], x[371], x[370], x[369], x[35]}), .y(y[329]));
  R2ind330 R2ind330_inst(.x({x[590], x[373], x[372], x[371], x[370], x[369], x[35]}), .y(y[330]));
  R2ind331 R2ind331_inst(.x({x[590], x[373], x[372], x[371], x[370], x[369], x[35]}), .y(y[331]));
  R2ind332 R2ind332_inst(.x({x[591], x[379], x[378], x[377], x[376], x[375], x[35]}), .y(y[332]));
  R2ind333 R2ind333_inst(.x({x[591], x[379], x[378], x[377], x[376], x[375], x[35]}), .y(y[333]));
  R2ind334 R2ind334_inst(.x({x[591], x[379], x[378], x[377], x[376], x[375], x[35]}), .y(y[334]));
  R2ind335 R2ind335_inst(.x({x[591], x[379], x[378], x[377], x[376], x[375], x[35]}), .y(y[335]));
  R2ind336 R2ind336_inst(.x({x[592], x[385], x[384], x[383], x[382], x[381], x[35]}), .y(y[336]));
  R2ind337 R2ind337_inst(.x({x[592], x[385], x[384], x[383], x[382], x[381], x[35]}), .y(y[337]));
  R2ind338 R2ind338_inst(.x({x[592], x[385], x[384], x[383], x[382], x[381], x[35]}), .y(y[338]));
  R2ind339 R2ind339_inst(.x({x[592], x[385], x[384], x[383], x[382], x[381], x[35]}), .y(y[339]));
  R2ind340 R2ind340_inst(.x({x[593], x[411], x[410], x[409], x[408], x[407], x[35]}), .y(y[340]));
  R2ind341 R2ind341_inst(.x({x[593], x[411], x[410], x[409], x[408], x[407], x[35]}), .y(y[341]));
  R2ind342 R2ind342_inst(.x({x[593], x[411], x[410], x[409], x[408], x[407], x[35]}), .y(y[342]));
  R2ind343 R2ind343_inst(.x({x[593], x[411], x[410], x[409], x[408], x[407], x[35]}), .y(y[343]));
  R2ind344 R2ind344_inst(.x({x[594], x[417], x[416], x[415], x[414], x[413], x[35]}), .y(y[344]));
  R2ind345 R2ind345_inst(.x({x[594], x[417], x[416], x[415], x[414], x[413], x[35]}), .y(y[345]));
  R2ind346 R2ind346_inst(.x({x[594], x[417], x[416], x[415], x[414], x[413], x[35]}), .y(y[346]));
  R2ind347 R2ind347_inst(.x({x[594], x[417], x[416], x[415], x[414], x[413], x[35]}), .y(y[347]));
  R2ind348 R2ind348_inst(.x({x[595], x[423], x[422], x[421], x[420], x[419], x[35]}), .y(y[348]));
  R2ind349 R2ind349_inst(.x({x[595], x[423], x[422], x[421], x[420], x[419], x[35]}), .y(y[349]));
  R2ind350 R2ind350_inst(.x({x[595], x[423], x[422], x[421], x[420], x[419], x[35]}), .y(y[350]));
  R2ind351 R2ind351_inst(.x({x[595], x[423], x[422], x[421], x[420], x[419], x[35]}), .y(y[351]));
  R2ind352 R2ind352_inst(.x({x[596], x[41], x[40], x[39], x[38], x[37], x[35]}), .y(y[352]));
  R2ind353 R2ind353_inst(.x({x[596], x[41], x[40], x[39], x[38], x[37], x[35]}), .y(y[353]));
  R2ind354 R2ind354_inst(.x({x[596], x[41], x[40], x[39], x[38], x[37], x[35]}), .y(y[354]));
  R2ind355 R2ind355_inst(.x({x[596], x[41], x[40], x[39], x[38], x[37], x[35]}), .y(y[355]));
  R2ind356 R2ind356_inst(.x({x[597], x[87], x[86], x[85], x[84], x[83], x[35]}), .y(y[356]));
  R2ind357 R2ind357_inst(.x({x[597], x[87], x[86], x[85], x[84], x[83], x[35]}), .y(y[357]));
  R2ind358 R2ind358_inst(.x({x[597], x[87], x[86], x[85], x[84], x[83], x[35]}), .y(y[358]));
  R2ind359 R2ind359_inst(.x({x[597], x[87], x[86], x[85], x[84], x[83], x[35]}), .y(y[359]));
  R2ind360 R2ind360_inst(.x({x[598], x[93], x[92], x[91], x[90], x[89], x[35]}), .y(y[360]));
  R2ind361 R2ind361_inst(.x({x[598], x[93], x[92], x[91], x[90], x[89], x[35]}), .y(y[361]));
  R2ind362 R2ind362_inst(.x({x[598], x[93], x[92], x[91], x[90], x[89], x[35]}), .y(y[362]));
  R2ind363 R2ind363_inst(.x({x[598], x[93], x[92], x[91], x[90], x[89], x[35]}), .y(y[363]));
  R2ind364 R2ind364_inst(.x({x[599], x[99], x[98], x[97], x[96], x[95], x[35]}), .y(y[364]));
  R2ind365 R2ind365_inst(.x({x[599], x[99], x[98], x[97], x[96], x[95], x[35]}), .y(y[365]));
  R2ind366 R2ind366_inst(.x({x[599], x[99], x[98], x[97], x[96], x[95], x[35]}), .y(y[366]));
  R2ind367 R2ind367_inst(.x({x[599], x[99], x[98], x[97], x[96], x[95], x[35]}), .y(y[367]));
  R2ind368 R2ind368_inst(.x({x[600], x[105], x[104], x[103], x[102], x[101], x[35]}), .y(y[368]));
  R2ind369 R2ind369_inst(.x({x[600], x[105], x[104], x[103], x[102], x[101], x[35]}), .y(y[369]));
  R2ind370 R2ind370_inst(.x({x[600], x[105], x[104], x[103], x[102], x[101], x[35]}), .y(y[370]));
  R2ind371 R2ind371_inst(.x({x[600], x[105], x[104], x[103], x[102], x[101], x[35]}), .y(y[371]));
  R2ind372 R2ind372_inst(.x({x[601], x[151], x[150], x[149], x[148], x[147], x[35]}), .y(y[372]));
  R2ind373 R2ind373_inst(.x({x[601], x[151], x[150], x[149], x[148], x[147], x[35]}), .y(y[373]));
  R2ind374 R2ind374_inst(.x({x[601], x[151], x[150], x[149], x[148], x[147], x[35]}), .y(y[374]));
  R2ind375 R2ind375_inst(.x({x[601], x[151], x[150], x[149], x[148], x[147], x[35]}), .y(y[375]));
  R2ind376 R2ind376_inst(.x({x[602], x[157], x[156], x[155], x[154], x[153], x[35]}), .y(y[376]));
  R2ind377 R2ind377_inst(.x({x[602], x[157], x[156], x[155], x[154], x[153], x[35]}), .y(y[377]));
  R2ind378 R2ind378_inst(.x({x[602], x[157], x[156], x[155], x[154], x[153], x[35]}), .y(y[378]));
  R2ind379 R2ind379_inst(.x({x[602], x[157], x[156], x[155], x[154], x[153], x[35]}), .y(y[379]));
  R2ind380 R2ind380_inst(.x({x[603], x[163], x[162], x[161], x[160], x[159], x[35]}), .y(y[380]));
  R2ind381 R2ind381_inst(.x({x[603], x[163], x[162], x[161], x[160], x[159], x[35]}), .y(y[381]));
  R2ind382 R2ind382_inst(.x({x[603], x[163], x[162], x[161], x[160], x[159], x[35]}), .y(y[382]));
  R2ind383 R2ind383_inst(.x({x[603], x[163], x[162], x[161], x[160], x[159], x[35]}), .y(y[383]));
  R2ind384 R2ind384_inst(.x({x[604], x[169], x[168], x[167], x[166], x[165], x[35]}), .y(y[384]));
  R2ind385 R2ind385_inst(.x({x[604], x[169], x[168], x[167], x[166], x[165], x[35]}), .y(y[385]));
  R2ind386 R2ind386_inst(.x({x[604], x[169], x[168], x[167], x[166], x[165], x[35]}), .y(y[386]));
  R2ind387 R2ind387_inst(.x({x[604], x[169], x[168], x[167], x[166], x[165], x[35]}), .y(y[387]));
  R2ind388 R2ind388_inst(.x({x[605], x[215], x[214], x[213], x[212], x[211], x[35]}), .y(y[388]));
  R2ind389 R2ind389_inst(.x({x[605], x[215], x[214], x[213], x[212], x[211], x[35]}), .y(y[389]));
  R2ind390 R2ind390_inst(.x({x[605], x[215], x[214], x[213], x[212], x[211], x[35]}), .y(y[390]));
  R2ind391 R2ind391_inst(.x({x[605], x[215], x[214], x[213], x[212], x[211], x[35]}), .y(y[391]));
  R2ind392 R2ind392_inst(.x({x[606], x[221], x[220], x[219], x[218], x[217], x[35]}), .y(y[392]));
  R2ind393 R2ind393_inst(.x({x[606], x[221], x[220], x[219], x[218], x[217], x[35]}), .y(y[393]));
  R2ind394 R2ind394_inst(.x({x[606], x[221], x[220], x[219], x[218], x[217], x[35]}), .y(y[394]));
  R2ind395 R2ind395_inst(.x({x[606], x[221], x[220], x[219], x[218], x[217], x[35]}), .y(y[395]));
  R2ind396 R2ind396_inst(.x({x[607], x[227], x[226], x[225], x[224], x[223], x[35]}), .y(y[396]));
  R2ind397 R2ind397_inst(.x({x[607], x[227], x[226], x[225], x[224], x[223], x[35]}), .y(y[397]));
  R2ind398 R2ind398_inst(.x({x[607], x[227], x[226], x[225], x[224], x[223], x[35]}), .y(y[398]));
  R2ind399 R2ind399_inst(.x({x[607], x[227], x[226], x[225], x[224], x[223], x[35]}), .y(y[399]));
  R2ind400 R2ind400_inst(.x({x[608], x[233], x[232], x[231], x[230], x[229], x[35]}), .y(y[400]));
  R2ind401 R2ind401_inst(.x({x[608], x[233], x[232], x[231], x[230], x[229], x[35]}), .y(y[401]));
  R2ind402 R2ind402_inst(.x({x[608], x[233], x[232], x[231], x[230], x[229], x[35]}), .y(y[402]));
  R2ind403 R2ind403_inst(.x({x[608], x[233], x[232], x[231], x[230], x[229], x[35]}), .y(y[403]));
  R2ind404 R2ind404_inst(.x({x[609], x[279], x[278], x[277], x[276], x[275], x[35]}), .y(y[404]));
  R2ind405 R2ind405_inst(.x({x[609], x[279], x[278], x[277], x[276], x[275], x[35]}), .y(y[405]));
  R2ind406 R2ind406_inst(.x({x[609], x[279], x[278], x[277], x[276], x[275], x[35]}), .y(y[406]));
  R2ind407 R2ind407_inst(.x({x[609], x[279], x[278], x[277], x[276], x[275], x[35]}), .y(y[407]));
  R2ind408 R2ind408_inst(.x({x[610], x[285], x[284], x[283], x[282], x[281], x[35]}), .y(y[408]));
  R2ind409 R2ind409_inst(.x({x[610], x[285], x[284], x[283], x[282], x[281], x[35]}), .y(y[409]));
  R2ind410 R2ind410_inst(.x({x[610], x[285], x[284], x[283], x[282], x[281], x[35]}), .y(y[410]));
  R2ind411 R2ind411_inst(.x({x[610], x[285], x[284], x[283], x[282], x[281], x[35]}), .y(y[411]));
  R2ind412 R2ind412_inst(.x({x[611], x[291], x[290], x[289], x[288], x[287], x[35]}), .y(y[412]));
  R2ind413 R2ind413_inst(.x({x[611], x[291], x[290], x[289], x[288], x[287], x[35]}), .y(y[413]));
  R2ind414 R2ind414_inst(.x({x[611], x[291], x[290], x[289], x[288], x[287], x[35]}), .y(y[414]));
  R2ind415 R2ind415_inst(.x({x[611], x[291], x[290], x[289], x[288], x[287], x[35]}), .y(y[415]));
  R2ind416 R2ind416_inst(.x({x[617], x[616], x[615], x[614], x[613], x[612], x[35]}), .y(y[416]));
  R2ind417 R2ind417_inst(.x({x[617], x[616], x[615], x[614], x[613], x[612], x[35]}), .y(y[417]));
  R2ind418 R2ind418_inst(.x({x[617], x[616], x[615], x[614], x[613], x[612], x[35]}), .y(y[418]));
  R2ind419 R2ind419_inst(.x({x[617], x[616], x[615], x[614], x[613], x[612], x[35]}), .y(y[419]));
  R2ind420 R2ind420_inst(.x({x[623], x[622], x[621], x[620], x[619], x[618], x[35]}), .y(y[420]));
  R2ind421 R2ind421_inst(.x({x[623], x[622], x[621], x[620], x[619], x[618], x[35]}), .y(y[421]));
  R2ind422 R2ind422_inst(.x({x[623], x[622], x[621], x[620], x[619], x[618], x[35]}), .y(y[422]));
  R2ind423 R2ind423_inst(.x({x[623], x[622], x[621], x[620], x[619], x[618], x[35]}), .y(y[423]));
  R2ind424 R2ind424_inst(.x({x[629], x[628], x[627], x[626], x[625], x[624], x[35]}), .y(y[424]));
  R2ind425 R2ind425_inst(.x({x[629], x[628], x[627], x[626], x[625], x[624], x[35]}), .y(y[425]));
  R2ind426 R2ind426_inst(.x({x[629], x[628], x[627], x[626], x[625], x[624], x[35]}), .y(y[426]));
  R2ind427 R2ind427_inst(.x({x[629], x[628], x[627], x[626], x[625], x[624], x[35]}), .y(y[427]));
  R2ind428 R2ind428_inst(.x({x[635], x[634], x[633], x[632], x[631], x[630], x[35]}), .y(y[428]));
  R2ind429 R2ind429_inst(.x({x[635], x[634], x[633], x[632], x[631], x[630], x[35]}), .y(y[429]));
  R2ind430 R2ind430_inst(.x({x[635], x[634], x[633], x[632], x[631], x[630], x[35]}), .y(y[430]));
  R2ind431 R2ind431_inst(.x({x[635], x[634], x[633], x[632], x[631], x[630], x[35]}), .y(y[431]));
  R2ind432 R2ind432_inst(.x({x[641], x[640], x[639], x[638], x[637], x[636], x[35]}), .y(y[432]));
  R2ind433 R2ind433_inst(.x({x[641], x[640], x[639], x[638], x[637], x[636], x[35]}), .y(y[433]));
  R2ind434 R2ind434_inst(.x({x[641], x[640], x[639], x[638], x[637], x[636], x[35]}), .y(y[434]));
  R2ind435 R2ind435_inst(.x({x[641], x[640], x[639], x[638], x[637], x[636], x[35]}), .y(y[435]));
  R2ind436 R2ind436_inst(.x({x[647], x[646], x[645], x[644], x[643], x[642], x[35]}), .y(y[436]));
  R2ind437 R2ind437_inst(.x({x[647], x[646], x[645], x[644], x[643], x[642], x[35]}), .y(y[437]));
  R2ind438 R2ind438_inst(.x({x[647], x[646], x[645], x[644], x[643], x[642], x[35]}), .y(y[438]));
  R2ind439 R2ind439_inst(.x({x[647], x[646], x[645], x[644], x[643], x[642], x[35]}), .y(y[439]));
  R2ind440 R2ind440_inst(.x({x[653], x[652], x[651], x[650], x[649], x[648], x[35]}), .y(y[440]));
  R2ind441 R2ind441_inst(.x({x[653], x[652], x[651], x[650], x[649], x[648], x[35]}), .y(y[441]));
  R2ind442 R2ind442_inst(.x({x[653], x[652], x[651], x[650], x[649], x[648], x[35]}), .y(y[442]));
  R2ind443 R2ind443_inst(.x({x[653], x[652], x[651], x[650], x[649], x[648], x[35]}), .y(y[443]));
  R2ind444 R2ind444_inst(.x({x[659], x[658], x[657], x[656], x[655], x[654], x[35]}), .y(y[444]));
  R2ind445 R2ind445_inst(.x({x[659], x[658], x[657], x[656], x[655], x[654], x[35]}), .y(y[445]));
  R2ind446 R2ind446_inst(.x({x[659], x[658], x[657], x[656], x[655], x[654], x[35]}), .y(y[446]));
  R2ind447 R2ind447_inst(.x({x[659], x[658], x[657], x[656], x[655], x[654], x[35]}), .y(y[447]));
  R2ind448 R2ind448_inst(.x({x[665], x[664], x[663], x[662], x[661], x[660], x[35]}), .y(y[448]));
  R2ind449 R2ind449_inst(.x({x[665], x[664], x[663], x[662], x[661], x[660], x[35]}), .y(y[449]));
  R2ind450 R2ind450_inst(.x({x[665], x[664], x[663], x[662], x[661], x[660], x[35]}), .y(y[450]));
  R2ind451 R2ind451_inst(.x({x[665], x[664], x[663], x[662], x[661], x[660], x[35]}), .y(y[451]));
  R2ind452 R2ind452_inst(.x({x[671], x[670], x[669], x[668], x[667], x[666], x[35]}), .y(y[452]));
  R2ind453 R2ind453_inst(.x({x[671], x[670], x[669], x[668], x[667], x[666], x[35]}), .y(y[453]));
  R2ind454 R2ind454_inst(.x({x[671], x[670], x[669], x[668], x[667], x[666], x[35]}), .y(y[454]));
  R2ind455 R2ind455_inst(.x({x[671], x[670], x[669], x[668], x[667], x[666], x[35]}), .y(y[455]));
  R2ind456 R2ind456_inst(.x({x[677], x[676], x[675], x[674], x[673], x[672], x[35]}), .y(y[456]));
  R2ind457 R2ind457_inst(.x({x[677], x[676], x[675], x[674], x[673], x[672], x[35]}), .y(y[457]));
  R2ind458 R2ind458_inst(.x({x[677], x[676], x[675], x[674], x[673], x[672], x[35]}), .y(y[458]));
  R2ind459 R2ind459_inst(.x({x[677], x[676], x[675], x[674], x[673], x[672], x[35]}), .y(y[459]));
  R2ind460 R2ind460_inst(.x({x[683], x[682], x[681], x[680], x[679], x[678], x[35]}), .y(y[460]));
  R2ind461 R2ind461_inst(.x({x[683], x[682], x[681], x[680], x[679], x[678], x[35]}), .y(y[461]));
  R2ind462 R2ind462_inst(.x({x[683], x[682], x[681], x[680], x[679], x[678], x[35]}), .y(y[462]));
  R2ind463 R2ind463_inst(.x({x[683], x[682], x[681], x[680], x[679], x[678], x[35]}), .y(y[463]));
  R2ind464 R2ind464_inst(.x({x[689], x[688], x[687], x[686], x[685], x[684], x[35]}), .y(y[464]));
  R2ind465 R2ind465_inst(.x({x[689], x[688], x[687], x[686], x[685], x[684], x[35]}), .y(y[465]));
  R2ind466 R2ind466_inst(.x({x[689], x[688], x[687], x[686], x[685], x[684], x[35]}), .y(y[466]));
  R2ind467 R2ind467_inst(.x({x[689], x[688], x[687], x[686], x[685], x[684], x[35]}), .y(y[467]));
  R2ind468 R2ind468_inst(.x({x[695], x[694], x[693], x[692], x[691], x[690], x[35]}), .y(y[468]));
  R2ind469 R2ind469_inst(.x({x[695], x[694], x[693], x[692], x[691], x[690], x[35]}), .y(y[469]));
  R2ind470 R2ind470_inst(.x({x[695], x[694], x[693], x[692], x[691], x[690], x[35]}), .y(y[470]));
  R2ind471 R2ind471_inst(.x({x[695], x[694], x[693], x[692], x[691], x[690], x[35]}), .y(y[471]));
  R2ind472 R2ind472_inst(.x({x[701], x[700], x[699], x[698], x[697], x[696], x[35]}), .y(y[472]));
  R2ind473 R2ind473_inst(.x({x[701], x[700], x[699], x[698], x[697], x[696], x[35]}), .y(y[473]));
  R2ind474 R2ind474_inst(.x({x[701], x[700], x[699], x[698], x[697], x[696], x[35]}), .y(y[474]));
  R2ind475 R2ind475_inst(.x({x[701], x[700], x[699], x[698], x[697], x[696], x[35]}), .y(y[475]));
  R2ind476 R2ind476_inst(.x({x[707], x[706], x[705], x[704], x[703], x[702], x[35]}), .y(y[476]));
  R2ind477 R2ind477_inst(.x({x[707], x[706], x[705], x[704], x[703], x[702], x[35]}), .y(y[477]));
  R2ind478 R2ind478_inst(.x({x[707], x[706], x[705], x[704], x[703], x[702], x[35]}), .y(y[478]));
  R2ind479 R2ind479_inst(.x({x[707], x[706], x[705], x[704], x[703], x[702], x[35]}), .y(y[479]));
  R2ind480 R2ind480_inst(.x({x[713], x[712], x[711], x[710], x[709], x[708], x[35]}), .y(y[480]));
  R2ind481 R2ind481_inst(.x({x[713], x[712], x[711], x[710], x[709], x[708], x[35]}), .y(y[481]));
  R2ind482 R2ind482_inst(.x({x[713], x[712], x[711], x[710], x[709], x[708], x[35]}), .y(y[482]));
  R2ind483 R2ind483_inst(.x({x[713], x[712], x[711], x[710], x[709], x[708], x[35]}), .y(y[483]));
  R2ind484 R2ind484_inst(.x({x[719], x[718], x[717], x[716], x[715], x[714], x[35]}), .y(y[484]));
  R2ind485 R2ind485_inst(.x({x[719], x[718], x[717], x[716], x[715], x[714], x[35]}), .y(y[485]));
  R2ind486 R2ind486_inst(.x({x[719], x[718], x[717], x[716], x[715], x[714], x[35]}), .y(y[486]));
  R2ind487 R2ind487_inst(.x({x[719], x[718], x[717], x[716], x[715], x[714], x[35]}), .y(y[487]));
  R2ind488 R2ind488_inst(.x({x[725], x[724], x[723], x[722], x[721], x[720], x[35]}), .y(y[488]));
  R2ind489 R2ind489_inst(.x({x[725], x[724], x[723], x[722], x[721], x[720], x[35]}), .y(y[489]));
  R2ind490 R2ind490_inst(.x({x[725], x[724], x[723], x[722], x[721], x[720], x[35]}), .y(y[490]));
  R2ind491 R2ind491_inst(.x({x[725], x[724], x[723], x[722], x[721], x[720], x[35]}), .y(y[491]));
  R2ind492 R2ind492_inst(.x({x[731], x[730], x[729], x[728], x[727], x[726], x[35]}), .y(y[492]));
  R2ind493 R2ind493_inst(.x({x[731], x[730], x[729], x[728], x[727], x[726], x[35]}), .y(y[493]));
  R2ind494 R2ind494_inst(.x({x[731], x[730], x[729], x[728], x[727], x[726], x[35]}), .y(y[494]));
  R2ind495 R2ind495_inst(.x({x[731], x[730], x[729], x[728], x[727], x[726], x[35]}), .y(y[495]));
  R2ind496 R2ind496_inst(.x({x[737], x[736], x[735], x[734], x[733], x[732], x[35]}), .y(y[496]));
  R2ind497 R2ind497_inst(.x({x[737], x[736], x[735], x[734], x[733], x[732], x[35]}), .y(y[497]));
  R2ind498 R2ind498_inst(.x({x[737], x[736], x[735], x[734], x[733], x[732], x[35]}), .y(y[498]));
  R2ind499 R2ind499_inst(.x({x[737], x[736], x[735], x[734], x[733], x[732], x[35]}), .y(y[499]));
  R2ind500 R2ind500_inst(.x({x[743], x[742], x[741], x[740], x[739], x[738], x[35]}), .y(y[500]));
  R2ind501 R2ind501_inst(.x({x[743], x[742], x[741], x[740], x[739], x[738], x[35]}), .y(y[501]));
  R2ind502 R2ind502_inst(.x({x[743], x[742], x[741], x[740], x[739], x[738], x[35]}), .y(y[502]));
  R2ind503 R2ind503_inst(.x({x[743], x[742], x[741], x[740], x[739], x[738], x[35]}), .y(y[503]));
  R2ind504 R2ind504_inst(.x({x[749], x[748], x[747], x[746], x[745], x[744], x[35]}), .y(y[504]));
  R2ind505 R2ind505_inst(.x({x[749], x[748], x[747], x[746], x[745], x[744], x[35]}), .y(y[505]));
  R2ind506 R2ind506_inst(.x({x[749], x[748], x[747], x[746], x[745], x[744], x[35]}), .y(y[506]));
  R2ind507 R2ind507_inst(.x({x[749], x[748], x[747], x[746], x[745], x[744], x[35]}), .y(y[507]));
  R2ind508 R2ind508_inst(.x({x[755], x[754], x[753], x[752], x[751], x[750], x[35]}), .y(y[508]));
  R2ind509 R2ind509_inst(.x({x[755], x[754], x[753], x[752], x[751], x[750], x[35]}), .y(y[509]));
  R2ind510 R2ind510_inst(.x({x[755], x[754], x[753], x[752], x[751], x[750], x[35]}), .y(y[510]));
  R2ind511 R2ind511_inst(.x({x[755], x[754], x[753], x[752], x[751], x[750], x[35]}), .y(y[511]));
  R2ind512 R2ind512_inst(.x({x[761], x[760], x[759], x[758], x[757], x[756], x[35]}), .y(y[512]));
  R2ind513 R2ind513_inst(.x({x[761], x[760], x[759], x[758], x[757], x[756], x[35]}), .y(y[513]));
  R2ind514 R2ind514_inst(.x({x[761], x[760], x[759], x[758], x[757], x[756], x[35]}), .y(y[514]));
  R2ind515 R2ind515_inst(.x({x[761], x[760], x[759], x[758], x[757], x[756], x[35]}), .y(y[515]));
  R2ind516 R2ind516_inst(.x({x[767], x[766], x[765], x[764], x[763], x[762], x[35]}), .y(y[516]));
  R2ind517 R2ind517_inst(.x({x[767], x[766], x[765], x[764], x[763], x[762], x[35]}), .y(y[517]));
  R2ind518 R2ind518_inst(.x({x[767], x[766], x[765], x[764], x[763], x[762], x[35]}), .y(y[518]));
  R2ind519 R2ind519_inst(.x({x[767], x[766], x[765], x[764], x[763], x[762], x[35]}), .y(y[519]));
  R2ind520 R2ind520_inst(.x({x[773], x[772], x[771], x[770], x[769], x[768], x[35]}), .y(y[520]));
  R2ind521 R2ind521_inst(.x({x[773], x[772], x[771], x[770], x[769], x[768], x[35]}), .y(y[521]));
  R2ind522 R2ind522_inst(.x({x[773], x[772], x[771], x[770], x[769], x[768], x[35]}), .y(y[522]));
  R2ind523 R2ind523_inst(.x({x[773], x[772], x[771], x[770], x[769], x[768], x[35]}), .y(y[523]));
  R2ind524 R2ind524_inst(.x({x[779], x[778], x[777], x[776], x[775], x[774], x[35]}), .y(y[524]));
  R2ind525 R2ind525_inst(.x({x[779], x[778], x[777], x[776], x[775], x[774], x[35]}), .y(y[525]));
  R2ind526 R2ind526_inst(.x({x[779], x[778], x[777], x[776], x[775], x[774], x[35]}), .y(y[526]));
  R2ind527 R2ind527_inst(.x({x[779], x[778], x[777], x[776], x[775], x[774], x[35]}), .y(y[527]));
  R2ind528 R2ind528_inst(.x({x[785], x[784], x[783], x[782], x[781], x[780], x[35]}), .y(y[528]));
  R2ind529 R2ind529_inst(.x({x[785], x[784], x[783], x[782], x[781], x[780], x[35]}), .y(y[529]));
  R2ind530 R2ind530_inst(.x({x[785], x[784], x[783], x[782], x[781], x[780], x[35]}), .y(y[530]));
  R2ind531 R2ind531_inst(.x({x[785], x[784], x[783], x[782], x[781], x[780], x[35]}), .y(y[531]));
  R2ind532 R2ind532_inst(.x({x[791], x[790], x[789], x[788], x[787], x[786], x[35]}), .y(y[532]));
  R2ind533 R2ind533_inst(.x({x[791], x[790], x[789], x[788], x[787], x[786], x[35]}), .y(y[533]));
  R2ind534 R2ind534_inst(.x({x[791], x[790], x[789], x[788], x[787], x[786], x[35]}), .y(y[534]));
  R2ind535 R2ind535_inst(.x({x[791], x[790], x[789], x[788], x[787], x[786], x[35]}), .y(y[535]));
  R2ind536 R2ind536_inst(.x({x[797], x[796], x[795], x[794], x[793], x[792], x[35]}), .y(y[536]));
  R2ind537 R2ind537_inst(.x({x[797], x[796], x[795], x[794], x[793], x[792], x[35]}), .y(y[537]));
  R2ind538 R2ind538_inst(.x({x[797], x[796], x[795], x[794], x[793], x[792], x[35]}), .y(y[538]));
  R2ind539 R2ind539_inst(.x({x[797], x[796], x[795], x[794], x[793], x[792], x[35]}), .y(y[539]));
  R2ind540 R2ind540_inst(.x({x[803], x[802], x[801], x[800], x[799], x[798], x[35]}), .y(y[540]));
  R2ind541 R2ind541_inst(.x({x[803], x[802], x[801], x[800], x[799], x[798], x[35]}), .y(y[541]));
  R2ind542 R2ind542_inst(.x({x[803], x[802], x[801], x[800], x[799], x[798], x[35]}), .y(y[542]));
  R2ind543 R2ind543_inst(.x({x[803], x[802], x[801], x[800], x[799], x[798], x[35]}), .y(y[543]));
endmodule

