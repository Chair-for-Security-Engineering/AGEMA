/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* 16 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 17 register stage(s) in total */

module sbox_HPC2_BDDcudd_Pipeline_d1 (X_s0, clk, X_s1, Fresh, Y_s0, Y_s1);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [410:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_169 ;
    wire signal_170 ;
    wire signal_171 ;
    wire signal_172 ;
    wire signal_173 ;
    wire signal_174 ;
    wire signal_175 ;
    wire signal_176 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_182 ;
    wire signal_183 ;
    wire signal_184 ;
    wire signal_185 ;
    wire signal_186 ;
    wire signal_187 ;
    wire signal_188 ;
    wire signal_189 ;
    wire signal_190 ;
    wire signal_191 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_555 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;

    /* cells in depth 0 */

    /* cells in depth 1 */
    buf_clk cell_547 ( .C (clk), .D (X_s0[5]), .Q (signal_1392) ) ;
    buf_clk cell_549 ( .C (clk), .D (X_s1[5]), .Q (signal_1394) ) ;
    buf_clk cell_551 ( .C (clk), .D (X_s0[6]), .Q (signal_1396) ) ;
    buf_clk cell_553 ( .C (clk), .D (X_s1[6]), .Q (signal_1398) ) ;
    buf_clk cell_575 ( .C (clk), .D (X_s0[3]), .Q (signal_1420) ) ;
    buf_clk cell_579 ( .C (clk), .D (X_s1[3]), .Q (signal_1424) ) ;
    buf_clk cell_691 ( .C (clk), .D (X_s0[1]), .Q (signal_1536) ) ;
    buf_clk cell_699 ( .C (clk), .D (X_s1[1]), .Q (signal_1544) ) ;
    buf_clk cell_731 ( .C (clk), .D (X_s0[2]), .Q (signal_1576) ) ;
    buf_clk cell_741 ( .C (clk), .D (X_s1[2]), .Q (signal_1586) ) ;
    buf_clk cell_751 ( .C (clk), .D (X_s0[4]), .Q (signal_1596) ) ;
    buf_clk cell_763 ( .C (clk), .D (X_s1[4]), .Q (signal_1608) ) ;
    buf_clk cell_775 ( .C (clk), .D (X_s0[7]), .Q (signal_1620) ) ;
    buf_clk cell_789 ( .C (clk), .D (X_s1[7]), .Q (signal_1634) ) ;

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_136 ( .s ({X_s1[5], X_s0[5]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[0]), .c ({signal_555, signal_151}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_137 ( .s ({X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[1]), .c ({signal_557, signal_152}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_138 ( .s ({X_s1[5], X_s0[5]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[2]), .c ({signal_558, signal_153}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_139 ( .s ({X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[3]), .c ({signal_560, signal_154}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_140 ( .s ({X_s1[0], X_s0[0]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[4]), .c ({signal_561, signal_155}) ) ;
    buf_clk cell_548 ( .C (clk), .D (signal_1392), .Q (signal_1393) ) ;
    buf_clk cell_550 ( .C (clk), .D (signal_1394), .Q (signal_1395) ) ;
    buf_clk cell_552 ( .C (clk), .D (signal_1396), .Q (signal_1397) ) ;
    buf_clk cell_554 ( .C (clk), .D (signal_1398), .Q (signal_1399) ) ;
    buf_clk cell_576 ( .C (clk), .D (signal_1420), .Q (signal_1421) ) ;
    buf_clk cell_580 ( .C (clk), .D (signal_1424), .Q (signal_1425) ) ;
    buf_clk cell_692 ( .C (clk), .D (signal_1536), .Q (signal_1537) ) ;
    buf_clk cell_700 ( .C (clk), .D (signal_1544), .Q (signal_1545) ) ;
    buf_clk cell_732 ( .C (clk), .D (signal_1576), .Q (signal_1577) ) ;
    buf_clk cell_742 ( .C (clk), .D (signal_1586), .Q (signal_1587) ) ;
    buf_clk cell_752 ( .C (clk), .D (signal_1596), .Q (signal_1597) ) ;
    buf_clk cell_764 ( .C (clk), .D (signal_1608), .Q (signal_1609) ) ;
    buf_clk cell_776 ( .C (clk), .D (signal_1620), .Q (signal_1621) ) ;
    buf_clk cell_790 ( .C (clk), .D (signal_1634), .Q (signal_1635) ) ;

    /* cells in depth 3 */
    buf_clk cell_555 ( .C (clk), .D (signal_1397), .Q (signal_1400) ) ;
    buf_clk cell_557 ( .C (clk), .D (signal_1399), .Q (signal_1402) ) ;
    buf_clk cell_559 ( .C (clk), .D (signal_153), .Q (signal_1404) ) ;
    buf_clk cell_561 ( .C (clk), .D (signal_558), .Q (signal_1406) ) ;
    buf_clk cell_563 ( .C (clk), .D (signal_154), .Q (signal_1408) ) ;
    buf_clk cell_565 ( .C (clk), .D (signal_560), .Q (signal_1410) ) ;
    buf_clk cell_567 ( .C (clk), .D (signal_151), .Q (signal_1412) ) ;
    buf_clk cell_569 ( .C (clk), .D (signal_555), .Q (signal_1414) ) ;
    buf_clk cell_571 ( .C (clk), .D (signal_155), .Q (signal_1416) ) ;
    buf_clk cell_573 ( .C (clk), .D (signal_561), .Q (signal_1418) ) ;
    buf_clk cell_577 ( .C (clk), .D (signal_1421), .Q (signal_1422) ) ;
    buf_clk cell_581 ( .C (clk), .D (signal_1425), .Q (signal_1426) ) ;
    buf_clk cell_583 ( .C (clk), .D (signal_152), .Q (signal_1428) ) ;
    buf_clk cell_585 ( .C (clk), .D (signal_557), .Q (signal_1430) ) ;
    buf_clk cell_693 ( .C (clk), .D (signal_1537), .Q (signal_1538) ) ;
    buf_clk cell_701 ( .C (clk), .D (signal_1545), .Q (signal_1546) ) ;
    buf_clk cell_733 ( .C (clk), .D (signal_1577), .Q (signal_1578) ) ;
    buf_clk cell_743 ( .C (clk), .D (signal_1587), .Q (signal_1588) ) ;
    buf_clk cell_753 ( .C (clk), .D (signal_1597), .Q (signal_1598) ) ;
    buf_clk cell_765 ( .C (clk), .D (signal_1609), .Q (signal_1610) ) ;
    buf_clk cell_777 ( .C (clk), .D (signal_1621), .Q (signal_1622) ) ;
    buf_clk cell_791 ( .C (clk), .D (signal_1635), .Q (signal_1636) ) ;

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_141 ( .s ({signal_1395, signal_1393}), .b ({signal_561, signal_155}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[5]), .c ({signal_562, signal_156}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_142 ( .s ({signal_1395, signal_1393}), .b ({1'b0, 1'b1}), .a ({signal_561, signal_155}), .clk (clk), .r (Fresh[6]), .c ({signal_563, signal_157}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_143 ( .s ({signal_1395, signal_1393}), .b ({signal_560, signal_154}), .a ({signal_561, signal_155}), .clk (clk), .r (Fresh[7]), .c ({signal_564, signal_158}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_144 ( .s ({signal_1399, signal_1397}), .b ({signal_558, signal_153}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[8]), .c ({signal_565, signal_159}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_145 ( .s ({signal_1399, signal_1397}), .b ({signal_561, signal_155}), .a ({signal_560, signal_154}), .clk (clk), .r (Fresh[9]), .c ({signal_566, signal_160}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_146 ( .s ({signal_1399, signal_1397}), .b ({signal_558, signal_153}), .a ({signal_560, signal_154}), .clk (clk), .r (Fresh[10]), .c ({signal_567, signal_161}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_147 ( .s ({signal_1395, signal_1393}), .b ({signal_561, signal_155}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[11]), .c ({signal_568, signal_162}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_148 ( .s ({signal_1399, signal_1397}), .b ({signal_555, signal_151}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[12]), .c ({signal_569, signal_163}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_149 ( .s ({signal_1399, signal_1397}), .b ({signal_558, signal_153}), .a ({signal_561, signal_155}), .clk (clk), .r (Fresh[13]), .c ({signal_570, signal_164}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_150 ( .s ({signal_1395, signal_1393}), .b ({signal_560, signal_154}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[14]), .c ({signal_571, signal_165}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_151 ( .s ({signal_1399, signal_1397}), .b ({signal_555, signal_151}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[15]), .c ({signal_572, signal_166}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_152 ( .s ({signal_1399, signal_1397}), .b ({signal_560, signal_154}), .a ({signal_555, signal_151}), .clk (clk), .r (Fresh[16]), .c ({signal_573, signal_167}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_153 ( .s ({signal_1395, signal_1393}), .b ({1'b0, 1'b0}), .a ({signal_560, signal_154}), .clk (clk), .r (Fresh[17]), .c ({signal_574, signal_168}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_154 ( .s ({signal_1395, signal_1393}), .b ({1'b0, 1'b1}), .a ({signal_560, signal_154}), .clk (clk), .r (Fresh[18]), .c ({signal_575, signal_169}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_155 ( .s ({signal_1399, signal_1397}), .b ({1'b0, 1'b1}), .a ({signal_560, signal_154}), .clk (clk), .r (Fresh[19]), .c ({signal_576, signal_170}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_156 ( .s ({signal_1399, signal_1397}), .b ({signal_555, signal_151}), .a ({signal_560, signal_154}), .clk (clk), .r (Fresh[20]), .c ({signal_577, signal_171}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_157 ( .s ({signal_1399, signal_1397}), .b ({1'b0, 1'b0}), .a ({signal_560, signal_154}), .clk (clk), .r (Fresh[21]), .c ({signal_578, signal_172}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_158 ( .s ({signal_1399, signal_1397}), .b ({signal_558, signal_153}), .a ({signal_555, signal_151}), .clk (clk), .r (Fresh[22]), .c ({signal_579, signal_173}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_159 ( .s ({signal_1395, signal_1393}), .b ({signal_560, signal_154}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[23]), .c ({signal_580, signal_174}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_160 ( .s ({signal_1395, signal_1393}), .b ({1'b0, 1'b0}), .a ({signal_561, signal_155}), .clk (clk), .r (Fresh[24]), .c ({signal_581, signal_175}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_161 ( .s ({signal_1399, signal_1397}), .b ({1'b0, 1'b0}), .a ({signal_558, signal_153}), .clk (clk), .r (Fresh[25]), .c ({signal_582, signal_176}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_162 ( .s ({signal_1395, signal_1393}), .b ({signal_561, signal_155}), .a ({signal_560, signal_154}), .clk (clk), .r (Fresh[26]), .c ({signal_583, signal_177}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_163 ( .s ({signal_1399, signal_1397}), .b ({signal_555, signal_151}), .a ({signal_558, signal_153}), .clk (clk), .r (Fresh[27]), .c ({signal_584, signal_178}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_164 ( .s ({signal_1399, signal_1397}), .b ({signal_560, signal_154}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[28]), .c ({signal_585, signal_179}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_165 ( .s ({signal_1399, signal_1397}), .b ({1'b0, 1'b1}), .a ({signal_561, signal_155}), .clk (clk), .r (Fresh[29]), .c ({signal_586, signal_180}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_166 ( .s ({signal_1399, signal_1397}), .b ({1'b0, 1'b0}), .a ({signal_561, signal_155}), .clk (clk), .r (Fresh[30]), .c ({signal_587, signal_181}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_167 ( .s ({signal_1399, signal_1397}), .b ({signal_561, signal_155}), .a ({signal_555, signal_151}), .clk (clk), .r (Fresh[31]), .c ({signal_588, signal_182}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_168 ( .s ({signal_1399, signal_1397}), .b ({signal_558, signal_153}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[32]), .c ({signal_589, signal_183}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_169 ( .s ({signal_1399, signal_1397}), .b ({1'b0, 1'b1}), .a ({signal_555, signal_151}), .clk (clk), .r (Fresh[33]), .c ({signal_590, signal_184}) ) ;
    buf_clk cell_556 ( .C (clk), .D (signal_1400), .Q (signal_1401) ) ;
    buf_clk cell_558 ( .C (clk), .D (signal_1402), .Q (signal_1403) ) ;
    buf_clk cell_560 ( .C (clk), .D (signal_1404), .Q (signal_1405) ) ;
    buf_clk cell_562 ( .C (clk), .D (signal_1406), .Q (signal_1407) ) ;
    buf_clk cell_564 ( .C (clk), .D (signal_1408), .Q (signal_1409) ) ;
    buf_clk cell_566 ( .C (clk), .D (signal_1410), .Q (signal_1411) ) ;
    buf_clk cell_568 ( .C (clk), .D (signal_1412), .Q (signal_1413) ) ;
    buf_clk cell_570 ( .C (clk), .D (signal_1414), .Q (signal_1415) ) ;
    buf_clk cell_572 ( .C (clk), .D (signal_1416), .Q (signal_1417) ) ;
    buf_clk cell_574 ( .C (clk), .D (signal_1418), .Q (signal_1419) ) ;
    buf_clk cell_578 ( .C (clk), .D (signal_1422), .Q (signal_1423) ) ;
    buf_clk cell_582 ( .C (clk), .D (signal_1426), .Q (signal_1427) ) ;
    buf_clk cell_584 ( .C (clk), .D (signal_1428), .Q (signal_1429) ) ;
    buf_clk cell_586 ( .C (clk), .D (signal_1430), .Q (signal_1431) ) ;
    buf_clk cell_694 ( .C (clk), .D (signal_1538), .Q (signal_1539) ) ;
    buf_clk cell_702 ( .C (clk), .D (signal_1546), .Q (signal_1547) ) ;
    buf_clk cell_734 ( .C (clk), .D (signal_1578), .Q (signal_1579) ) ;
    buf_clk cell_744 ( .C (clk), .D (signal_1588), .Q (signal_1589) ) ;
    buf_clk cell_754 ( .C (clk), .D (signal_1598), .Q (signal_1599) ) ;
    buf_clk cell_766 ( .C (clk), .D (signal_1610), .Q (signal_1611) ) ;
    buf_clk cell_778 ( .C (clk), .D (signal_1622), .Q (signal_1623) ) ;
    buf_clk cell_792 ( .C (clk), .D (signal_1636), .Q (signal_1637) ) ;

    /* cells in depth 5 */
    buf_clk cell_587 ( .C (clk), .D (signal_1423), .Q (signal_1432) ) ;
    buf_clk cell_589 ( .C (clk), .D (signal_1427), .Q (signal_1434) ) ;
    buf_clk cell_591 ( .C (clk), .D (signal_1413), .Q (signal_1436) ) ;
    buf_clk cell_593 ( .C (clk), .D (signal_1415), .Q (signal_1438) ) ;
    buf_clk cell_595 ( .C (clk), .D (signal_1429), .Q (signal_1440) ) ;
    buf_clk cell_597 ( .C (clk), .D (signal_1431), .Q (signal_1442) ) ;
    buf_clk cell_599 ( .C (clk), .D (signal_182), .Q (signal_1444) ) ;
    buf_clk cell_601 ( .C (clk), .D (signal_588), .Q (signal_1446) ) ;
    buf_clk cell_603 ( .C (clk), .D (signal_175), .Q (signal_1448) ) ;
    buf_clk cell_605 ( .C (clk), .D (signal_581), .Q (signal_1450) ) ;
    buf_clk cell_607 ( .C (clk), .D (signal_177), .Q (signal_1452) ) ;
    buf_clk cell_609 ( .C (clk), .D (signal_583), .Q (signal_1454) ) ;
    buf_clk cell_611 ( .C (clk), .D (signal_169), .Q (signal_1456) ) ;
    buf_clk cell_613 ( .C (clk), .D (signal_575), .Q (signal_1458) ) ;
    buf_clk cell_615 ( .C (clk), .D (signal_178), .Q (signal_1460) ) ;
    buf_clk cell_617 ( .C (clk), .D (signal_584), .Q (signal_1462) ) ;
    buf_clk cell_619 ( .C (clk), .D (signal_167), .Q (signal_1464) ) ;
    buf_clk cell_621 ( .C (clk), .D (signal_573), .Q (signal_1466) ) ;
    buf_clk cell_623 ( .C (clk), .D (signal_171), .Q (signal_1468) ) ;
    buf_clk cell_625 ( .C (clk), .D (signal_577), .Q (signal_1470) ) ;
    buf_clk cell_627 ( .C (clk), .D (signal_183), .Q (signal_1472) ) ;
    buf_clk cell_629 ( .C (clk), .D (signal_589), .Q (signal_1474) ) ;
    buf_clk cell_631 ( .C (clk), .D (signal_184), .Q (signal_1476) ) ;
    buf_clk cell_633 ( .C (clk), .D (signal_590), .Q (signal_1478) ) ;
    buf_clk cell_635 ( .C (clk), .D (signal_180), .Q (signal_1480) ) ;
    buf_clk cell_637 ( .C (clk), .D (signal_586), .Q (signal_1482) ) ;
    buf_clk cell_639 ( .C (clk), .D (signal_172), .Q (signal_1484) ) ;
    buf_clk cell_641 ( .C (clk), .D (signal_578), .Q (signal_1486) ) ;
    buf_clk cell_643 ( .C (clk), .D (signal_163), .Q (signal_1488) ) ;
    buf_clk cell_645 ( .C (clk), .D (signal_569), .Q (signal_1490) ) ;
    buf_clk cell_647 ( .C (clk), .D (signal_168), .Q (signal_1492) ) ;
    buf_clk cell_649 ( .C (clk), .D (signal_574), .Q (signal_1494) ) ;
    buf_clk cell_651 ( .C (clk), .D (signal_170), .Q (signal_1496) ) ;
    buf_clk cell_653 ( .C (clk), .D (signal_576), .Q (signal_1498) ) ;
    buf_clk cell_655 ( .C (clk), .D (signal_161), .Q (signal_1500) ) ;
    buf_clk cell_657 ( .C (clk), .D (signal_567), .Q (signal_1502) ) ;
    buf_clk cell_659 ( .C (clk), .D (signal_164), .Q (signal_1504) ) ;
    buf_clk cell_661 ( .C (clk), .D (signal_570), .Q (signal_1506) ) ;
    buf_clk cell_663 ( .C (clk), .D (signal_162), .Q (signal_1508) ) ;
    buf_clk cell_665 ( .C (clk), .D (signal_568), .Q (signal_1510) ) ;
    buf_clk cell_667 ( .C (clk), .D (signal_173), .Q (signal_1512) ) ;
    buf_clk cell_669 ( .C (clk), .D (signal_579), .Q (signal_1514) ) ;
    buf_clk cell_671 ( .C (clk), .D (signal_158), .Q (signal_1516) ) ;
    buf_clk cell_673 ( .C (clk), .D (signal_564), .Q (signal_1518) ) ;
    buf_clk cell_675 ( .C (clk), .D (signal_181), .Q (signal_1520) ) ;
    buf_clk cell_677 ( .C (clk), .D (signal_587), .Q (signal_1522) ) ;
    buf_clk cell_679 ( .C (clk), .D (signal_176), .Q (signal_1524) ) ;
    buf_clk cell_681 ( .C (clk), .D (signal_582), .Q (signal_1526) ) ;
    buf_clk cell_683 ( .C (clk), .D (signal_157), .Q (signal_1528) ) ;
    buf_clk cell_685 ( .C (clk), .D (signal_563), .Q (signal_1530) ) ;
    buf_clk cell_687 ( .C (clk), .D (signal_166), .Q (signal_1532) ) ;
    buf_clk cell_689 ( .C (clk), .D (signal_572), .Q (signal_1534) ) ;
    buf_clk cell_695 ( .C (clk), .D (signal_1539), .Q (signal_1540) ) ;
    buf_clk cell_703 ( .C (clk), .D (signal_1547), .Q (signal_1548) ) ;
    buf_clk cell_735 ( .C (clk), .D (signal_1579), .Q (signal_1580) ) ;
    buf_clk cell_745 ( .C (clk), .D (signal_1589), .Q (signal_1590) ) ;
    buf_clk cell_755 ( .C (clk), .D (signal_1599), .Q (signal_1600) ) ;
    buf_clk cell_767 ( .C (clk), .D (signal_1611), .Q (signal_1612) ) ;
    buf_clk cell_779 ( .C (clk), .D (signal_1623), .Q (signal_1624) ) ;
    buf_clk cell_793 ( .C (clk), .D (signal_1637), .Q (signal_1638) ) ;

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_170 ( .s ({signal_1403, signal_1401}), .b ({signal_562, signal_156}), .a ({signal_1407, signal_1405}), .clk (clk), .r (Fresh[34]), .c ({signal_591, signal_185}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_171 ( .s ({signal_1403, signal_1401}), .b ({signal_581, signal_175}), .a ({signal_574, signal_168}), .clk (clk), .r (Fresh[35]), .c ({signal_592, signal_186}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_172 ( .s ({signal_1403, signal_1401}), .b ({signal_574, signal_168}), .a ({signal_564, signal_158}), .clk (clk), .r (Fresh[36]), .c ({signal_593, signal_187}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_173 ( .s ({signal_1403, signal_1401}), .b ({signal_575, signal_169}), .a ({signal_571, signal_165}), .clk (clk), .r (Fresh[37]), .c ({signal_594, signal_188}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_174 ( .s ({signal_1403, signal_1401}), .b ({signal_574, signal_168}), .a ({signal_575, signal_169}), .clk (clk), .r (Fresh[38]), .c ({signal_595, signal_189}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_175 ( .s ({signal_1403, signal_1401}), .b ({signal_1411, signal_1409}), .a ({signal_583, signal_177}), .clk (clk), .r (Fresh[39]), .c ({signal_596, signal_190}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_176 ( .s ({signal_1403, signal_1401}), .b ({signal_1407, signal_1405}), .a ({signal_571, signal_165}), .clk (clk), .r (Fresh[40]), .c ({signal_597, signal_191}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_177 ( .s ({signal_1403, signal_1401}), .b ({signal_1407, signal_1405}), .a ({signal_580, signal_174}), .clk (clk), .r (Fresh[41]), .c ({signal_598, signal_192}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_178 ( .s ({signal_1403, signal_1401}), .b ({signal_1415, signal_1413}), .a ({signal_581, signal_175}), .clk (clk), .r (Fresh[42]), .c ({signal_599, signal_193}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_179 ( .s ({signal_1403, signal_1401}), .b ({1'b0, 1'b0}), .a ({signal_574, signal_168}), .clk (clk), .r (Fresh[43]), .c ({signal_600, signal_194}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_180 ( .s ({signal_1403, signal_1401}), .b ({signal_580, signal_174}), .a ({signal_1419, signal_1417}), .clk (clk), .r (Fresh[44]), .c ({signal_601, signal_195}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_181 ( .s ({signal_1403, signal_1401}), .b ({signal_575, signal_169}), .a ({signal_574, signal_168}), .clk (clk), .r (Fresh[45]), .c ({signal_602, signal_196}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_182 ( .s ({signal_1403, signal_1401}), .b ({signal_580, signal_174}), .a ({signal_563, signal_157}), .clk (clk), .r (Fresh[46]), .c ({signal_603, signal_197}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_183 ( .s ({signal_1403, signal_1401}), .b ({signal_580, signal_174}), .a ({signal_581, signal_175}), .clk (clk), .r (Fresh[47]), .c ({signal_604, signal_198}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_184 ( .s ({signal_1403, signal_1401}), .b ({signal_580, signal_174}), .a ({signal_562, signal_156}), .clk (clk), .r (Fresh[48]), .c ({signal_605, signal_199}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_185 ( .s ({signal_1403, signal_1401}), .b ({signal_574, signal_168}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[49]), .c ({signal_606, signal_200}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_186 ( .s ({signal_1403, signal_1401}), .b ({signal_1411, signal_1409}), .a ({signal_564, signal_158}), .clk (clk), .r (Fresh[50]), .c ({signal_607, signal_201}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_187 ( .s ({signal_1403, signal_1401}), .b ({signal_563, signal_157}), .a ({signal_571, signal_165}), .clk (clk), .r (Fresh[51]), .c ({signal_608, signal_202}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_188 ( .s ({signal_1403, signal_1401}), .b ({signal_575, signal_169}), .a ({signal_568, signal_162}), .clk (clk), .r (Fresh[52]), .c ({signal_609, signal_203}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_189 ( .s ({signal_1403, signal_1401}), .b ({signal_562, signal_156}), .a ({signal_1419, signal_1417}), .clk (clk), .r (Fresh[53]), .c ({signal_610, signal_204}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_190 ( .s ({signal_1403, signal_1401}), .b ({signal_1411, signal_1409}), .a ({signal_575, signal_169}), .clk (clk), .r (Fresh[54]), .c ({signal_611, signal_205}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_191 ( .s ({signal_1403, signal_1401}), .b ({signal_568, signal_162}), .a ({signal_1415, signal_1413}), .clk (clk), .r (Fresh[55]), .c ({signal_612, signal_206}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_192 ( .s ({signal_1403, signal_1401}), .b ({signal_581, signal_175}), .a ({signal_1415, signal_1413}), .clk (clk), .r (Fresh[56]), .c ({signal_613, signal_207}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_193 ( .s ({signal_1403, signal_1401}), .b ({signal_580, signal_174}), .a ({signal_575, signal_169}), .clk (clk), .r (Fresh[57]), .c ({signal_614, signal_208}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_194 ( .s ({signal_1403, signal_1401}), .b ({signal_568, signal_162}), .a ({signal_583, signal_177}), .clk (clk), .r (Fresh[58]), .c ({signal_615, signal_209}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_195 ( .s ({signal_1403, signal_1401}), .b ({1'b0, 1'b1}), .a ({signal_563, signal_157}), .clk (clk), .r (Fresh[59]), .c ({signal_616, signal_210}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_196 ( .s ({signal_1403, signal_1401}), .b ({signal_580, signal_174}), .a ({signal_564, signal_158}), .clk (clk), .r (Fresh[60]), .c ({signal_617, signal_211}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_197 ( .s ({signal_1403, signal_1401}), .b ({signal_1419, signal_1417}), .a ({signal_580, signal_174}), .clk (clk), .r (Fresh[61]), .c ({signal_618, signal_212}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_198 ( .s ({signal_1403, signal_1401}), .b ({signal_564, signal_158}), .a ({signal_1407, signal_1405}), .clk (clk), .r (Fresh[62]), .c ({signal_619, signal_213}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_199 ( .s ({signal_1403, signal_1401}), .b ({signal_564, signal_158}), .a ({signal_574, signal_168}), .clk (clk), .r (Fresh[63]), .c ({signal_620, signal_214}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_200 ( .s ({signal_1403, signal_1401}), .b ({signal_574, signal_168}), .a ({signal_583, signal_177}), .clk (clk), .r (Fresh[64]), .c ({signal_621, signal_215}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_201 ( .s ({signal_1403, signal_1401}), .b ({signal_581, signal_175}), .a ({signal_564, signal_158}), .clk (clk), .r (Fresh[65]), .c ({signal_622, signal_216}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_202 ( .s ({signal_1403, signal_1401}), .b ({signal_571, signal_165}), .a ({signal_581, signal_175}), .clk (clk), .r (Fresh[66]), .c ({signal_623, signal_217}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_203 ( .s ({signal_1403, signal_1401}), .b ({signal_575, signal_169}), .a ({signal_1407, signal_1405}), .clk (clk), .r (Fresh[67]), .c ({signal_624, signal_218}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_204 ( .s ({signal_1403, signal_1401}), .b ({signal_1419, signal_1417}), .a ({signal_575, signal_169}), .clk (clk), .r (Fresh[68]), .c ({signal_625, signal_219}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_205 ( .s ({signal_1403, signal_1401}), .b ({signal_1419, signal_1417}), .a ({signal_564, signal_158}), .clk (clk), .r (Fresh[69]), .c ({signal_626, signal_220}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_206 ( .s ({signal_1403, signal_1401}), .b ({signal_574, signal_168}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[70]), .c ({signal_627, signal_221}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_207 ( .s ({signal_1403, signal_1401}), .b ({signal_562, signal_156}), .a ({signal_580, signal_174}), .clk (clk), .r (Fresh[71]), .c ({signal_628, signal_222}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_208 ( .s ({signal_1403, signal_1401}), .b ({signal_564, signal_158}), .a ({signal_1419, signal_1417}), .clk (clk), .r (Fresh[72]), .c ({signal_629, signal_223}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_209 ( .s ({signal_1403, signal_1401}), .b ({signal_583, signal_177}), .a ({signal_1411, signal_1409}), .clk (clk), .r (Fresh[73]), .c ({signal_630, signal_224}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_210 ( .s ({signal_1403, signal_1401}), .b ({signal_562, signal_156}), .a ({signal_568, signal_162}), .clk (clk), .r (Fresh[74]), .c ({signal_631, signal_225}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_211 ( .s ({signal_1403, signal_1401}), .b ({signal_562, signal_156}), .a ({signal_581, signal_175}), .clk (clk), .r (Fresh[75]), .c ({signal_632, signal_226}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_212 ( .s ({signal_1403, signal_1401}), .b ({signal_564, signal_158}), .a ({signal_571, signal_165}), .clk (clk), .r (Fresh[76]), .c ({signal_633, signal_227}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_213 ( .s ({signal_1403, signal_1401}), .b ({signal_1407, signal_1405}), .a ({signal_583, signal_177}), .clk (clk), .r (Fresh[77]), .c ({signal_634, signal_228}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_214 ( .s ({signal_1403, signal_1401}), .b ({signal_563, signal_157}), .a ({signal_583, signal_177}), .clk (clk), .r (Fresh[78]), .c ({signal_635, signal_229}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_215 ( .s ({signal_1403, signal_1401}), .b ({1'b0, 1'b0}), .a ({signal_564, signal_158}), .clk (clk), .r (Fresh[79]), .c ({signal_636, signal_230}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_216 ( .s ({signal_1403, signal_1401}), .b ({signal_562, signal_156}), .a ({signal_1411, signal_1409}), .clk (clk), .r (Fresh[80]), .c ({signal_637, signal_231}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_217 ( .s ({signal_1403, signal_1401}), .b ({signal_575, signal_169}), .a ({signal_1411, signal_1409}), .clk (clk), .r (Fresh[81]), .c ({signal_638, signal_232}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_218 ( .s ({signal_1403, signal_1401}), .b ({1'b0, 1'b1}), .a ({signal_564, signal_158}), .clk (clk), .r (Fresh[82]), .c ({signal_639, signal_233}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_219 ( .s ({signal_1403, signal_1401}), .b ({signal_575, signal_169}), .a ({signal_580, signal_174}), .clk (clk), .r (Fresh[83]), .c ({signal_640, signal_234}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_220 ( .s ({signal_1403, signal_1401}), .b ({signal_1415, signal_1413}), .a ({signal_574, signal_168}), .clk (clk), .r (Fresh[84]), .c ({signal_641, signal_235}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_221 ( .s ({signal_1403, signal_1401}), .b ({1'b0, 1'b0}), .a ({signal_563, signal_157}), .clk (clk), .r (Fresh[85]), .c ({signal_642, signal_236}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_222 ( .s ({signal_1403, signal_1401}), .b ({signal_583, signal_177}), .a ({signal_571, signal_165}), .clk (clk), .r (Fresh[86]), .c ({signal_643, signal_237}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_223 ( .s ({signal_1403, signal_1401}), .b ({signal_568, signal_162}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[87]), .c ({signal_644, signal_238}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_224 ( .s ({signal_1403, signal_1401}), .b ({signal_568, signal_162}), .a ({signal_562, signal_156}), .clk (clk), .r (Fresh[88]), .c ({signal_645, signal_239}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_225 ( .s ({signal_1403, signal_1401}), .b ({signal_1419, signal_1417}), .a ({signal_571, signal_165}), .clk (clk), .r (Fresh[89]), .c ({signal_646, signal_240}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_226 ( .s ({signal_1403, signal_1401}), .b ({signal_575, signal_169}), .a ({signal_562, signal_156}), .clk (clk), .r (Fresh[90]), .c ({signal_647, signal_241}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_227 ( .s ({signal_1403, signal_1401}), .b ({signal_571, signal_165}), .a ({signal_1411, signal_1409}), .clk (clk), .r (Fresh[91]), .c ({signal_648, signal_242}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_228 ( .s ({signal_1403, signal_1401}), .b ({signal_575, signal_169}), .a ({signal_1415, signal_1413}), .clk (clk), .r (Fresh[92]), .c ({signal_649, signal_243}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_229 ( .s ({signal_1427, signal_1423}), .b ({signal_566, signal_160}), .a ({signal_582, signal_176}), .clk (clk), .r (Fresh[93]), .c ({signal_651, signal_244}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_230 ( .s ({signal_1403, signal_1401}), .b ({1'b0, 1'b1}), .a ({signal_568, signal_162}), .clk (clk), .r (Fresh[94]), .c ({signal_652, signal_245}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_231 ( .s ({signal_1403, signal_1401}), .b ({signal_574, signal_168}), .a ({signal_580, signal_174}), .clk (clk), .r (Fresh[95]), .c ({signal_653, signal_246}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_232 ( .s ({signal_1403, signal_1401}), .b ({signal_583, signal_177}), .a ({signal_563, signal_157}), .clk (clk), .r (Fresh[96]), .c ({signal_654, signal_247}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_233 ( .s ({signal_1403, signal_1401}), .b ({1'b0, 1'b1}), .a ({signal_574, signal_168}), .clk (clk), .r (Fresh[97]), .c ({signal_655, signal_248}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_234 ( .s ({signal_1403, signal_1401}), .b ({signal_581, signal_175}), .a ({signal_575, signal_169}), .clk (clk), .r (Fresh[98]), .c ({signal_656, signal_249}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_235 ( .s ({signal_1403, signal_1401}), .b ({signal_568, signal_162}), .a ({signal_563, signal_157}), .clk (clk), .r (Fresh[99]), .c ({signal_657, signal_250}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_236 ( .s ({signal_1403, signal_1401}), .b ({signal_581, signal_175}), .a ({signal_562, signal_156}), .clk (clk), .r (Fresh[100]), .c ({signal_658, signal_251}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_237 ( .s ({signal_1403, signal_1401}), .b ({signal_580, signal_174}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[101]), .c ({signal_659, signal_252}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_238 ( .s ({signal_1403, signal_1401}), .b ({1'b0, 1'b1}), .a ({signal_583, signal_177}), .clk (clk), .r (Fresh[102]), .c ({signal_660, signal_253}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_239 ( .s ({signal_1403, signal_1401}), .b ({signal_563, signal_157}), .a ({signal_1411, signal_1409}), .clk (clk), .r (Fresh[103]), .c ({signal_661, signal_254}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_240 ( .s ({signal_1403, signal_1401}), .b ({signal_574, signal_168}), .a ({signal_581, signal_175}), .clk (clk), .r (Fresh[104]), .c ({signal_662, signal_255}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_241 ( .s ({signal_1403, signal_1401}), .b ({signal_1411, signal_1409}), .a ({signal_563, signal_157}), .clk (clk), .r (Fresh[105]), .c ({signal_663, signal_256}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_242 ( .s ({signal_1403, signal_1401}), .b ({signal_1419, signal_1417}), .a ({signal_562, signal_156}), .clk (clk), .r (Fresh[106]), .c ({signal_664, signal_257}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_243 ( .s ({signal_1403, signal_1401}), .b ({signal_583, signal_177}), .a ({signal_564, signal_158}), .clk (clk), .r (Fresh[107]), .c ({signal_665, signal_258}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_244 ( .s ({signal_1403, signal_1401}), .b ({signal_562, signal_156}), .a ({signal_575, signal_169}), .clk (clk), .r (Fresh[108]), .c ({signal_666, signal_259}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_245 ( .s ({signal_1403, signal_1401}), .b ({signal_581, signal_175}), .a ({signal_1419, signal_1417}), .clk (clk), .r (Fresh[109]), .c ({signal_667, signal_260}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_246 ( .s ({signal_1403, signal_1401}), .b ({signal_580, signal_174}), .a ({signal_1411, signal_1409}), .clk (clk), .r (Fresh[110]), .c ({signal_668, signal_261}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_247 ( .s ({signal_1403, signal_1401}), .b ({signal_1415, signal_1413}), .a ({signal_571, signal_165}), .clk (clk), .r (Fresh[111]), .c ({signal_669, signal_262}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_248 ( .s ({signal_1403, signal_1401}), .b ({signal_571, signal_165}), .a ({signal_574, signal_168}), .clk (clk), .r (Fresh[112]), .c ({signal_670, signal_263}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_249 ( .s ({signal_1403, signal_1401}), .b ({signal_563, signal_157}), .a ({signal_1415, signal_1413}), .clk (clk), .r (Fresh[113]), .c ({signal_671, signal_264}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_250 ( .s ({signal_1403, signal_1401}), .b ({signal_568, signal_162}), .a ({signal_1407, signal_1405}), .clk (clk), .r (Fresh[114]), .c ({signal_672, signal_265}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_251 ( .s ({signal_1403, signal_1401}), .b ({signal_1407, signal_1405}), .a ({signal_562, signal_156}), .clk (clk), .r (Fresh[115]), .c ({signal_673, signal_266}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_252 ( .s ({signal_1403, signal_1401}), .b ({signal_1419, signal_1417}), .a ({signal_583, signal_177}), .clk (clk), .r (Fresh[116]), .c ({signal_674, signal_267}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_253 ( .s ({signal_1403, signal_1401}), .b ({signal_1415, signal_1413}), .a ({signal_568, signal_162}), .clk (clk), .r (Fresh[117]), .c ({signal_675, signal_268}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_254 ( .s ({signal_1403, signal_1401}), .b ({signal_1415, signal_1413}), .a ({signal_575, signal_169}), .clk (clk), .r (Fresh[118]), .c ({signal_676, signal_269}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_255 ( .s ({signal_1403, signal_1401}), .b ({signal_571, signal_165}), .a ({signal_564, signal_158}), .clk (clk), .r (Fresh[119]), .c ({signal_677, signal_270}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_256 ( .s ({signal_1403, signal_1401}), .b ({signal_564, signal_158}), .a ({signal_562, signal_156}), .clk (clk), .r (Fresh[120]), .c ({signal_678, signal_271}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_257 ( .s ({signal_1403, signal_1401}), .b ({signal_574, signal_168}), .a ({signal_1411, signal_1409}), .clk (clk), .r (Fresh[121]), .c ({signal_679, signal_272}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_258 ( .s ({signal_1403, signal_1401}), .b ({signal_575, signal_169}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[122]), .c ({signal_680, signal_273}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_259 ( .s ({signal_1427, signal_1423}), .b ({signal_1419, signal_1417}), .a ({signal_570, signal_164}), .clk (clk), .r (Fresh[123]), .c ({signal_681, signal_274}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_260 ( .s ({signal_1403, signal_1401}), .b ({signal_563, signal_157}), .a ({signal_1407, signal_1405}), .clk (clk), .r (Fresh[124]), .c ({signal_682, signal_275}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_261 ( .s ({signal_1403, signal_1401}), .b ({signal_580, signal_174}), .a ({signal_1407, signal_1405}), .clk (clk), .r (Fresh[125]), .c ({signal_683, signal_276}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_262 ( .s ({signal_1403, signal_1401}), .b ({signal_581, signal_175}), .a ({signal_568, signal_162}), .clk (clk), .r (Fresh[126]), .c ({signal_684, signal_277}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_263 ( .s ({signal_1403, signal_1401}), .b ({signal_583, signal_177}), .a ({signal_568, signal_162}), .clk (clk), .r (Fresh[127]), .c ({signal_685, signal_278}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_264 ( .s ({signal_1403, signal_1401}), .b ({signal_580, signal_174}), .a ({signal_571, signal_165}), .clk (clk), .r (Fresh[128]), .c ({signal_686, signal_279}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_265 ( .s ({signal_1403, signal_1401}), .b ({signal_583, signal_177}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[129]), .c ({signal_687, signal_280}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_266 ( .s ({signal_1403, signal_1401}), .b ({signal_581, signal_175}), .a ({signal_580, signal_174}), .clk (clk), .r (Fresh[130]), .c ({signal_688, signal_281}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_267 ( .s ({signal_1427, signal_1423}), .b ({signal_562, signal_156}), .a ({signal_1431, signal_1429}), .clk (clk), .r (Fresh[131]), .c ({signal_689, signal_282}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_268 ( .s ({signal_1403, signal_1401}), .b ({signal_563, signal_157}), .a ({signal_574, signal_168}), .clk (clk), .r (Fresh[132]), .c ({signal_690, signal_283}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_269 ( .s ({signal_1403, signal_1401}), .b ({signal_568, signal_162}), .a ({signal_581, signal_175}), .clk (clk), .r (Fresh[133]), .c ({signal_691, signal_284}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_270 ( .s ({signal_1403, signal_1401}), .b ({signal_575, signal_169}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[134]), .c ({signal_692, signal_285}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_271 ( .s ({signal_1403, signal_1401}), .b ({1'b0, 1'b0}), .a ({signal_562, signal_156}), .clk (clk), .r (Fresh[135]), .c ({signal_693, signal_286}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_272 ( .s ({signal_1403, signal_1401}), .b ({signal_562, signal_156}), .a ({signal_564, signal_158}), .clk (clk), .r (Fresh[136]), .c ({signal_694, signal_287}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_273 ( .s ({signal_1403, signal_1401}), .b ({signal_1411, signal_1409}), .a ({signal_571, signal_165}), .clk (clk), .r (Fresh[137]), .c ({signal_695, signal_288}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_274 ( .s ({signal_1403, signal_1401}), .b ({signal_568, signal_162}), .a ({signal_571, signal_165}), .clk (clk), .r (Fresh[138]), .c ({signal_696, signal_289}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_275 ( .s ({signal_1403, signal_1401}), .b ({signal_583, signal_177}), .a ({signal_580, signal_174}), .clk (clk), .r (Fresh[139]), .c ({signal_697, signal_290}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_276 ( .s ({signal_1403, signal_1401}), .b ({signal_562, signal_156}), .a ({signal_583, signal_177}), .clk (clk), .r (Fresh[140]), .c ({signal_698, signal_291}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_277 ( .s ({signal_1403, signal_1401}), .b ({signal_571, signal_165}), .a ({signal_1415, signal_1413}), .clk (clk), .r (Fresh[141]), .c ({signal_699, signal_292}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_278 ( .s ({signal_1403, signal_1401}), .b ({signal_581, signal_175}), .a ({signal_563, signal_157}), .clk (clk), .r (Fresh[142]), .c ({signal_700, signal_293}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_279 ( .s ({signal_1403, signal_1401}), .b ({signal_575, signal_169}), .a ({signal_564, signal_158}), .clk (clk), .r (Fresh[143]), .c ({signal_701, signal_294}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_280 ( .s ({signal_1403, signal_1401}), .b ({signal_580, signal_174}), .a ({signal_568, signal_162}), .clk (clk), .r (Fresh[144]), .c ({signal_702, signal_295}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_281 ( .s ({signal_1403, signal_1401}), .b ({1'b0, 1'b1}), .a ({signal_575, signal_169}), .clk (clk), .r (Fresh[145]), .c ({signal_703, signal_296}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_282 ( .s ({signal_1403, signal_1401}), .b ({signal_580, signal_174}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[146]), .c ({signal_704, signal_297}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_283 ( .s ({signal_1403, signal_1401}), .b ({1'b0, 1'b1}), .a ({signal_571, signal_165}), .clk (clk), .r (Fresh[147]), .c ({signal_705, signal_298}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_284 ( .s ({signal_1427, signal_1423}), .b ({signal_588, signal_182}), .a ({signal_1407, signal_1405}), .clk (clk), .r (Fresh[148]), .c ({signal_706, signal_299}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_285 ( .s ({signal_1403, signal_1401}), .b ({signal_583, signal_177}), .a ({signal_581, signal_175}), .clk (clk), .r (Fresh[149]), .c ({signal_707, signal_300}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_286 ( .s ({signal_1403, signal_1401}), .b ({signal_564, signal_158}), .a ({signal_568, signal_162}), .clk (clk), .r (Fresh[150]), .c ({signal_708, signal_301}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_287 ( .s ({signal_1427, signal_1423}), .b ({signal_565, signal_159}), .a ({signal_567, signal_161}), .clk (clk), .r (Fresh[151]), .c ({signal_709, signal_302}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_288 ( .s ({signal_1403, signal_1401}), .b ({signal_575, signal_169}), .a ({signal_583, signal_177}), .clk (clk), .r (Fresh[152]), .c ({signal_710, signal_303}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_289 ( .s ({signal_1403, signal_1401}), .b ({signal_1407, signal_1405}), .a ({signal_574, signal_168}), .clk (clk), .r (Fresh[153]), .c ({signal_711, signal_304}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_290 ( .s ({signal_1403, signal_1401}), .b ({signal_575, signal_169}), .a ({signal_1419, signal_1417}), .clk (clk), .r (Fresh[154]), .c ({signal_712, signal_305}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_291 ( .s ({signal_1427, signal_1423}), .b ({signal_585, signal_179}), .a ({signal_562, signal_156}), .clk (clk), .r (Fresh[155]), .c ({signal_713, signal_306}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_292 ( .s ({signal_1403, signal_1401}), .b ({signal_1419, signal_1417}), .a ({signal_574, signal_168}), .clk (clk), .r (Fresh[156]), .c ({signal_714, signal_307}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_293 ( .s ({signal_1403, signal_1401}), .b ({signal_574, signal_168}), .a ({signal_571, signal_165}), .clk (clk), .r (Fresh[157]), .c ({signal_715, signal_308}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_294 ( .s ({signal_1403, signal_1401}), .b ({signal_1415, signal_1413}), .a ({signal_583, signal_177}), .clk (clk), .r (Fresh[158]), .c ({signal_716, signal_309}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_295 ( .s ({signal_1403, signal_1401}), .b ({signal_574, signal_168}), .a ({signal_568, signal_162}), .clk (clk), .r (Fresh[159]), .c ({signal_717, signal_310}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_296 ( .s ({signal_1403, signal_1401}), .b ({signal_1407, signal_1405}), .a ({signal_575, signal_169}), .clk (clk), .r (Fresh[160]), .c ({signal_718, signal_311}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_297 ( .s ({signal_1403, signal_1401}), .b ({signal_568, signal_162}), .a ({signal_580, signal_174}), .clk (clk), .r (Fresh[161]), .c ({signal_719, signal_312}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_298 ( .s ({signal_1403, signal_1401}), .b ({signal_564, signal_158}), .a ({signal_580, signal_174}), .clk (clk), .r (Fresh[162]), .c ({signal_720, signal_313}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_299 ( .s ({signal_1403, signal_1401}), .b ({signal_1411, signal_1409}), .a ({signal_562, signal_156}), .clk (clk), .r (Fresh[163]), .c ({signal_721, signal_314}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_300 ( .s ({signal_1403, signal_1401}), .b ({signal_1415, signal_1413}), .a ({signal_564, signal_158}), .clk (clk), .r (Fresh[164]), .c ({signal_722, signal_315}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_301 ( .s ({signal_1403, signal_1401}), .b ({1'b0, 1'b1}), .a ({signal_580, signal_174}), .clk (clk), .r (Fresh[165]), .c ({signal_723, signal_316}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_302 ( .s ({signal_1403, signal_1401}), .b ({signal_580, signal_174}), .a ({signal_574, signal_168}), .clk (clk), .r (Fresh[166]), .c ({signal_724, signal_317}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_303 ( .s ({signal_1403, signal_1401}), .b ({signal_571, signal_165}), .a ({signal_575, signal_169}), .clk (clk), .r (Fresh[167]), .c ({signal_725, signal_318}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_304 ( .s ({signal_1403, signal_1401}), .b ({signal_581, signal_175}), .a ({signal_1407, signal_1405}), .clk (clk), .r (Fresh[168]), .c ({signal_726, signal_319}) ) ;
    buf_clk cell_588 ( .C (clk), .D (signal_1432), .Q (signal_1433) ) ;
    buf_clk cell_590 ( .C (clk), .D (signal_1434), .Q (signal_1435) ) ;
    buf_clk cell_592 ( .C (clk), .D (signal_1436), .Q (signal_1437) ) ;
    buf_clk cell_594 ( .C (clk), .D (signal_1438), .Q (signal_1439) ) ;
    buf_clk cell_596 ( .C (clk), .D (signal_1440), .Q (signal_1441) ) ;
    buf_clk cell_598 ( .C (clk), .D (signal_1442), .Q (signal_1443) ) ;
    buf_clk cell_600 ( .C (clk), .D (signal_1444), .Q (signal_1445) ) ;
    buf_clk cell_602 ( .C (clk), .D (signal_1446), .Q (signal_1447) ) ;
    buf_clk cell_604 ( .C (clk), .D (signal_1448), .Q (signal_1449) ) ;
    buf_clk cell_606 ( .C (clk), .D (signal_1450), .Q (signal_1451) ) ;
    buf_clk cell_608 ( .C (clk), .D (signal_1452), .Q (signal_1453) ) ;
    buf_clk cell_610 ( .C (clk), .D (signal_1454), .Q (signal_1455) ) ;
    buf_clk cell_612 ( .C (clk), .D (signal_1456), .Q (signal_1457) ) ;
    buf_clk cell_614 ( .C (clk), .D (signal_1458), .Q (signal_1459) ) ;
    buf_clk cell_616 ( .C (clk), .D (signal_1460), .Q (signal_1461) ) ;
    buf_clk cell_618 ( .C (clk), .D (signal_1462), .Q (signal_1463) ) ;
    buf_clk cell_620 ( .C (clk), .D (signal_1464), .Q (signal_1465) ) ;
    buf_clk cell_622 ( .C (clk), .D (signal_1466), .Q (signal_1467) ) ;
    buf_clk cell_624 ( .C (clk), .D (signal_1468), .Q (signal_1469) ) ;
    buf_clk cell_626 ( .C (clk), .D (signal_1470), .Q (signal_1471) ) ;
    buf_clk cell_628 ( .C (clk), .D (signal_1472), .Q (signal_1473) ) ;
    buf_clk cell_630 ( .C (clk), .D (signal_1474), .Q (signal_1475) ) ;
    buf_clk cell_632 ( .C (clk), .D (signal_1476), .Q (signal_1477) ) ;
    buf_clk cell_634 ( .C (clk), .D (signal_1478), .Q (signal_1479) ) ;
    buf_clk cell_636 ( .C (clk), .D (signal_1480), .Q (signal_1481) ) ;
    buf_clk cell_638 ( .C (clk), .D (signal_1482), .Q (signal_1483) ) ;
    buf_clk cell_640 ( .C (clk), .D (signal_1484), .Q (signal_1485) ) ;
    buf_clk cell_642 ( .C (clk), .D (signal_1486), .Q (signal_1487) ) ;
    buf_clk cell_644 ( .C (clk), .D (signal_1488), .Q (signal_1489) ) ;
    buf_clk cell_646 ( .C (clk), .D (signal_1490), .Q (signal_1491) ) ;
    buf_clk cell_648 ( .C (clk), .D (signal_1492), .Q (signal_1493) ) ;
    buf_clk cell_650 ( .C (clk), .D (signal_1494), .Q (signal_1495) ) ;
    buf_clk cell_652 ( .C (clk), .D (signal_1496), .Q (signal_1497) ) ;
    buf_clk cell_654 ( .C (clk), .D (signal_1498), .Q (signal_1499) ) ;
    buf_clk cell_656 ( .C (clk), .D (signal_1500), .Q (signal_1501) ) ;
    buf_clk cell_658 ( .C (clk), .D (signal_1502), .Q (signal_1503) ) ;
    buf_clk cell_660 ( .C (clk), .D (signal_1504), .Q (signal_1505) ) ;
    buf_clk cell_662 ( .C (clk), .D (signal_1506), .Q (signal_1507) ) ;
    buf_clk cell_664 ( .C (clk), .D (signal_1508), .Q (signal_1509) ) ;
    buf_clk cell_666 ( .C (clk), .D (signal_1510), .Q (signal_1511) ) ;
    buf_clk cell_668 ( .C (clk), .D (signal_1512), .Q (signal_1513) ) ;
    buf_clk cell_670 ( .C (clk), .D (signal_1514), .Q (signal_1515) ) ;
    buf_clk cell_672 ( .C (clk), .D (signal_1516), .Q (signal_1517) ) ;
    buf_clk cell_674 ( .C (clk), .D (signal_1518), .Q (signal_1519) ) ;
    buf_clk cell_676 ( .C (clk), .D (signal_1520), .Q (signal_1521) ) ;
    buf_clk cell_678 ( .C (clk), .D (signal_1522), .Q (signal_1523) ) ;
    buf_clk cell_680 ( .C (clk), .D (signal_1524), .Q (signal_1525) ) ;
    buf_clk cell_682 ( .C (clk), .D (signal_1526), .Q (signal_1527) ) ;
    buf_clk cell_684 ( .C (clk), .D (signal_1528), .Q (signal_1529) ) ;
    buf_clk cell_686 ( .C (clk), .D (signal_1530), .Q (signal_1531) ) ;
    buf_clk cell_688 ( .C (clk), .D (signal_1532), .Q (signal_1533) ) ;
    buf_clk cell_690 ( .C (clk), .D (signal_1534), .Q (signal_1535) ) ;
    buf_clk cell_696 ( .C (clk), .D (signal_1540), .Q (signal_1541) ) ;
    buf_clk cell_704 ( .C (clk), .D (signal_1548), .Q (signal_1549) ) ;
    buf_clk cell_736 ( .C (clk), .D (signal_1580), .Q (signal_1581) ) ;
    buf_clk cell_746 ( .C (clk), .D (signal_1590), .Q (signal_1591) ) ;
    buf_clk cell_756 ( .C (clk), .D (signal_1600), .Q (signal_1601) ) ;
    buf_clk cell_768 ( .C (clk), .D (signal_1612), .Q (signal_1613) ) ;
    buf_clk cell_780 ( .C (clk), .D (signal_1624), .Q (signal_1625) ) ;
    buf_clk cell_794 ( .C (clk), .D (signal_1638), .Q (signal_1639) ) ;

    /* cells in depth 7 */
    buf_clk cell_697 ( .C (clk), .D (signal_1541), .Q (signal_1542) ) ;
    buf_clk cell_705 ( .C (clk), .D (signal_1549), .Q (signal_1550) ) ;
    buf_clk cell_707 ( .C (clk), .D (signal_282), .Q (signal_1552) ) ;
    buf_clk cell_709 ( .C (clk), .D (signal_689), .Q (signal_1554) ) ;
    buf_clk cell_711 ( .C (clk), .D (signal_274), .Q (signal_1556) ) ;
    buf_clk cell_713 ( .C (clk), .D (signal_681), .Q (signal_1558) ) ;
    buf_clk cell_715 ( .C (clk), .D (signal_306), .Q (signal_1560) ) ;
    buf_clk cell_717 ( .C (clk), .D (signal_713), .Q (signal_1562) ) ;
    buf_clk cell_719 ( .C (clk), .D (signal_299), .Q (signal_1564) ) ;
    buf_clk cell_721 ( .C (clk), .D (signal_706), .Q (signal_1566) ) ;
    buf_clk cell_723 ( .C (clk), .D (signal_244), .Q (signal_1568) ) ;
    buf_clk cell_725 ( .C (clk), .D (signal_651), .Q (signal_1570) ) ;
    buf_clk cell_727 ( .C (clk), .D (signal_302), .Q (signal_1572) ) ;
    buf_clk cell_729 ( .C (clk), .D (signal_709), .Q (signal_1574) ) ;
    buf_clk cell_737 ( .C (clk), .D (signal_1581), .Q (signal_1582) ) ;
    buf_clk cell_747 ( .C (clk), .D (signal_1591), .Q (signal_1592) ) ;
    buf_clk cell_757 ( .C (clk), .D (signal_1601), .Q (signal_1602) ) ;
    buf_clk cell_769 ( .C (clk), .D (signal_1613), .Q (signal_1614) ) ;
    buf_clk cell_781 ( .C (clk), .D (signal_1625), .Q (signal_1626) ) ;
    buf_clk cell_795 ( .C (clk), .D (signal_1639), .Q (signal_1640) ) ;

    /* cells in depth 8 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_305 ( .s ({signal_1435, signal_1433}), .b ({signal_1439, signal_1437}), .a ({signal_635, signal_229}), .clk (clk), .r (Fresh[169]), .c ({signal_727, signal_320}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_306 ( .s ({signal_1435, signal_1433}), .b ({signal_724, signal_317}), .a ({signal_641, signal_235}), .clk (clk), .r (Fresh[170]), .c ({signal_728, signal_321}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_307 ( .s ({signal_1435, signal_1433}), .b ({signal_711, signal_304}), .a ({signal_698, signal_291}), .clk (clk), .r (Fresh[171]), .c ({signal_729, signal_322}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_308 ( .s ({signal_1435, signal_1433}), .b ({signal_718, signal_311}), .a ({signal_1443, signal_1441}), .clk (clk), .r (Fresh[172]), .c ({signal_730, signal_323}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_309 ( .s ({signal_1435, signal_1433}), .b ({signal_619, signal_213}), .a ({signal_660, signal_253}), .clk (clk), .r (Fresh[173]), .c ({signal_731, signal_324}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_310 ( .s ({signal_1435, signal_1433}), .b ({signal_652, signal_245}), .a ({signal_704, signal_297}), .clk (clk), .r (Fresh[174]), .c ({signal_732, signal_325}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_311 ( .s ({signal_1435, signal_1433}), .b ({1'b0, 1'b1}), .a ({signal_592, signal_186}), .clk (clk), .r (Fresh[175]), .c ({signal_733, signal_326}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_312 ( .s ({signal_1435, signal_1433}), .b ({signal_1447, signal_1445}), .a ({signal_673, signal_266}), .clk (clk), .r (Fresh[176]), .c ({signal_734, signal_327}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_313 ( .s ({signal_1435, signal_1433}), .b ({signal_605, signal_199}), .a ({signal_632, signal_226}), .clk (clk), .r (Fresh[177]), .c ({signal_735, signal_328}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_314 ( .s ({signal_1435, signal_1433}), .b ({signal_666, signal_259}), .a ({signal_695, signal_288}), .clk (clk), .r (Fresh[178]), .c ({signal_736, signal_329}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_315 ( .s ({signal_1435, signal_1433}), .b ({signal_697, signal_290}), .a ({signal_670, signal_263}), .clk (clk), .r (Fresh[179]), .c ({signal_737, signal_330}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_316 ( .s ({signal_1435, signal_1433}), .b ({signal_699, signal_292}), .a ({signal_724, signal_317}), .clk (clk), .r (Fresh[180]), .c ({signal_738, signal_331}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_317 ( .s ({signal_1435, signal_1433}), .b ({signal_621, signal_215}), .a ({signal_1451, signal_1449}), .clk (clk), .r (Fresh[181]), .c ({signal_739, signal_332}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_318 ( .s ({signal_1435, signal_1433}), .b ({signal_628, signal_222}), .a ({signal_665, signal_258}), .clk (clk), .r (Fresh[182]), .c ({signal_740, signal_333}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_319 ( .s ({signal_1435, signal_1433}), .b ({signal_611, signal_205}), .a ({signal_1455, signal_1453}), .clk (clk), .r (Fresh[183]), .c ({signal_741, signal_334}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_320 ( .s ({signal_1435, signal_1433}), .b ({signal_644, signal_238}), .a ({signal_640, signal_234}), .clk (clk), .r (Fresh[184]), .c ({signal_742, signal_335}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_321 ( .s ({signal_1435, signal_1433}), .b ({signal_625, signal_219}), .a ({signal_619, signal_213}), .clk (clk), .r (Fresh[185]), .c ({signal_743, signal_336}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_322 ( .s ({signal_1435, signal_1433}), .b ({signal_722, signal_315}), .a ({signal_688, signal_281}), .clk (clk), .r (Fresh[186]), .c ({signal_744, signal_337}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_323 ( .s ({signal_1435, signal_1433}), .b ({signal_700, signal_293}), .a ({signal_608, signal_202}), .clk (clk), .r (Fresh[187]), .c ({signal_745, signal_338}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_324 ( .s ({signal_1435, signal_1433}), .b ({signal_720, signal_313}), .a ({signal_1459, signal_1457}), .clk (clk), .r (Fresh[188]), .c ({signal_746, signal_339}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_325 ( .s ({signal_1435, signal_1433}), .b ({signal_626, signal_220}), .a ({signal_635, signal_229}), .clk (clk), .r (Fresh[189]), .c ({signal_747, signal_340}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_326 ( .s ({signal_1435, signal_1433}), .b ({signal_649, signal_243}), .a ({signal_643, signal_237}), .clk (clk), .r (Fresh[190]), .c ({signal_748, signal_341}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_327 ( .s ({signal_1435, signal_1433}), .b ({signal_648, signal_242}), .a ({signal_696, signal_289}), .clk (clk), .r (Fresh[191]), .c ({signal_749, signal_342}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_328 ( .s ({signal_1435, signal_1433}), .b ({signal_622, signal_216}), .a ({signal_723, signal_316}), .clk (clk), .r (Fresh[192]), .c ({signal_750, signal_343}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_329 ( .s ({signal_1435, signal_1433}), .b ({signal_643, signal_237}), .a ({signal_690, signal_283}), .clk (clk), .r (Fresh[193]), .c ({signal_751, signal_344}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_330 ( .s ({signal_1435, signal_1433}), .b ({signal_726, signal_319}), .a ({signal_656, signal_249}), .clk (clk), .r (Fresh[194]), .c ({signal_752, signal_345}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_331 ( .s ({signal_1435, signal_1433}), .b ({signal_662, signal_255}), .a ({signal_649, signal_243}), .clk (clk), .r (Fresh[195]), .c ({signal_753, signal_346}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_332 ( .s ({signal_1435, signal_1433}), .b ({signal_613, signal_207}), .a ({signal_1463, signal_1461}), .clk (clk), .r (Fresh[196]), .c ({signal_754, signal_347}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_333 ( .s ({signal_1435, signal_1433}), .b ({signal_677, signal_270}), .a ({signal_661, signal_254}), .clk (clk), .r (Fresh[197]), .c ({signal_755, signal_348}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_334 ( .s ({signal_1435, signal_1433}), .b ({signal_668, signal_261}), .a ({signal_722, signal_315}), .clk (clk), .r (Fresh[198]), .c ({signal_756, signal_349}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_335 ( .s ({signal_1435, signal_1433}), .b ({signal_1443, signal_1441}), .a ({signal_656, signal_249}), .clk (clk), .r (Fresh[199]), .c ({signal_757, signal_350}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_336 ( .s ({signal_1435, signal_1433}), .b ({signal_662, signal_255}), .a ({signal_687, signal_280}), .clk (clk), .r (Fresh[200]), .c ({signal_758, signal_351}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_337 ( .s ({signal_1435, signal_1433}), .b ({signal_638, signal_232}), .a ({signal_597, signal_191}), .clk (clk), .r (Fresh[201]), .c ({signal_759, signal_352}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_338 ( .s ({signal_1435, signal_1433}), .b ({signal_717, signal_310}), .a ({signal_699, signal_292}), .clk (clk), .r (Fresh[202]), .c ({signal_760, signal_353}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_339 ( .s ({signal_1435, signal_1433}), .b ({signal_655, signal_248}), .a ({signal_637, signal_231}), .clk (clk), .r (Fresh[203]), .c ({signal_761, signal_354}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_340 ( .s ({signal_1435, signal_1433}), .b ({signal_707, signal_300}), .a ({signal_716, signal_309}), .clk (clk), .r (Fresh[204]), .c ({signal_762, signal_355}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_341 ( .s ({signal_1435, signal_1433}), .b ({signal_629, signal_223}), .a ({signal_692, signal_285}), .clk (clk), .r (Fresh[205]), .c ({signal_763, signal_356}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_342 ( .s ({signal_1435, signal_1433}), .b ({signal_644, signal_238}), .a ({signal_657, signal_250}), .clk (clk), .r (Fresh[206]), .c ({signal_764, signal_357}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_343 ( .s ({signal_1435, signal_1433}), .b ({signal_642, signal_236}), .a ({signal_1467, signal_1465}), .clk (clk), .r (Fresh[207]), .c ({signal_765, signal_358}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_344 ( .s ({signal_1435, signal_1433}), .b ({signal_679, signal_272}), .a ({signal_638, signal_232}), .clk (clk), .r (Fresh[208]), .c ({signal_766, signal_359}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_345 ( .s ({signal_1435, signal_1433}), .b ({signal_1471, signal_1469}), .a ({signal_711, signal_304}), .clk (clk), .r (Fresh[209]), .c ({signal_767, signal_360}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_346 ( .s ({signal_1435, signal_1433}), .b ({signal_688, signal_281}), .a ({signal_692, signal_285}), .clk (clk), .r (Fresh[210]), .c ({signal_768, signal_361}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_347 ( .s ({signal_1435, signal_1433}), .b ({signal_598, signal_192}), .a ({signal_656, signal_249}), .clk (clk), .r (Fresh[211]), .c ({signal_769, signal_362}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_348 ( .s ({signal_1435, signal_1433}), .b ({signal_705, signal_298}), .a ({signal_1475, signal_1473}), .clk (clk), .r (Fresh[212]), .c ({signal_770, signal_363}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_349 ( .s ({signal_1435, signal_1433}), .b ({signal_631, signal_225}), .a ({signal_1479, signal_1477}), .clk (clk), .r (Fresh[213]), .c ({signal_771, signal_364}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_350 ( .s ({signal_1435, signal_1433}), .b ({signal_1463, signal_1461}), .a ({signal_694, signal_287}), .clk (clk), .r (Fresh[214]), .c ({signal_772, signal_365}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_351 ( .s ({signal_1435, signal_1433}), .b ({signal_630, signal_224}), .a ({signal_1483, signal_1481}), .clk (clk), .r (Fresh[215]), .c ({signal_773, signal_366}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_352 ( .s ({signal_1435, signal_1433}), .b ({signal_596, signal_190}), .a ({signal_1487, signal_1485}), .clk (clk), .r (Fresh[216]), .c ({signal_774, signal_367}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_353 ( .s ({signal_1435, signal_1433}), .b ({signal_664, signal_257}), .a ({signal_603, signal_197}), .clk (clk), .r (Fresh[217]), .c ({signal_775, signal_368}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_354 ( .s ({signal_1435, signal_1433}), .b ({signal_1491, signal_1489}), .a ({signal_671, signal_264}), .clk (clk), .r (Fresh[218]), .c ({signal_776, signal_369}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_355 ( .s ({signal_1435, signal_1433}), .b ({signal_669, signal_262}), .a ({signal_1495, signal_1493}), .clk (clk), .r (Fresh[219]), .c ({signal_777, signal_370}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_356 ( .s ({signal_1435, signal_1433}), .b ({signal_595, signal_189}), .a ({signal_715, signal_308}), .clk (clk), .r (Fresh[220]), .c ({signal_778, signal_371}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_357 ( .s ({signal_1435, signal_1433}), .b ({signal_1439, signal_1437}), .a ({signal_657, signal_250}), .clk (clk), .r (Fresh[221]), .c ({signal_779, signal_372}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_358 ( .s ({signal_1435, signal_1433}), .b ({signal_672, signal_265}), .a ({signal_670, signal_263}), .clk (clk), .r (Fresh[222]), .c ({signal_780, signal_373}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_359 ( .s ({signal_1435, signal_1433}), .b ({signal_685, signal_278}), .a ({signal_645, signal_239}), .clk (clk), .r (Fresh[223]), .c ({signal_781, signal_374}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_360 ( .s ({signal_1435, signal_1433}), .b ({signal_593, signal_187}), .a ({signal_620, signal_214}), .clk (clk), .r (Fresh[224]), .c ({signal_782, signal_375}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_361 ( .s ({signal_1435, signal_1433}), .b ({signal_596, signal_190}), .a ({signal_602, signal_196}), .clk (clk), .r (Fresh[225]), .c ({signal_783, signal_376}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_362 ( .s ({signal_1435, signal_1433}), .b ({signal_690, signal_283}), .a ({signal_1499, signal_1497}), .clk (clk), .r (Fresh[226]), .c ({signal_784, signal_377}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_363 ( .s ({signal_1435, signal_1433}), .b ({signal_668, signal_261}), .a ({signal_702, signal_295}), .clk (clk), .r (Fresh[227]), .c ({signal_785, signal_378}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_364 ( .s ({signal_1435, signal_1433}), .b ({signal_624, signal_218}), .a ({signal_594, signal_188}), .clk (clk), .r (Fresh[228]), .c ({signal_786, signal_379}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_365 ( .s ({signal_1435, signal_1433}), .b ({signal_691, signal_284}), .a ({signal_607, signal_201}), .clk (clk), .r (Fresh[229]), .c ({signal_787, signal_380}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_366 ( .s ({signal_1435, signal_1433}), .b ({signal_1503, signal_1501}), .a ({signal_680, signal_273}), .clk (clk), .r (Fresh[230]), .c ({signal_788, signal_381}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_367 ( .s ({signal_1435, signal_1433}), .b ({signal_1503, signal_1501}), .a ({signal_603, signal_197}), .clk (clk), .r (Fresh[231]), .c ({signal_789, signal_382}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_368 ( .s ({signal_1435, signal_1433}), .b ({signal_606, signal_200}), .a ({signal_1507, signal_1505}), .clk (clk), .r (Fresh[232]), .c ({signal_790, signal_383}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_369 ( .s ({signal_1435, signal_1433}), .b ({signal_710, signal_303}), .a ({signal_676, signal_269}), .clk (clk), .r (Fresh[233]), .c ({signal_791, signal_384}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_370 ( .s ({signal_1435, signal_1433}), .b ({signal_655, signal_248}), .a ({signal_663, signal_256}), .clk (clk), .r (Fresh[234]), .c ({signal_792, signal_385}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_371 ( .s ({signal_1435, signal_1433}), .b ({signal_1499, signal_1497}), .a ({signal_668, signal_261}), .clk (clk), .r (Fresh[235]), .c ({signal_793, signal_386}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_372 ( .s ({signal_1435, signal_1433}), .b ({signal_641, signal_235}), .a ({signal_712, signal_305}), .clk (clk), .r (Fresh[236]), .c ({signal_794, signal_387}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_373 ( .s ({signal_1435, signal_1433}), .b ({signal_631, signal_225}), .a ({signal_1483, signal_1481}), .clk (clk), .r (Fresh[237]), .c ({signal_795, signal_388}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_374 ( .s ({signal_1435, signal_1433}), .b ({signal_621, signal_215}), .a ({signal_1499, signal_1497}), .clk (clk), .r (Fresh[238]), .c ({signal_796, signal_389}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_375 ( .s ({signal_1435, signal_1433}), .b ({signal_654, signal_247}), .a ({signal_683, signal_276}), .clk (clk), .r (Fresh[239]), .c ({signal_797, signal_390}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_376 ( .s ({signal_1435, signal_1433}), .b ({signal_623, signal_217}), .a ({signal_625, signal_219}), .clk (clk), .r (Fresh[240]), .c ({signal_798, signal_391}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_377 ( .s ({signal_1435, signal_1433}), .b ({signal_627, signal_221}), .a ({signal_618, signal_212}), .clk (clk), .r (Fresh[241]), .c ({signal_799, signal_392}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_378 ( .s ({signal_1435, signal_1433}), .b ({signal_1511, signal_1509}), .a ({signal_659, signal_252}), .clk (clk), .r (Fresh[242]), .c ({signal_800, signal_393}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_379 ( .s ({signal_1435, signal_1433}), .b ({signal_597, signal_191}), .a ({signal_609, signal_203}), .clk (clk), .r (Fresh[243]), .c ({signal_801, signal_394}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_380 ( .s ({signal_1435, signal_1433}), .b ({signal_704, signal_297}), .a ({signal_642, signal_236}), .clk (clk), .r (Fresh[244]), .c ({signal_802, signal_395}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_381 ( .s ({signal_1435, signal_1433}), .b ({signal_620, signal_214}), .a ({signal_1443, signal_1441}), .clk (clk), .r (Fresh[245]), .c ({signal_803, signal_396}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_382 ( .s ({signal_1435, signal_1433}), .b ({signal_661, signal_254}), .a ({signal_595, signal_189}), .clk (clk), .r (Fresh[246]), .c ({signal_804, signal_397}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_383 ( .s ({signal_1435, signal_1433}), .b ({signal_661, signal_254}), .a ({signal_625, signal_219}), .clk (clk), .r (Fresh[247]), .c ({signal_805, signal_398}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_384 ( .s ({signal_1435, signal_1433}), .b ({signal_616, signal_210}), .a ({signal_598, signal_192}), .clk (clk), .r (Fresh[248]), .c ({signal_806, signal_399}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_385 ( .s ({signal_1435, signal_1433}), .b ({signal_685, signal_278}), .a ({signal_674, signal_267}), .clk (clk), .r (Fresh[249]), .c ({signal_807, signal_400}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_386 ( .s ({signal_1435, signal_1433}), .b ({signal_618, signal_212}), .a ({signal_621, signal_215}), .clk (clk), .r (Fresh[250]), .c ({signal_808, signal_401}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_387 ( .s ({signal_1435, signal_1433}), .b ({signal_703, signal_296}), .a ({signal_678, signal_271}), .clk (clk), .r (Fresh[251]), .c ({signal_809, signal_402}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_388 ( .s ({signal_1435, signal_1433}), .b ({signal_1515, signal_1513}), .a ({signal_599, signal_193}), .clk (clk), .r (Fresh[252]), .c ({signal_810, signal_403}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_389 ( .s ({signal_1435, signal_1433}), .b ({signal_615, signal_209}), .a ({signal_686, signal_279}), .clk (clk), .r (Fresh[253]), .c ({signal_811, signal_404}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_390 ( .s ({signal_1435, signal_1433}), .b ({signal_658, signal_251}), .a ({signal_704, signal_297}), .clk (clk), .r (Fresh[254]), .c ({signal_812, signal_405}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_391 ( .s ({signal_1435, signal_1433}), .b ({signal_609, signal_203}), .a ({signal_1519, signal_1517}), .clk (clk), .r (Fresh[255]), .c ({signal_813, signal_406}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_392 ( .s ({signal_1435, signal_1433}), .b ({signal_649, signal_243}), .a ({signal_693, signal_286}), .clk (clk), .r (Fresh[256]), .c ({signal_814, signal_407}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_393 ( .s ({signal_1435, signal_1433}), .b ({signal_640, signal_234}), .a ({signal_1523, signal_1521}), .clk (clk), .r (Fresh[257]), .c ({signal_815, signal_408}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_394 ( .s ({signal_1435, signal_1433}), .b ({signal_701, signal_294}), .a ({signal_662, signal_255}), .clk (clk), .r (Fresh[258]), .c ({signal_816, signal_409}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_395 ( .s ({signal_1435, signal_1433}), .b ({signal_640, signal_234}), .a ({signal_675, signal_268}), .clk (clk), .r (Fresh[259]), .c ({signal_817, signal_410}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_396 ( .s ({signal_1435, signal_1433}), .b ({signal_647, signal_241}), .a ({signal_1499, signal_1497}), .clk (clk), .r (Fresh[260]), .c ({signal_818, signal_411}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_397 ( .s ({signal_1435, signal_1433}), .b ({signal_597, signal_191}), .a ({signal_639, signal_233}), .clk (clk), .r (Fresh[261]), .c ({signal_819, signal_412}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_398 ( .s ({signal_1435, signal_1433}), .b ({signal_670, signal_263}), .a ({signal_599, signal_193}), .clk (clk), .r (Fresh[262]), .c ({signal_820, signal_413}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_399 ( .s ({signal_1435, signal_1433}), .b ({signal_723, signal_316}), .a ({signal_625, signal_219}), .clk (clk), .r (Fresh[263]), .c ({signal_821, signal_414}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_400 ( .s ({signal_1435, signal_1433}), .b ({signal_636, signal_230}), .a ({signal_719, signal_312}), .clk (clk), .r (Fresh[264]), .c ({signal_822, signal_415}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_401 ( .s ({signal_1435, signal_1433}), .b ({signal_684, signal_277}), .a ({signal_623, signal_217}), .clk (clk), .r (Fresh[265]), .c ({signal_823, signal_416}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_402 ( .s ({signal_1435, signal_1433}), .b ({signal_704, signal_297}), .a ({signal_710, signal_303}), .clk (clk), .r (Fresh[266]), .c ({signal_824, signal_417}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_403 ( .s ({signal_1435, signal_1433}), .b ({signal_708, signal_301}), .a ({signal_682, signal_275}), .clk (clk), .r (Fresh[267]), .c ({signal_825, signal_418}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_404 ( .s ({signal_1435, signal_1433}), .b ({signal_671, signal_264}), .a ({signal_610, signal_204}), .clk (clk), .r (Fresh[268]), .c ({signal_826, signal_419}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_405 ( .s ({signal_1435, signal_1433}), .b ({signal_601, signal_195}), .a ({signal_628, signal_222}), .clk (clk), .r (Fresh[269]), .c ({signal_827, signal_420}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_406 ( .s ({signal_1435, signal_1433}), .b ({signal_634, signal_228}), .a ({signal_648, signal_242}), .clk (clk), .r (Fresh[270]), .c ({signal_828, signal_421}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_407 ( .s ({signal_1435, signal_1433}), .b ({signal_659, signal_252}), .a ({signal_724, signal_317}), .clk (clk), .r (Fresh[271]), .c ({signal_829, signal_422}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_408 ( .s ({signal_1435, signal_1433}), .b ({signal_625, signal_219}), .a ({signal_593, signal_187}), .clk (clk), .r (Fresh[272]), .c ({signal_830, signal_423}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_409 ( .s ({signal_1435, signal_1433}), .b ({signal_704, signal_297}), .a ({signal_1455, signal_1453}), .clk (clk), .r (Fresh[273]), .c ({signal_831, signal_424}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_410 ( .s ({signal_1435, signal_1433}), .b ({signal_593, signal_187}), .a ({signal_1527, signal_1525}), .clk (clk), .r (Fresh[274]), .c ({signal_832, signal_425}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_411 ( .s ({signal_1435, signal_1433}), .b ({signal_596, signal_190}), .a ({signal_633, signal_227}), .clk (clk), .r (Fresh[275]), .c ({signal_833, signal_426}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_412 ( .s ({signal_1435, signal_1433}), .b ({signal_683, signal_276}), .a ({signal_1531, signal_1529}), .clk (clk), .r (Fresh[276]), .c ({signal_834, signal_427}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_413 ( .s ({signal_1435, signal_1433}), .b ({signal_648, signal_242}), .a ({signal_616, signal_210}), .clk (clk), .r (Fresh[277]), .c ({signal_835, signal_428}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_414 ( .s ({signal_1435, signal_1433}), .b ({signal_604, signal_198}), .a ({signal_613, signal_207}), .clk (clk), .r (Fresh[278]), .c ({signal_836, signal_429}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_415 ( .s ({signal_1435, signal_1433}), .b ({signal_671, signal_264}), .a ({signal_725, signal_318}), .clk (clk), .r (Fresh[279]), .c ({signal_837, signal_430}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_416 ( .s ({signal_1435, signal_1433}), .b ({signal_1527, signal_1525}), .a ({signal_679, signal_272}), .clk (clk), .r (Fresh[280]), .c ({signal_838, signal_431}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_417 ( .s ({signal_1435, signal_1433}), .b ({signal_705, signal_298}), .a ({signal_612, signal_206}), .clk (clk), .r (Fresh[281]), .c ({signal_839, signal_432}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_418 ( .s ({signal_1435, signal_1433}), .b ({signal_646, signal_240}), .a ({signal_591, signal_185}), .clk (clk), .r (Fresh[282]), .c ({signal_840, signal_433}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_419 ( .s ({signal_1435, signal_1433}), .b ({signal_697, signal_290}), .a ({signal_646, signal_240}), .clk (clk), .r (Fresh[283]), .c ({signal_841, signal_434}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_420 ( .s ({signal_1435, signal_1433}), .b ({signal_721, signal_314}), .a ({signal_619, signal_213}), .clk (clk), .r (Fresh[284]), .c ({signal_842, signal_435}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_421 ( .s ({signal_1435, signal_1433}), .b ({signal_667, signal_260}), .a ({signal_623, signal_217}), .clk (clk), .r (Fresh[285]), .c ({signal_843, signal_436}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_422 ( .s ({signal_1435, signal_1433}), .b ({signal_600, signal_194}), .a ({signal_645, signal_239}), .clk (clk), .r (Fresh[286]), .c ({signal_844, signal_437}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_423 ( .s ({signal_1435, signal_1433}), .b ({signal_617, signal_211}), .a ({signal_614, signal_208}), .clk (clk), .r (Fresh[287]), .c ({signal_845, signal_438}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_424 ( .s ({signal_1435, signal_1433}), .b ({signal_664, signal_257}), .a ({signal_616, signal_210}), .clk (clk), .r (Fresh[288]), .c ({signal_846, signal_439}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_425 ( .s ({signal_1435, signal_1433}), .b ({signal_1535, signal_1533}), .a ({signal_702, signal_295}), .clk (clk), .r (Fresh[289]), .c ({signal_847, signal_440}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_426 ( .s ({signal_1435, signal_1433}), .b ({signal_714, signal_307}), .a ({signal_653, signal_246}), .clk (clk), .r (Fresh[290]), .c ({signal_848, signal_441}) ) ;
    buf_clk cell_698 ( .C (clk), .D (signal_1542), .Q (signal_1543) ) ;
    buf_clk cell_706 ( .C (clk), .D (signal_1550), .Q (signal_1551) ) ;
    buf_clk cell_708 ( .C (clk), .D (signal_1552), .Q (signal_1553) ) ;
    buf_clk cell_710 ( .C (clk), .D (signal_1554), .Q (signal_1555) ) ;
    buf_clk cell_712 ( .C (clk), .D (signal_1556), .Q (signal_1557) ) ;
    buf_clk cell_714 ( .C (clk), .D (signal_1558), .Q (signal_1559) ) ;
    buf_clk cell_716 ( .C (clk), .D (signal_1560), .Q (signal_1561) ) ;
    buf_clk cell_718 ( .C (clk), .D (signal_1562), .Q (signal_1563) ) ;
    buf_clk cell_720 ( .C (clk), .D (signal_1564), .Q (signal_1565) ) ;
    buf_clk cell_722 ( .C (clk), .D (signal_1566), .Q (signal_1567) ) ;
    buf_clk cell_724 ( .C (clk), .D (signal_1568), .Q (signal_1569) ) ;
    buf_clk cell_726 ( .C (clk), .D (signal_1570), .Q (signal_1571) ) ;
    buf_clk cell_728 ( .C (clk), .D (signal_1572), .Q (signal_1573) ) ;
    buf_clk cell_730 ( .C (clk), .D (signal_1574), .Q (signal_1575) ) ;
    buf_clk cell_738 ( .C (clk), .D (signal_1582), .Q (signal_1583) ) ;
    buf_clk cell_748 ( .C (clk), .D (signal_1592), .Q (signal_1593) ) ;
    buf_clk cell_758 ( .C (clk), .D (signal_1602), .Q (signal_1603) ) ;
    buf_clk cell_770 ( .C (clk), .D (signal_1614), .Q (signal_1615) ) ;
    buf_clk cell_782 ( .C (clk), .D (signal_1626), .Q (signal_1627) ) ;
    buf_clk cell_796 ( .C (clk), .D (signal_1640), .Q (signal_1641) ) ;

    /* cells in depth 9 */
    buf_clk cell_739 ( .C (clk), .D (signal_1583), .Q (signal_1584) ) ;
    buf_clk cell_749 ( .C (clk), .D (signal_1593), .Q (signal_1594) ) ;
    buf_clk cell_759 ( .C (clk), .D (signal_1603), .Q (signal_1604) ) ;
    buf_clk cell_771 ( .C (clk), .D (signal_1615), .Q (signal_1616) ) ;
    buf_clk cell_783 ( .C (clk), .D (signal_1627), .Q (signal_1628) ) ;
    buf_clk cell_797 ( .C (clk), .D (signal_1641), .Q (signal_1642) ) ;

    /* cells in depth 10 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_427 ( .s ({signal_1551, signal_1543}), .b ({signal_753, signal_346}), .a ({signal_800, signal_393}), .clk (clk), .r (Fresh[291]), .c ({signal_850, signal_442}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_428 ( .s ({signal_1551, signal_1543}), .b ({signal_751, signal_344}), .a ({signal_833, signal_426}), .clk (clk), .r (Fresh[292]), .c ({signal_851, signal_443}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_429 ( .s ({signal_1551, signal_1543}), .b ({signal_796, signal_389}), .a ({signal_812, signal_405}), .clk (clk), .r (Fresh[293]), .c ({signal_852, signal_444}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_430 ( .s ({signal_1551, signal_1543}), .b ({signal_771, signal_364}), .a ({signal_843, signal_436}), .clk (clk), .r (Fresh[294]), .c ({signal_853, signal_445}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_431 ( .s ({signal_1551, signal_1543}), .b ({signal_840, signal_433}), .a ({signal_831, signal_424}), .clk (clk), .r (Fresh[295]), .c ({signal_854, signal_446}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_432 ( .s ({signal_1551, signal_1543}), .b ({signal_744, signal_337}), .a ({signal_790, signal_383}), .clk (clk), .r (Fresh[296]), .c ({signal_855, signal_447}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_433 ( .s ({signal_1551, signal_1543}), .b ({signal_774, signal_367}), .a ({signal_829, signal_422}), .clk (clk), .r (Fresh[297]), .c ({signal_856, signal_448}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_434 ( .s ({signal_1551, signal_1543}), .b ({signal_750, signal_343}), .a ({signal_809, signal_402}), .clk (clk), .r (Fresh[298]), .c ({signal_857, signal_449}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_435 ( .s ({signal_1551, signal_1543}), .b ({signal_847, signal_440}), .a ({signal_731, signal_324}), .clk (clk), .r (Fresh[299]), .c ({signal_858, signal_450}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_436 ( .s ({signal_1551, signal_1543}), .b ({signal_766, signal_359}), .a ({signal_848, signal_441}), .clk (clk), .r (Fresh[300]), .c ({signal_859, signal_451}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_437 ( .s ({signal_1551, signal_1543}), .b ({signal_764, signal_357}), .a ({signal_789, signal_382}), .clk (clk), .r (Fresh[301]), .c ({signal_860, signal_452}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_438 ( .s ({signal_1551, signal_1543}), .b ({signal_799, signal_392}), .a ({signal_793, signal_386}), .clk (clk), .r (Fresh[302]), .c ({signal_861, signal_453}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_439 ( .s ({signal_1551, signal_1543}), .b ({signal_738, signal_331}), .a ({signal_827, signal_420}), .clk (clk), .r (Fresh[303]), .c ({signal_862, signal_454}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_440 ( .s ({signal_1551, signal_1543}), .b ({signal_822, signal_415}), .a ({signal_823, signal_416}), .clk (clk), .r (Fresh[304]), .c ({signal_863, signal_455}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_441 ( .s ({signal_1551, signal_1543}), .b ({signal_803, signal_396}), .a ({signal_1555, signal_1553}), .clk (clk), .r (Fresh[305]), .c ({signal_864, signal_456}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_442 ( .s ({signal_1551, signal_1543}), .b ({signal_842, signal_435}), .a ({signal_826, signal_419}), .clk (clk), .r (Fresh[306]), .c ({signal_865, signal_457}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_443 ( .s ({signal_1551, signal_1543}), .b ({signal_730, signal_323}), .a ({signal_755, signal_348}), .clk (clk), .r (Fresh[307]), .c ({signal_866, signal_458}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_444 ( .s ({signal_1551, signal_1543}), .b ({signal_806, signal_399}), .a ({signal_1559, signal_1557}), .clk (clk), .r (Fresh[308]), .c ({signal_867, signal_459}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_445 ( .s ({signal_1551, signal_1543}), .b ({signal_839, signal_432}), .a ({signal_1563, signal_1561}), .clk (clk), .r (Fresh[309]), .c ({signal_868, signal_460}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_446 ( .s ({signal_1551, signal_1543}), .b ({signal_786, signal_379}), .a ({signal_733, signal_326}), .clk (clk), .r (Fresh[310]), .c ({signal_869, signal_461}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_447 ( .s ({signal_1551, signal_1543}), .b ({signal_775, signal_368}), .a ({signal_758, signal_351}), .clk (clk), .r (Fresh[311]), .c ({signal_870, signal_462}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_448 ( .s ({signal_1551, signal_1543}), .b ({signal_741, signal_334}), .a ({signal_781, signal_374}), .clk (clk), .r (Fresh[312]), .c ({signal_871, signal_463}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_449 ( .s ({signal_1551, signal_1543}), .b ({signal_819, signal_412}), .a ({signal_732, signal_325}), .clk (clk), .r (Fresh[313]), .c ({signal_872, signal_464}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_450 ( .s ({signal_1551, signal_1543}), .b ({signal_768, signal_361}), .a ({signal_808, signal_401}), .clk (clk), .r (Fresh[314]), .c ({signal_873, signal_465}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_451 ( .s ({signal_1551, signal_1543}), .b ({signal_734, signal_327}), .a ({signal_737, signal_330}), .clk (clk), .r (Fresh[315]), .c ({signal_874, signal_466}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_452 ( .s ({signal_1551, signal_1543}), .b ({signal_727, signal_320}), .a ({signal_752, signal_345}), .clk (clk), .r (Fresh[316]), .c ({signal_875, signal_467}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_453 ( .s ({signal_1551, signal_1543}), .b ({signal_815, signal_408}), .a ({signal_845, signal_438}), .clk (clk), .r (Fresh[317]), .c ({signal_876, signal_468}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_454 ( .s ({signal_1551, signal_1543}), .b ({signal_837, signal_430}), .a ({signal_824, signal_417}), .clk (clk), .r (Fresh[318]), .c ({signal_877, signal_469}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_455 ( .s ({signal_1551, signal_1543}), .b ({signal_821, signal_414}), .a ({signal_747, signal_340}), .clk (clk), .r (Fresh[319]), .c ({signal_878, signal_470}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_456 ( .s ({signal_1551, signal_1543}), .b ({signal_778, signal_371}), .a ({signal_1567, signal_1565}), .clk (clk), .r (Fresh[320]), .c ({signal_879, signal_471}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_457 ( .s ({signal_1551, signal_1543}), .b ({signal_756, signal_349}), .a ({signal_757, signal_350}), .clk (clk), .r (Fresh[321]), .c ({signal_880, signal_472}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_458 ( .s ({signal_1551, signal_1543}), .b ({signal_791, signal_384}), .a ({signal_794, signal_387}), .clk (clk), .r (Fresh[322]), .c ({signal_881, signal_473}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_459 ( .s ({signal_1551, signal_1543}), .b ({signal_782, signal_375}), .a ({signal_748, signal_341}), .clk (clk), .r (Fresh[323]), .c ({signal_882, signal_474}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_460 ( .s ({signal_1551, signal_1543}), .b ({signal_795, signal_388}), .a ({signal_817, signal_410}), .clk (clk), .r (Fresh[324]), .c ({signal_883, signal_475}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_461 ( .s ({signal_1551, signal_1543}), .b ({signal_767, signal_360}), .a ({signal_792, signal_385}), .clk (clk), .r (Fresh[325]), .c ({signal_884, signal_476}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_462 ( .s ({signal_1551, signal_1543}), .b ({signal_844, signal_437}), .a ({signal_746, signal_339}), .clk (clk), .r (Fresh[326]), .c ({signal_885, signal_477}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_463 ( .s ({signal_1551, signal_1543}), .b ({signal_810, signal_403}), .a ({signal_739, signal_332}), .clk (clk), .r (Fresh[327]), .c ({signal_886, signal_478}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_464 ( .s ({signal_1551, signal_1543}), .b ({signal_742, signal_335}), .a ({signal_749, signal_342}), .clk (clk), .r (Fresh[328]), .c ({signal_887, signal_479}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_465 ( .s ({signal_1551, signal_1543}), .b ({signal_743, signal_336}), .a ({signal_772, signal_365}), .clk (clk), .r (Fresh[329]), .c ({signal_888, signal_480}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_466 ( .s ({signal_1551, signal_1543}), .b ({signal_763, signal_356}), .a ({signal_835, signal_428}), .clk (clk), .r (Fresh[330]), .c ({signal_889, signal_481}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_467 ( .s ({signal_1551, signal_1543}), .b ({signal_776, signal_369}), .a ({signal_785, signal_378}), .clk (clk), .r (Fresh[331]), .c ({signal_890, signal_482}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_468 ( .s ({signal_1551, signal_1543}), .b ({signal_798, signal_391}), .a ({signal_804, signal_397}), .clk (clk), .r (Fresh[332]), .c ({signal_891, signal_483}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_469 ( .s ({signal_1551, signal_1543}), .b ({signal_780, signal_373}), .a ({signal_735, signal_328}), .clk (clk), .r (Fresh[333]), .c ({signal_892, signal_484}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_470 ( .s ({signal_1551, signal_1543}), .b ({signal_828, signal_421}), .a ({signal_783, signal_376}), .clk (clk), .r (Fresh[334]), .c ({signal_893, signal_485}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_471 ( .s ({signal_1551, signal_1543}), .b ({signal_759, signal_352}), .a ({signal_773, signal_366}), .clk (clk), .r (Fresh[335]), .c ({signal_894, signal_486}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_472 ( .s ({signal_1551, signal_1543}), .b ({signal_838, signal_431}), .a ({signal_825, signal_418}), .clk (clk), .r (Fresh[336]), .c ({signal_895, signal_487}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_473 ( .s ({signal_1551, signal_1543}), .b ({signal_805, signal_398}), .a ({signal_832, signal_425}), .clk (clk), .r (Fresh[337]), .c ({signal_896, signal_488}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_474 ( .s ({signal_1551, signal_1543}), .b ({signal_761, signal_354}), .a ({signal_818, signal_411}), .clk (clk), .r (Fresh[338]), .c ({signal_897, signal_489}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_475 ( .s ({signal_1551, signal_1543}), .b ({signal_760, signal_353}), .a ({signal_740, signal_333}), .clk (clk), .r (Fresh[339]), .c ({signal_898, signal_490}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_476 ( .s ({signal_1551, signal_1543}), .b ({signal_769, signal_362}), .a ({signal_788, signal_381}), .clk (clk), .r (Fresh[340]), .c ({signal_899, signal_491}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_477 ( .s ({signal_1551, signal_1543}), .b ({signal_787, signal_380}), .a ({signal_811, signal_404}), .clk (clk), .r (Fresh[341]), .c ({signal_900, signal_492}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_478 ( .s ({signal_1551, signal_1543}), .b ({signal_1571, signal_1569}), .a ({signal_770, signal_363}), .clk (clk), .r (Fresh[342]), .c ({signal_901, signal_493}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_479 ( .s ({signal_1551, signal_1543}), .b ({signal_765, signal_358}), .a ({signal_802, signal_395}), .clk (clk), .r (Fresh[343]), .c ({signal_902, signal_494}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_480 ( .s ({signal_1551, signal_1543}), .b ({signal_846, signal_439}), .a ({signal_836, signal_429}), .clk (clk), .r (Fresh[344]), .c ({signal_903, signal_495}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_481 ( .s ({signal_1551, signal_1543}), .b ({signal_814, signal_407}), .a ({signal_729, signal_322}), .clk (clk), .r (Fresh[345]), .c ({signal_904, signal_496}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_482 ( .s ({signal_1551, signal_1543}), .b ({signal_762, signal_355}), .a ({signal_841, signal_434}), .clk (clk), .r (Fresh[346]), .c ({signal_905, signal_497}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_483 ( .s ({signal_1551, signal_1543}), .b ({signal_797, signal_390}), .a ({signal_816, signal_409}), .clk (clk), .r (Fresh[347]), .c ({signal_906, signal_498}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_484 ( .s ({signal_1551, signal_1543}), .b ({signal_736, signal_329}), .a ({signal_784, signal_377}), .clk (clk), .r (Fresh[348]), .c ({signal_907, signal_499}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_485 ( .s ({signal_1551, signal_1543}), .b ({signal_728, signal_321}), .a ({signal_830, signal_423}), .clk (clk), .r (Fresh[349]), .c ({signal_908, signal_500}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_486 ( .s ({signal_1551, signal_1543}), .b ({signal_820, signal_413}), .a ({signal_807, signal_400}), .clk (clk), .r (Fresh[350]), .c ({signal_909, signal_501}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_487 ( .s ({signal_1551, signal_1543}), .b ({signal_779, signal_372}), .a ({signal_813, signal_406}), .clk (clk), .r (Fresh[351]), .c ({signal_910, signal_502}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_488 ( .s ({signal_1551, signal_1543}), .b ({signal_1575, signal_1573}), .a ({signal_834, signal_427}), .clk (clk), .r (Fresh[352]), .c ({signal_911, signal_503}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_489 ( .s ({signal_1551, signal_1543}), .b ({signal_777, signal_370}), .a ({signal_754, signal_347}), .clk (clk), .r (Fresh[353]), .c ({signal_912, signal_504}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_490 ( .s ({signal_1551, signal_1543}), .b ({signal_801, signal_394}), .a ({signal_745, signal_338}), .clk (clk), .r (Fresh[354]), .c ({signal_913, signal_505}) ) ;
    buf_clk cell_740 ( .C (clk), .D (signal_1584), .Q (signal_1585) ) ;
    buf_clk cell_750 ( .C (clk), .D (signal_1594), .Q (signal_1595) ) ;
    buf_clk cell_760 ( .C (clk), .D (signal_1604), .Q (signal_1605) ) ;
    buf_clk cell_772 ( .C (clk), .D (signal_1616), .Q (signal_1617) ) ;
    buf_clk cell_784 ( .C (clk), .D (signal_1628), .Q (signal_1629) ) ;
    buf_clk cell_798 ( .C (clk), .D (signal_1642), .Q (signal_1643) ) ;

    /* cells in depth 11 */
    buf_clk cell_761 ( .C (clk), .D (signal_1605), .Q (signal_1606) ) ;
    buf_clk cell_773 ( .C (clk), .D (signal_1617), .Q (signal_1618) ) ;
    buf_clk cell_785 ( .C (clk), .D (signal_1629), .Q (signal_1630) ) ;
    buf_clk cell_799 ( .C (clk), .D (signal_1643), .Q (signal_1644) ) ;

    /* cells in depth 12 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_491 ( .s ({signal_1595, signal_1585}), .b ({signal_883, signal_475}), .a ({signal_852, signal_444}), .clk (clk), .r (Fresh[355]), .c ({signal_915, signal_506}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_492 ( .s ({signal_1595, signal_1585}), .b ({signal_858, signal_450}), .a ({signal_863, signal_455}), .clk (clk), .r (Fresh[356]), .c ({signal_916, signal_507}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_493 ( .s ({signal_1595, signal_1585}), .b ({signal_897, signal_489}), .a ({signal_878, signal_470}), .clk (clk), .r (Fresh[357]), .c ({signal_917, signal_508}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_494 ( .s ({signal_1595, signal_1585}), .b ({signal_891, signal_483}), .a ({signal_853, signal_445}), .clk (clk), .r (Fresh[358]), .c ({signal_918, signal_509}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_495 ( .s ({signal_1595, signal_1585}), .b ({signal_907, signal_499}), .a ({signal_865, signal_457}), .clk (clk), .r (Fresh[359]), .c ({signal_919, signal_510}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_496 ( .s ({signal_1595, signal_1585}), .b ({signal_888, signal_480}), .a ({signal_886, signal_478}), .clk (clk), .r (Fresh[360]), .c ({signal_920, signal_511}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_497 ( .s ({signal_1595, signal_1585}), .b ({signal_909, signal_501}), .a ({signal_884, signal_476}), .clk (clk), .r (Fresh[361]), .c ({signal_921, signal_512}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_498 ( .s ({signal_1595, signal_1585}), .b ({signal_898, signal_490}), .a ({signal_876, signal_468}), .clk (clk), .r (Fresh[362]), .c ({signal_922, signal_513}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_499 ( .s ({signal_1595, signal_1585}), .b ({signal_911, signal_503}), .a ({signal_869, signal_461}), .clk (clk), .r (Fresh[363]), .c ({signal_923, signal_514}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_500 ( .s ({signal_1595, signal_1585}), .b ({signal_866, signal_458}), .a ({signal_870, signal_462}), .clk (clk), .r (Fresh[364]), .c ({signal_924, signal_515}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_501 ( .s ({signal_1595, signal_1585}), .b ({signal_857, signal_449}), .a ({signal_875, signal_467}), .clk (clk), .r (Fresh[365]), .c ({signal_925, signal_516}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_502 ( .s ({signal_1595, signal_1585}), .b ({signal_906, signal_498}), .a ({signal_899, signal_491}), .clk (clk), .r (Fresh[366]), .c ({signal_926, signal_517}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_503 ( .s ({signal_1595, signal_1585}), .b ({signal_860, signal_452}), .a ({signal_896, signal_488}), .clk (clk), .r (Fresh[367]), .c ({signal_927, signal_518}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_504 ( .s ({signal_1595, signal_1585}), .b ({signal_900, signal_492}), .a ({signal_877, signal_469}), .clk (clk), .r (Fresh[368]), .c ({signal_928, signal_519}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_505 ( .s ({signal_1595, signal_1585}), .b ({signal_903, signal_495}), .a ({signal_880, signal_472}), .clk (clk), .r (Fresh[369]), .c ({signal_929, signal_520}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_506 ( .s ({signal_1595, signal_1585}), .b ({signal_904, signal_496}), .a ({signal_872, signal_464}), .clk (clk), .r (Fresh[370]), .c ({signal_930, signal_521}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_507 ( .s ({signal_1595, signal_1585}), .b ({signal_902, signal_494}), .a ({signal_868, signal_460}), .clk (clk), .r (Fresh[371]), .c ({signal_931, signal_522}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_508 ( .s ({signal_1595, signal_1585}), .b ({signal_881, signal_473}), .a ({signal_905, signal_497}), .clk (clk), .r (Fresh[372]), .c ({signal_932, signal_523}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_509 ( .s ({signal_1595, signal_1585}), .b ({signal_901, signal_493}), .a ({signal_867, signal_459}), .clk (clk), .r (Fresh[373]), .c ({signal_933, signal_524}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_510 ( .s ({signal_1595, signal_1585}), .b ({signal_862, signal_454}), .a ({signal_910, signal_502}), .clk (clk), .r (Fresh[374]), .c ({signal_934, signal_525}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_511 ( .s ({signal_1595, signal_1585}), .b ({signal_912, signal_504}), .a ({signal_887, signal_479}), .clk (clk), .r (Fresh[375]), .c ({signal_935, signal_526}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_512 ( .s ({signal_1595, signal_1585}), .b ({signal_864, signal_456}), .a ({signal_855, signal_447}), .clk (clk), .r (Fresh[376]), .c ({signal_936, signal_527}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_513 ( .s ({signal_1595, signal_1585}), .b ({signal_854, signal_446}), .a ({signal_874, signal_466}), .clk (clk), .r (Fresh[377]), .c ({signal_937, signal_528}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_514 ( .s ({signal_1595, signal_1585}), .b ({signal_879, signal_471}), .a ({signal_893, signal_485}), .clk (clk), .r (Fresh[378]), .c ({signal_938, signal_529}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_515 ( .s ({signal_1595, signal_1585}), .b ({signal_890, signal_482}), .a ({signal_859, signal_451}), .clk (clk), .r (Fresh[379]), .c ({signal_939, signal_530}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_516 ( .s ({signal_1595, signal_1585}), .b ({signal_856, signal_448}), .a ({signal_871, signal_463}), .clk (clk), .r (Fresh[380]), .c ({signal_940, signal_531}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_517 ( .s ({signal_1595, signal_1585}), .b ({signal_873, signal_465}), .a ({signal_913, signal_505}), .clk (clk), .r (Fresh[381]), .c ({signal_941, signal_532}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_518 ( .s ({signal_1595, signal_1585}), .b ({signal_861, signal_453}), .a ({signal_908, signal_500}), .clk (clk), .r (Fresh[382]), .c ({signal_942, signal_533}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_519 ( .s ({signal_1595, signal_1585}), .b ({signal_882, signal_474}), .a ({signal_889, signal_481}), .clk (clk), .r (Fresh[383]), .c ({signal_943, signal_534}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_520 ( .s ({signal_1595, signal_1585}), .b ({signal_885, signal_477}), .a ({signal_892, signal_484}), .clk (clk), .r (Fresh[384]), .c ({signal_944, signal_535}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_521 ( .s ({signal_1595, signal_1585}), .b ({signal_895, signal_487}), .a ({signal_850, signal_442}), .clk (clk), .r (Fresh[385]), .c ({signal_945, signal_536}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_522 ( .s ({signal_1595, signal_1585}), .b ({signal_894, signal_486}), .a ({signal_851, signal_443}), .clk (clk), .r (Fresh[386]), .c ({signal_946, signal_537}) ) ;
    buf_clk cell_762 ( .C (clk), .D (signal_1606), .Q (signal_1607) ) ;
    buf_clk cell_774 ( .C (clk), .D (signal_1618), .Q (signal_1619) ) ;
    buf_clk cell_786 ( .C (clk), .D (signal_1630), .Q (signal_1631) ) ;
    buf_clk cell_800 ( .C (clk), .D (signal_1644), .Q (signal_1645) ) ;

    /* cells in depth 13 */
    buf_clk cell_787 ( .C (clk), .D (signal_1631), .Q (signal_1632) ) ;
    buf_clk cell_801 ( .C (clk), .D (signal_1645), .Q (signal_1646) ) ;

    /* cells in depth 14 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_523 ( .s ({signal_1619, signal_1607}), .b ({signal_940, signal_531}), .a ({signal_927, signal_518}), .clk (clk), .r (Fresh[387]), .c ({signal_948, signal_538}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_524 ( .s ({signal_1619, signal_1607}), .b ({signal_917, signal_508}), .a ({signal_944, signal_535}), .clk (clk), .r (Fresh[388]), .c ({signal_949, signal_539}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_525 ( .s ({signal_1619, signal_1607}), .b ({signal_933, signal_524}), .a ({signal_932, signal_523}), .clk (clk), .r (Fresh[389]), .c ({signal_950, signal_540}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_526 ( .s ({signal_1619, signal_1607}), .b ({signal_928, signal_519}), .a ({signal_936, signal_527}), .clk (clk), .r (Fresh[390]), .c ({signal_951, signal_541}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_527 ( .s ({signal_1619, signal_1607}), .b ({signal_937, signal_528}), .a ({signal_915, signal_506}), .clk (clk), .r (Fresh[391]), .c ({signal_952, signal_542}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_528 ( .s ({signal_1619, signal_1607}), .b ({signal_935, signal_526}), .a ({signal_946, signal_537}), .clk (clk), .r (Fresh[392]), .c ({signal_953, signal_543}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_529 ( .s ({signal_1619, signal_1607}), .b ({signal_919, signal_510}), .a ({signal_942, signal_533}), .clk (clk), .r (Fresh[393]), .c ({signal_954, signal_544}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_530 ( .s ({signal_1619, signal_1607}), .b ({signal_916, signal_507}), .a ({signal_920, signal_511}), .clk (clk), .r (Fresh[394]), .c ({signal_955, signal_545}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_531 ( .s ({signal_1619, signal_1607}), .b ({signal_923, signal_514}), .a ({signal_925, signal_516}), .clk (clk), .r (Fresh[395]), .c ({signal_956, signal_546}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_532 ( .s ({signal_1619, signal_1607}), .b ({signal_929, signal_520}), .a ({signal_934, signal_525}), .clk (clk), .r (Fresh[396]), .c ({signal_957, signal_547}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_533 ( .s ({signal_1619, signal_1607}), .b ({signal_921, signal_512}), .a ({signal_939, signal_530}), .clk (clk), .r (Fresh[397]), .c ({signal_958, signal_548}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_534 ( .s ({signal_1619, signal_1607}), .b ({signal_924, signal_515}), .a ({signal_943, signal_534}), .clk (clk), .r (Fresh[398]), .c ({signal_959, signal_549}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_535 ( .s ({signal_1619, signal_1607}), .b ({signal_930, signal_521}), .a ({signal_926, signal_517}), .clk (clk), .r (Fresh[399]), .c ({signal_960, signal_550}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_536 ( .s ({signal_1619, signal_1607}), .b ({signal_938, signal_529}), .a ({signal_945, signal_536}), .clk (clk), .r (Fresh[400]), .c ({signal_961, signal_551}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_537 ( .s ({signal_1619, signal_1607}), .b ({signal_922, signal_513}), .a ({signal_941, signal_532}), .clk (clk), .r (Fresh[401]), .c ({signal_962, signal_552}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_538 ( .s ({signal_1619, signal_1607}), .b ({signal_918, signal_509}), .a ({signal_931, signal_522}), .clk (clk), .r (Fresh[402]), .c ({signal_963, signal_553}) ) ;
    buf_clk cell_788 ( .C (clk), .D (signal_1632), .Q (signal_1633) ) ;
    buf_clk cell_802 ( .C (clk), .D (signal_1646), .Q (signal_1647) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_539 ( .s ({signal_1647, signal_1633}), .b ({signal_949, signal_539}), .a ({signal_955, signal_545}), .clk (clk), .r (Fresh[403]), .c ({signal_965, signal_145}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_540 ( .s ({signal_1647, signal_1633}), .b ({signal_958, signal_548}), .a ({signal_956, signal_546}), .clk (clk), .r (Fresh[404]), .c ({signal_966, signal_148}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_541 ( .s ({signal_1647, signal_1633}), .b ({signal_953, signal_543}), .a ({signal_957, signal_547}), .clk (clk), .r (Fresh[405]), .c ({signal_967, signal_143}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_542 ( .s ({signal_1647, signal_1633}), .b ({signal_963, signal_553}), .a ({signal_961, signal_551}), .clk (clk), .r (Fresh[406]), .c ({signal_968, signal_146}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_543 ( .s ({signal_1647, signal_1633}), .b ({signal_950, signal_540}), .a ({signal_962, signal_552}), .clk (clk), .r (Fresh[407]), .c ({signal_969, signal_149}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_544 ( .s ({signal_1647, signal_1633}), .b ({signal_960, signal_550}), .a ({signal_952, signal_542}), .clk (clk), .r (Fresh[408]), .c ({signal_970, signal_144}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_545 ( .s ({signal_1647, signal_1633}), .b ({signal_948, signal_538}), .a ({signal_959, signal_549}), .clk (clk), .r (Fresh[409]), .c ({signal_971, signal_147}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_546 ( .s ({signal_1647, signal_1633}), .b ({signal_954, signal_544}), .a ({signal_951, signal_541}), .clk (clk), .r (Fresh[410]), .c ({signal_972, signal_150}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(1)) cell_0 ( .clk (clk), .D ({signal_967, signal_143}), .Q ({Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1 ( .clk (clk), .D ({signal_970, signal_144}), .Q ({Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_2 ( .clk (clk), .D ({signal_965, signal_145}), .Q ({Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3 ( .clk (clk), .D ({signal_968, signal_146}), .Q ({Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_4 ( .clk (clk), .D ({signal_971, signal_147}), .Q ({Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_5 ( .clk (clk), .D ({signal_966, signal_148}), .Q ({Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_6 ( .clk (clk), .D ({signal_969, signal_149}), .Q ({Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_7 ( .clk (clk), .D ({signal_972, signal_150}), .Q ({Y_s1[0], Y_s0[0]}) ) ;
endmodule
