
module SkinnyTop_HPC2_Pipeline_d2 ( Plaintext_s0, Key_s0, clk, rst, Key_s1, 
        Key_s2, Plaintext_s1, Plaintext_s2, Fresh, Ciphertext_s0, done, 
        Ciphertext_s1, Ciphertext_s2 );
  input [63:0] Plaintext_s0;
  input [63:0] Key_s0;
  input [63:0] Key_s1;
  input [63:0] Key_s2;
  input [63:0] Plaintext_s1;
  input [63:0] Plaintext_s2;
  input [191:0] Fresh;
  output [63:0] Ciphertext_s0;
  output [63:0] Ciphertext_s1;
  output [63:0] Ciphertext_s2;
  input clk, rst;
  output done;
  wire   SubCellInst_SboxInst_0_n3, new_AGEMA_signal_1171,
         new_AGEMA_signal_1170, SubCellInst_SboxInst_0_XX_1_,
         new_AGEMA_signal_1175, new_AGEMA_signal_1174,
         SubCellInst_SboxInst_0_XX_2_, new_AGEMA_signal_1743,
         new_AGEMA_signal_1742, SubCellInst_SboxInst_0_Q0,
         new_AGEMA_signal_1745, new_AGEMA_signal_1744,
         SubCellInst_SboxInst_0_Q1, new_AGEMA_signal_1747,
         new_AGEMA_signal_1746, SubCellInst_SboxInst_0_Q4,
         new_AGEMA_signal_1749, new_AGEMA_signal_1748,
         SubCellInst_SboxInst_0_Q6, new_AGEMA_signal_1937,
         new_AGEMA_signal_1936, SubCellInst_SboxInst_0_L1,
         new_AGEMA_signal_1751, new_AGEMA_signal_1750,
         SubCellInst_SboxInst_0_L2, SubCellInst_SboxInst_1_n3,
         new_AGEMA_signal_1183, new_AGEMA_signal_1182,
         SubCellInst_SboxInst_1_XX_1_, new_AGEMA_signal_1187,
         new_AGEMA_signal_1186, SubCellInst_SboxInst_1_XX_2_,
         new_AGEMA_signal_1755, new_AGEMA_signal_1754,
         SubCellInst_SboxInst_1_Q0, new_AGEMA_signal_1757,
         new_AGEMA_signal_1756, SubCellInst_SboxInst_1_Q1,
         new_AGEMA_signal_1759, new_AGEMA_signal_1758,
         SubCellInst_SboxInst_1_Q4, new_AGEMA_signal_1761,
         new_AGEMA_signal_1760, SubCellInst_SboxInst_1_Q6,
         new_AGEMA_signal_1943, new_AGEMA_signal_1942,
         SubCellInst_SboxInst_1_L1, new_AGEMA_signal_1763,
         new_AGEMA_signal_1762, SubCellInst_SboxInst_1_L2,
         SubCellInst_SboxInst_2_n3, new_AGEMA_signal_1195,
         new_AGEMA_signal_1194, SubCellInst_SboxInst_2_XX_1_,
         new_AGEMA_signal_1199, new_AGEMA_signal_1198,
         SubCellInst_SboxInst_2_XX_2_, new_AGEMA_signal_1767,
         new_AGEMA_signal_1766, SubCellInst_SboxInst_2_Q0,
         new_AGEMA_signal_1769, new_AGEMA_signal_1768,
         SubCellInst_SboxInst_2_Q1, new_AGEMA_signal_1771,
         new_AGEMA_signal_1770, SubCellInst_SboxInst_2_Q4,
         new_AGEMA_signal_1773, new_AGEMA_signal_1772,
         SubCellInst_SboxInst_2_Q6, new_AGEMA_signal_1949,
         new_AGEMA_signal_1948, SubCellInst_SboxInst_2_L1,
         new_AGEMA_signal_1775, new_AGEMA_signal_1774,
         SubCellInst_SboxInst_2_L2, SubCellInst_SboxInst_3_n3,
         new_AGEMA_signal_1207, new_AGEMA_signal_1206,
         SubCellInst_SboxInst_3_XX_1_, new_AGEMA_signal_1211,
         new_AGEMA_signal_1210, SubCellInst_SboxInst_3_XX_2_,
         new_AGEMA_signal_1779, new_AGEMA_signal_1778,
         SubCellInst_SboxInst_3_Q0, new_AGEMA_signal_1781,
         new_AGEMA_signal_1780, SubCellInst_SboxInst_3_Q1,
         new_AGEMA_signal_1783, new_AGEMA_signal_1782,
         SubCellInst_SboxInst_3_Q4, new_AGEMA_signal_1785,
         new_AGEMA_signal_1784, SubCellInst_SboxInst_3_Q6,
         new_AGEMA_signal_1955, new_AGEMA_signal_1954,
         SubCellInst_SboxInst_3_L1, new_AGEMA_signal_1787,
         new_AGEMA_signal_1786, SubCellInst_SboxInst_3_L2,
         SubCellInst_SboxInst_4_n3, new_AGEMA_signal_1219,
         new_AGEMA_signal_1218, SubCellInst_SboxInst_4_XX_1_,
         new_AGEMA_signal_1223, new_AGEMA_signal_1222,
         SubCellInst_SboxInst_4_XX_2_, new_AGEMA_signal_1791,
         new_AGEMA_signal_1790, SubCellInst_SboxInst_4_Q0,
         new_AGEMA_signal_1793, new_AGEMA_signal_1792,
         SubCellInst_SboxInst_4_Q1, new_AGEMA_signal_1795,
         new_AGEMA_signal_1794, SubCellInst_SboxInst_4_Q4,
         new_AGEMA_signal_1797, new_AGEMA_signal_1796,
         SubCellInst_SboxInst_4_Q6, new_AGEMA_signal_1961,
         new_AGEMA_signal_1960, SubCellInst_SboxInst_4_L1,
         new_AGEMA_signal_1799, new_AGEMA_signal_1798,
         SubCellInst_SboxInst_4_L2, SubCellInst_SboxInst_5_n3,
         new_AGEMA_signal_1231, new_AGEMA_signal_1230,
         SubCellInst_SboxInst_5_XX_1_, new_AGEMA_signal_1235,
         new_AGEMA_signal_1234, SubCellInst_SboxInst_5_XX_2_,
         new_AGEMA_signal_1803, new_AGEMA_signal_1802,
         SubCellInst_SboxInst_5_Q0, new_AGEMA_signal_1805,
         new_AGEMA_signal_1804, SubCellInst_SboxInst_5_Q1,
         new_AGEMA_signal_1807, new_AGEMA_signal_1806,
         SubCellInst_SboxInst_5_Q4, new_AGEMA_signal_1809,
         new_AGEMA_signal_1808, SubCellInst_SboxInst_5_Q6,
         new_AGEMA_signal_1967, new_AGEMA_signal_1966,
         SubCellInst_SboxInst_5_L1, new_AGEMA_signal_1811,
         new_AGEMA_signal_1810, SubCellInst_SboxInst_5_L2,
         SubCellInst_SboxInst_6_n3, new_AGEMA_signal_1243,
         new_AGEMA_signal_1242, SubCellInst_SboxInst_6_XX_1_,
         new_AGEMA_signal_1247, new_AGEMA_signal_1246,
         SubCellInst_SboxInst_6_XX_2_, new_AGEMA_signal_1815,
         new_AGEMA_signal_1814, SubCellInst_SboxInst_6_Q0,
         new_AGEMA_signal_1817, new_AGEMA_signal_1816,
         SubCellInst_SboxInst_6_Q1, new_AGEMA_signal_1819,
         new_AGEMA_signal_1818, SubCellInst_SboxInst_6_Q4,
         new_AGEMA_signal_1821, new_AGEMA_signal_1820,
         SubCellInst_SboxInst_6_Q6, new_AGEMA_signal_1973,
         new_AGEMA_signal_1972, SubCellInst_SboxInst_6_L1,
         new_AGEMA_signal_1823, new_AGEMA_signal_1822,
         SubCellInst_SboxInst_6_L2, SubCellInst_SboxInst_7_n3,
         new_AGEMA_signal_1255, new_AGEMA_signal_1254,
         SubCellInst_SboxInst_7_XX_1_, new_AGEMA_signal_1259,
         new_AGEMA_signal_1258, SubCellInst_SboxInst_7_XX_2_,
         new_AGEMA_signal_1827, new_AGEMA_signal_1826,
         SubCellInst_SboxInst_7_Q0, new_AGEMA_signal_1829,
         new_AGEMA_signal_1828, SubCellInst_SboxInst_7_Q1,
         new_AGEMA_signal_1831, new_AGEMA_signal_1830,
         SubCellInst_SboxInst_7_Q4, new_AGEMA_signal_1833,
         new_AGEMA_signal_1832, SubCellInst_SboxInst_7_Q6,
         new_AGEMA_signal_1979, new_AGEMA_signal_1978,
         SubCellInst_SboxInst_7_L1, new_AGEMA_signal_1835,
         new_AGEMA_signal_1834, SubCellInst_SboxInst_7_L2,
         SubCellInst_SboxInst_8_n3, new_AGEMA_signal_1267,
         new_AGEMA_signal_1266, SubCellInst_SboxInst_8_XX_1_,
         new_AGEMA_signal_1271, new_AGEMA_signal_1270,
         SubCellInst_SboxInst_8_XX_2_, new_AGEMA_signal_1839,
         new_AGEMA_signal_1838, SubCellInst_SboxInst_8_Q0,
         new_AGEMA_signal_1841, new_AGEMA_signal_1840,
         SubCellInst_SboxInst_8_Q1, new_AGEMA_signal_1843,
         new_AGEMA_signal_1842, SubCellInst_SboxInst_8_Q4,
         new_AGEMA_signal_1845, new_AGEMA_signal_1844,
         SubCellInst_SboxInst_8_Q6, new_AGEMA_signal_1985,
         new_AGEMA_signal_1984, SubCellInst_SboxInst_8_L1,
         new_AGEMA_signal_1847, new_AGEMA_signal_1846,
         SubCellInst_SboxInst_8_L2, SubCellInst_SboxInst_9_n3,
         new_AGEMA_signal_1279, new_AGEMA_signal_1278,
         SubCellInst_SboxInst_9_XX_1_, new_AGEMA_signal_1283,
         new_AGEMA_signal_1282, SubCellInst_SboxInst_9_XX_2_,
         new_AGEMA_signal_1851, new_AGEMA_signal_1850,
         SubCellInst_SboxInst_9_Q0, new_AGEMA_signal_1853,
         new_AGEMA_signal_1852, SubCellInst_SboxInst_9_Q1,
         new_AGEMA_signal_1855, new_AGEMA_signal_1854,
         SubCellInst_SboxInst_9_Q4, new_AGEMA_signal_1857,
         new_AGEMA_signal_1856, SubCellInst_SboxInst_9_Q6,
         new_AGEMA_signal_1991, new_AGEMA_signal_1990,
         SubCellInst_SboxInst_9_L1, new_AGEMA_signal_1859,
         new_AGEMA_signal_1858, SubCellInst_SboxInst_9_L2,
         SubCellInst_SboxInst_10_n3, new_AGEMA_signal_1291,
         new_AGEMA_signal_1290, SubCellInst_SboxInst_10_XX_1_,
         new_AGEMA_signal_1295, new_AGEMA_signal_1294,
         SubCellInst_SboxInst_10_XX_2_, new_AGEMA_signal_1863,
         new_AGEMA_signal_1862, SubCellInst_SboxInst_10_Q0,
         new_AGEMA_signal_1865, new_AGEMA_signal_1864,
         SubCellInst_SboxInst_10_Q1, new_AGEMA_signal_1867,
         new_AGEMA_signal_1866, SubCellInst_SboxInst_10_Q4,
         new_AGEMA_signal_1869, new_AGEMA_signal_1868,
         SubCellInst_SboxInst_10_Q6, new_AGEMA_signal_1997,
         new_AGEMA_signal_1996, SubCellInst_SboxInst_10_L1,
         new_AGEMA_signal_1871, new_AGEMA_signal_1870,
         SubCellInst_SboxInst_10_L2, SubCellInst_SboxInst_11_n3,
         new_AGEMA_signal_1303, new_AGEMA_signal_1302,
         SubCellInst_SboxInst_11_XX_1_, new_AGEMA_signal_1307,
         new_AGEMA_signal_1306, SubCellInst_SboxInst_11_XX_2_,
         new_AGEMA_signal_1875, new_AGEMA_signal_1874,
         SubCellInst_SboxInst_11_Q0, new_AGEMA_signal_1877,
         new_AGEMA_signal_1876, SubCellInst_SboxInst_11_Q1,
         new_AGEMA_signal_1879, new_AGEMA_signal_1878,
         SubCellInst_SboxInst_11_Q4, new_AGEMA_signal_1881,
         new_AGEMA_signal_1880, SubCellInst_SboxInst_11_Q6,
         new_AGEMA_signal_2003, new_AGEMA_signal_2002,
         SubCellInst_SboxInst_11_L1, new_AGEMA_signal_1883,
         new_AGEMA_signal_1882, SubCellInst_SboxInst_11_L2,
         SubCellInst_SboxInst_12_n3, new_AGEMA_signal_1315,
         new_AGEMA_signal_1314, SubCellInst_SboxInst_12_XX_1_,
         new_AGEMA_signal_1319, new_AGEMA_signal_1318,
         SubCellInst_SboxInst_12_XX_2_, new_AGEMA_signal_1887,
         new_AGEMA_signal_1886, SubCellInst_SboxInst_12_Q0,
         new_AGEMA_signal_1889, new_AGEMA_signal_1888,
         SubCellInst_SboxInst_12_Q1, new_AGEMA_signal_1891,
         new_AGEMA_signal_1890, SubCellInst_SboxInst_12_Q4,
         new_AGEMA_signal_1893, new_AGEMA_signal_1892,
         SubCellInst_SboxInst_12_Q6, new_AGEMA_signal_2009,
         new_AGEMA_signal_2008, SubCellInst_SboxInst_12_L1,
         new_AGEMA_signal_1895, new_AGEMA_signal_1894,
         SubCellInst_SboxInst_12_L2, SubCellInst_SboxInst_13_n3,
         new_AGEMA_signal_1327, new_AGEMA_signal_1326,
         SubCellInst_SboxInst_13_XX_1_, new_AGEMA_signal_1331,
         new_AGEMA_signal_1330, SubCellInst_SboxInst_13_XX_2_,
         new_AGEMA_signal_1899, new_AGEMA_signal_1898,
         SubCellInst_SboxInst_13_Q0, new_AGEMA_signal_1901,
         new_AGEMA_signal_1900, SubCellInst_SboxInst_13_Q1,
         new_AGEMA_signal_1903, new_AGEMA_signal_1902,
         SubCellInst_SboxInst_13_Q4, new_AGEMA_signal_1905,
         new_AGEMA_signal_1904, SubCellInst_SboxInst_13_Q6,
         new_AGEMA_signal_2015, new_AGEMA_signal_2014,
         SubCellInst_SboxInst_13_L1, new_AGEMA_signal_1907,
         new_AGEMA_signal_1906, SubCellInst_SboxInst_13_L2,
         SubCellInst_SboxInst_14_n3, new_AGEMA_signal_1339,
         new_AGEMA_signal_1338, SubCellInst_SboxInst_14_XX_1_,
         new_AGEMA_signal_1343, new_AGEMA_signal_1342,
         SubCellInst_SboxInst_14_XX_2_, new_AGEMA_signal_1911,
         new_AGEMA_signal_1910, SubCellInst_SboxInst_14_Q0,
         new_AGEMA_signal_1913, new_AGEMA_signal_1912,
         SubCellInst_SboxInst_14_Q1, new_AGEMA_signal_1915,
         new_AGEMA_signal_1914, SubCellInst_SboxInst_14_Q4,
         new_AGEMA_signal_1917, new_AGEMA_signal_1916,
         SubCellInst_SboxInst_14_Q6, new_AGEMA_signal_2021,
         new_AGEMA_signal_2020, SubCellInst_SboxInst_14_L1,
         new_AGEMA_signal_1919, new_AGEMA_signal_1918,
         SubCellInst_SboxInst_14_L2, SubCellInst_SboxInst_15_n3,
         new_AGEMA_signal_1351, new_AGEMA_signal_1350,
         SubCellInst_SboxInst_15_XX_1_, new_AGEMA_signal_1355,
         new_AGEMA_signal_1354, SubCellInst_SboxInst_15_XX_2_,
         new_AGEMA_signal_1923, new_AGEMA_signal_1922,
         SubCellInst_SboxInst_15_Q0, new_AGEMA_signal_1925,
         new_AGEMA_signal_1924, SubCellInst_SboxInst_15_Q1,
         new_AGEMA_signal_1927, new_AGEMA_signal_1926,
         SubCellInst_SboxInst_15_Q4, new_AGEMA_signal_1929,
         new_AGEMA_signal_1928, SubCellInst_SboxInst_15_Q6,
         new_AGEMA_signal_2027, new_AGEMA_signal_2026,
         SubCellInst_SboxInst_15_L1, new_AGEMA_signal_1931,
         new_AGEMA_signal_1930, SubCellInst_SboxInst_15_L2,
         new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1357,
         new_AGEMA_signal_1356, new_AGEMA_signal_1367, new_AGEMA_signal_1366,
         new_AGEMA_signal_1363, new_AGEMA_signal_1362, new_AGEMA_signal_1373,
         new_AGEMA_signal_1372, new_AGEMA_signal_1369, new_AGEMA_signal_1368,
         new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1375,
         new_AGEMA_signal_1374, new_AGEMA_signal_1385, new_AGEMA_signal_1384,
         new_AGEMA_signal_1381, new_AGEMA_signal_1380, new_AGEMA_signal_1391,
         new_AGEMA_signal_1390, new_AGEMA_signal_1387, new_AGEMA_signal_1386,
         new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1393,
         new_AGEMA_signal_1392, new_AGEMA_signal_1403, new_AGEMA_signal_1402,
         new_AGEMA_signal_1399, new_AGEMA_signal_1398, new_AGEMA_signal_1409,
         new_AGEMA_signal_1408, new_AGEMA_signal_1405, new_AGEMA_signal_1404,
         new_AGEMA_signal_1415, new_AGEMA_signal_1414, new_AGEMA_signal_1411,
         new_AGEMA_signal_1410, new_AGEMA_signal_1421, new_AGEMA_signal_1420,
         new_AGEMA_signal_1417, new_AGEMA_signal_1416, new_AGEMA_signal_1427,
         new_AGEMA_signal_1426, new_AGEMA_signal_1423, new_AGEMA_signal_1422,
         new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1429,
         new_AGEMA_signal_1428, new_AGEMA_signal_1439, new_AGEMA_signal_1438,
         new_AGEMA_signal_1435, new_AGEMA_signal_1434, new_AGEMA_signal_1445,
         new_AGEMA_signal_1444, new_AGEMA_signal_1441, new_AGEMA_signal_1440,
         new_AGEMA_signal_1451, new_AGEMA_signal_1450, new_AGEMA_signal_1447,
         new_AGEMA_signal_1446, new_AGEMA_signal_1457, new_AGEMA_signal_1456,
         new_AGEMA_signal_1453, new_AGEMA_signal_1452, new_AGEMA_signal_1463,
         new_AGEMA_signal_1462, new_AGEMA_signal_1459, new_AGEMA_signal_1458,
         new_AGEMA_signal_1469, new_AGEMA_signal_1468, new_AGEMA_signal_1465,
         new_AGEMA_signal_1464, new_AGEMA_signal_1475, new_AGEMA_signal_1474,
         new_AGEMA_signal_1471, new_AGEMA_signal_1470, new_AGEMA_signal_1481,
         new_AGEMA_signal_1480, new_AGEMA_signal_1477, new_AGEMA_signal_1476,
         new_AGEMA_signal_1487, new_AGEMA_signal_1486, new_AGEMA_signal_1483,
         new_AGEMA_signal_1482, new_AGEMA_signal_1493, new_AGEMA_signal_1492,
         new_AGEMA_signal_1489, new_AGEMA_signal_1488, new_AGEMA_signal_1499,
         new_AGEMA_signal_1498, new_AGEMA_signal_1495, new_AGEMA_signal_1494,
         new_AGEMA_signal_1505, new_AGEMA_signal_1504, new_AGEMA_signal_1501,
         new_AGEMA_signal_1500, new_AGEMA_signal_1511, new_AGEMA_signal_1510,
         new_AGEMA_signal_1507, new_AGEMA_signal_1506, new_AGEMA_signal_1517,
         new_AGEMA_signal_1516, new_AGEMA_signal_1513, new_AGEMA_signal_1512,
         new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1519,
         new_AGEMA_signal_1518, new_AGEMA_signal_1529, new_AGEMA_signal_1528,
         new_AGEMA_signal_1525, new_AGEMA_signal_1524, new_AGEMA_signal_1535,
         new_AGEMA_signal_1534, new_AGEMA_signal_1531, new_AGEMA_signal_1530,
         new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1537,
         new_AGEMA_signal_1536, new_AGEMA_signal_1547, new_AGEMA_signal_1546,
         new_AGEMA_signal_1543, new_AGEMA_signal_1542, new_AGEMA_signal_1553,
         new_AGEMA_signal_1552, new_AGEMA_signal_1549, new_AGEMA_signal_1548,
         new_AGEMA_signal_1559, new_AGEMA_signal_1558, new_AGEMA_signal_1555,
         new_AGEMA_signal_1554, new_AGEMA_signal_1565, new_AGEMA_signal_1564,
         new_AGEMA_signal_1561, new_AGEMA_signal_1560, new_AGEMA_signal_1571,
         new_AGEMA_signal_1570, new_AGEMA_signal_1567, new_AGEMA_signal_1566,
         new_AGEMA_signal_1577, new_AGEMA_signal_1576, new_AGEMA_signal_1573,
         new_AGEMA_signal_1572, new_AGEMA_signal_1583, new_AGEMA_signal_1582,
         new_AGEMA_signal_1579, new_AGEMA_signal_1578, new_AGEMA_signal_1589,
         new_AGEMA_signal_1588, new_AGEMA_signal_1585, new_AGEMA_signal_1584,
         new_AGEMA_signal_1595, new_AGEMA_signal_1594, new_AGEMA_signal_1591,
         new_AGEMA_signal_1590, new_AGEMA_signal_1601, new_AGEMA_signal_1600,
         new_AGEMA_signal_1597, new_AGEMA_signal_1596, new_AGEMA_signal_1607,
         new_AGEMA_signal_1606, new_AGEMA_signal_1603, new_AGEMA_signal_1602,
         new_AGEMA_signal_1613, new_AGEMA_signal_1612, new_AGEMA_signal_1609,
         new_AGEMA_signal_1608, new_AGEMA_signal_1619, new_AGEMA_signal_1618,
         new_AGEMA_signal_1615, new_AGEMA_signal_1614, new_AGEMA_signal_1625,
         new_AGEMA_signal_1624, new_AGEMA_signal_1621, new_AGEMA_signal_1620,
         new_AGEMA_signal_1631, new_AGEMA_signal_1630, new_AGEMA_signal_1627,
         new_AGEMA_signal_1626, new_AGEMA_signal_1637, new_AGEMA_signal_1636,
         new_AGEMA_signal_1633, new_AGEMA_signal_1632, new_AGEMA_signal_1643,
         new_AGEMA_signal_1642, new_AGEMA_signal_1639, new_AGEMA_signal_1638,
         new_AGEMA_signal_1649, new_AGEMA_signal_1648, new_AGEMA_signal_1645,
         new_AGEMA_signal_1644, new_AGEMA_signal_1655, new_AGEMA_signal_1654,
         new_AGEMA_signal_1651, new_AGEMA_signal_1650, new_AGEMA_signal_1661,
         new_AGEMA_signal_1660, new_AGEMA_signal_1657, new_AGEMA_signal_1656,
         new_AGEMA_signal_1667, new_AGEMA_signal_1666, new_AGEMA_signal_1663,
         new_AGEMA_signal_1662, new_AGEMA_signal_1673, new_AGEMA_signal_1672,
         new_AGEMA_signal_1669, new_AGEMA_signal_1668, new_AGEMA_signal_1679,
         new_AGEMA_signal_1678, new_AGEMA_signal_1675, new_AGEMA_signal_1674,
         new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1681,
         new_AGEMA_signal_1680, new_AGEMA_signal_1691, new_AGEMA_signal_1690,
         new_AGEMA_signal_1687, new_AGEMA_signal_1686, new_AGEMA_signal_1697,
         new_AGEMA_signal_1696, new_AGEMA_signal_1693, new_AGEMA_signal_1692,
         new_AGEMA_signal_1703, new_AGEMA_signal_1702, new_AGEMA_signal_1699,
         new_AGEMA_signal_1698, new_AGEMA_signal_1709, new_AGEMA_signal_1708,
         new_AGEMA_signal_1705, new_AGEMA_signal_1704, new_AGEMA_signal_1715,
         new_AGEMA_signal_1714, new_AGEMA_signal_1711, new_AGEMA_signal_1710,
         new_AGEMA_signal_1721, new_AGEMA_signal_1720, new_AGEMA_signal_1717,
         new_AGEMA_signal_1716, new_AGEMA_signal_1727, new_AGEMA_signal_1726,
         new_AGEMA_signal_1723, new_AGEMA_signal_1722, new_AGEMA_signal_1733,
         new_AGEMA_signal_1732, new_AGEMA_signal_1729, new_AGEMA_signal_1728,
         new_AGEMA_signal_1739, new_AGEMA_signal_1738, new_AGEMA_signal_1735,
         new_AGEMA_signal_1734, FSM_1, new_AGEMA_signal_3278,
         new_AGEMA_signal_3280, new_AGEMA_signal_3282, new_AGEMA_signal_3284,
         new_AGEMA_signal_3286, new_AGEMA_signal_3288, new_AGEMA_signal_3290,
         new_AGEMA_signal_3292, new_AGEMA_signal_3294, new_AGEMA_signal_3296,
         new_AGEMA_signal_3298, new_AGEMA_signal_3300, new_AGEMA_signal_3302,
         new_AGEMA_signal_3304, new_AGEMA_signal_3306, new_AGEMA_signal_3308,
         new_AGEMA_signal_3310, new_AGEMA_signal_3312, new_AGEMA_signal_3314,
         new_AGEMA_signal_3316, new_AGEMA_signal_3318, new_AGEMA_signal_3320,
         new_AGEMA_signal_3322, new_AGEMA_signal_3324, new_AGEMA_signal_3326,
         new_AGEMA_signal_3328, new_AGEMA_signal_3330, new_AGEMA_signal_3332,
         new_AGEMA_signal_3334, new_AGEMA_signal_3336, new_AGEMA_signal_3338,
         new_AGEMA_signal_3340, new_AGEMA_signal_3342, new_AGEMA_signal_3344,
         new_AGEMA_signal_3346, new_AGEMA_signal_3348, new_AGEMA_signal_3350,
         new_AGEMA_signal_3352, new_AGEMA_signal_3354, new_AGEMA_signal_3356,
         new_AGEMA_signal_3358, new_AGEMA_signal_3360, new_AGEMA_signal_3362,
         new_AGEMA_signal_3364, new_AGEMA_signal_3366, new_AGEMA_signal_3368,
         new_AGEMA_signal_3370, new_AGEMA_signal_3372, new_AGEMA_signal_3374,
         new_AGEMA_signal_3376, new_AGEMA_signal_3378, new_AGEMA_signal_3380,
         new_AGEMA_signal_3382, new_AGEMA_signal_3384, new_AGEMA_signal_3386,
         new_AGEMA_signal_3388, new_AGEMA_signal_3390, new_AGEMA_signal_3392,
         new_AGEMA_signal_3394, new_AGEMA_signal_3396, new_AGEMA_signal_3398,
         new_AGEMA_signal_3400, new_AGEMA_signal_3402, new_AGEMA_signal_3404,
         new_AGEMA_signal_3406, new_AGEMA_signal_3408, new_AGEMA_signal_3410,
         new_AGEMA_signal_3412, new_AGEMA_signal_3414, new_AGEMA_signal_3416,
         new_AGEMA_signal_3418, new_AGEMA_signal_3420, new_AGEMA_signal_3422,
         new_AGEMA_signal_3424, new_AGEMA_signal_3426, new_AGEMA_signal_3428,
         new_AGEMA_signal_3430, new_AGEMA_signal_3432, new_AGEMA_signal_3434,
         new_AGEMA_signal_3436, new_AGEMA_signal_3438, new_AGEMA_signal_3440,
         new_AGEMA_signal_3442, new_AGEMA_signal_3444, new_AGEMA_signal_3446,
         new_AGEMA_signal_3448, new_AGEMA_signal_3450, new_AGEMA_signal_3452,
         new_AGEMA_signal_3454, new_AGEMA_signal_3456, new_AGEMA_signal_3458,
         new_AGEMA_signal_3460, new_AGEMA_signal_3462, new_AGEMA_signal_3464,
         new_AGEMA_signal_3466, new_AGEMA_signal_3468, new_AGEMA_signal_3470,
         new_AGEMA_signal_3472, new_AGEMA_signal_3474, new_AGEMA_signal_3476,
         new_AGEMA_signal_3478, new_AGEMA_signal_3480, new_AGEMA_signal_3482,
         new_AGEMA_signal_3484, new_AGEMA_signal_3486, new_AGEMA_signal_3488,
         new_AGEMA_signal_3490, new_AGEMA_signal_3492, new_AGEMA_signal_3494,
         new_AGEMA_signal_3496, new_AGEMA_signal_3498, new_AGEMA_signal_3500,
         new_AGEMA_signal_3502, new_AGEMA_signal_3504, new_AGEMA_signal_3506,
         new_AGEMA_signal_3508, new_AGEMA_signal_3510, new_AGEMA_signal_3512,
         new_AGEMA_signal_3514, new_AGEMA_signal_3516, new_AGEMA_signal_3518,
         new_AGEMA_signal_3520, new_AGEMA_signal_3522, new_AGEMA_signal_3524,
         new_AGEMA_signal_3526, new_AGEMA_signal_3528, new_AGEMA_signal_3530,
         new_AGEMA_signal_3532, new_AGEMA_signal_3534, new_AGEMA_signal_3536,
         new_AGEMA_signal_3538, new_AGEMA_signal_3540, new_AGEMA_signal_3542,
         new_AGEMA_signal_3544, new_AGEMA_signal_3546, new_AGEMA_signal_3548,
         new_AGEMA_signal_3550, new_AGEMA_signal_3552, new_AGEMA_signal_3554,
         new_AGEMA_signal_3556, new_AGEMA_signal_3558, new_AGEMA_signal_3560,
         new_AGEMA_signal_3562, new_AGEMA_signal_3564, new_AGEMA_signal_3566,
         new_AGEMA_signal_3568, new_AGEMA_signal_3570, new_AGEMA_signal_3572,
         new_AGEMA_signal_3574, new_AGEMA_signal_3576, new_AGEMA_signal_3578,
         new_AGEMA_signal_3580, new_AGEMA_signal_3582, new_AGEMA_signal_3584,
         new_AGEMA_signal_3586, new_AGEMA_signal_3588, new_AGEMA_signal_3590,
         new_AGEMA_signal_3592, new_AGEMA_signal_3594, new_AGEMA_signal_3596,
         new_AGEMA_signal_3598, new_AGEMA_signal_3600, new_AGEMA_signal_3602,
         new_AGEMA_signal_3604, new_AGEMA_signal_3606, new_AGEMA_signal_3608,
         new_AGEMA_signal_3610, new_AGEMA_signal_3612, new_AGEMA_signal_3614,
         new_AGEMA_signal_3616, new_AGEMA_signal_3618, new_AGEMA_signal_3620,
         new_AGEMA_signal_3622, new_AGEMA_signal_3624, new_AGEMA_signal_3626,
         new_AGEMA_signal_3628, new_AGEMA_signal_3630, new_AGEMA_signal_3632,
         new_AGEMA_signal_3634, new_AGEMA_signal_3636, new_AGEMA_signal_3638,
         new_AGEMA_signal_3640, new_AGEMA_signal_3642, new_AGEMA_signal_3644,
         new_AGEMA_signal_3646, new_AGEMA_signal_3648, new_AGEMA_signal_3650,
         new_AGEMA_signal_3652, new_AGEMA_signal_3654, new_AGEMA_signal_3656,
         new_AGEMA_signal_3658, new_AGEMA_signal_3660, new_AGEMA_signal_3662,
         new_AGEMA_signal_3664, new_AGEMA_signal_3666, new_AGEMA_signal_3668,
         new_AGEMA_signal_3670, new_AGEMA_signal_3672, new_AGEMA_signal_3674,
         new_AGEMA_signal_3676, new_AGEMA_signal_3678, new_AGEMA_signal_3680,
         new_AGEMA_signal_3682, new_AGEMA_signal_3684, new_AGEMA_signal_3686,
         new_AGEMA_signal_3688, new_AGEMA_signal_3690, new_AGEMA_signal_3692,
         new_AGEMA_signal_3694, new_AGEMA_signal_3696, new_AGEMA_signal_3698,
         new_AGEMA_signal_3700, new_AGEMA_signal_3702, new_AGEMA_signal_3704,
         new_AGEMA_signal_3706, new_AGEMA_signal_3708, new_AGEMA_signal_3710,
         new_AGEMA_signal_3712, new_AGEMA_signal_3714, new_AGEMA_signal_3716,
         new_AGEMA_signal_3718, new_AGEMA_signal_3720, new_AGEMA_signal_3722,
         new_AGEMA_signal_3724, new_AGEMA_signal_3726, new_AGEMA_signal_3728,
         new_AGEMA_signal_3730, new_AGEMA_signal_3732, new_AGEMA_signal_3734,
         new_AGEMA_signal_3736, new_AGEMA_signal_3738, new_AGEMA_signal_3740,
         new_AGEMA_signal_3742, new_AGEMA_signal_3744, new_AGEMA_signal_3746,
         new_AGEMA_signal_3748, new_AGEMA_signal_3750, new_AGEMA_signal_3752,
         new_AGEMA_signal_3754, new_AGEMA_signal_3756, new_AGEMA_signal_3758,
         new_AGEMA_signal_3760, new_AGEMA_signal_3762, new_AGEMA_signal_3764,
         new_AGEMA_signal_3766, new_AGEMA_signal_3768, new_AGEMA_signal_3770,
         new_AGEMA_signal_3772, new_AGEMA_signal_3774, new_AGEMA_signal_3776,
         new_AGEMA_signal_3778, new_AGEMA_signal_3780, new_AGEMA_signal_3782,
         new_AGEMA_signal_3784, new_AGEMA_signal_3786, new_AGEMA_signal_3788,
         new_AGEMA_signal_3790, new_AGEMA_signal_3792, new_AGEMA_signal_3794,
         new_AGEMA_signal_3796, new_AGEMA_signal_3798, new_AGEMA_signal_3800,
         new_AGEMA_signal_3802, new_AGEMA_signal_3804, new_AGEMA_signal_3806,
         new_AGEMA_signal_3808, new_AGEMA_signal_3810, new_AGEMA_signal_3812,
         new_AGEMA_signal_3814, new_AGEMA_signal_3816, new_AGEMA_signal_3818,
         new_AGEMA_signal_3820, new_AGEMA_signal_3822, new_AGEMA_signal_3824,
         new_AGEMA_signal_3826, new_AGEMA_signal_3828, new_AGEMA_signal_3830,
         new_AGEMA_signal_3832, new_AGEMA_signal_3834, new_AGEMA_signal_3836,
         new_AGEMA_signal_3838, new_AGEMA_signal_3840, new_AGEMA_signal_3842,
         new_AGEMA_signal_3844, new_AGEMA_signal_3846, new_AGEMA_signal_3848,
         new_AGEMA_signal_3850, new_AGEMA_signal_3852, new_AGEMA_signal_3854,
         new_AGEMA_signal_3856, new_AGEMA_signal_3858, new_AGEMA_signal_3860,
         new_AGEMA_signal_3862, new_AGEMA_signal_3864, new_AGEMA_signal_3866,
         new_AGEMA_signal_3868, new_AGEMA_signal_3870, new_AGEMA_signal_3872,
         new_AGEMA_signal_3874, new_AGEMA_signal_3876, new_AGEMA_signal_3878,
         new_AGEMA_signal_3880, new_AGEMA_signal_3882, new_AGEMA_signal_3884,
         new_AGEMA_signal_3886, new_AGEMA_signal_3888, new_AGEMA_signal_3890,
         new_AGEMA_signal_3892, new_AGEMA_signal_3894, new_AGEMA_signal_3896,
         new_AGEMA_signal_3898, new_AGEMA_signal_3900, new_AGEMA_signal_3902,
         new_AGEMA_signal_3904, new_AGEMA_signal_3906, new_AGEMA_signal_3908,
         new_AGEMA_signal_3910, new_AGEMA_signal_3912, new_AGEMA_signal_3914,
         new_AGEMA_signal_3916, new_AGEMA_signal_3918, new_AGEMA_signal_3920,
         new_AGEMA_signal_3922, new_AGEMA_signal_3924, new_AGEMA_signal_3926,
         new_AGEMA_signal_3928, new_AGEMA_signal_3930, new_AGEMA_signal_3932,
         new_AGEMA_signal_3934, new_AGEMA_signal_3936, new_AGEMA_signal_3938,
         new_AGEMA_signal_3940, new_AGEMA_signal_3942, new_AGEMA_signal_3944,
         new_AGEMA_signal_3946, new_AGEMA_signal_3948, new_AGEMA_signal_3950,
         new_AGEMA_signal_3952, new_AGEMA_signal_3954, new_AGEMA_signal_3958,
         new_AGEMA_signal_3962, new_AGEMA_signal_3966, new_AGEMA_signal_3970,
         new_AGEMA_signal_3974, new_AGEMA_signal_3978, new_AGEMA_signal_3982,
         new_AGEMA_signal_3986, new_AGEMA_signal_3990, new_AGEMA_signal_3994,
         new_AGEMA_signal_3998, new_AGEMA_signal_4002, new_AGEMA_signal_4006,
         new_AGEMA_signal_4010, new_AGEMA_signal_4014, new_AGEMA_signal_4018,
         new_AGEMA_signal_4022, new_AGEMA_signal_4026, new_AGEMA_signal_4030,
         new_AGEMA_signal_4034, new_AGEMA_signal_4038, new_AGEMA_signal_4042,
         new_AGEMA_signal_4046, new_AGEMA_signal_4050, new_AGEMA_signal_4054,
         new_AGEMA_signal_4058, new_AGEMA_signal_4062, new_AGEMA_signal_4066,
         new_AGEMA_signal_4070, new_AGEMA_signal_4074, new_AGEMA_signal_4078,
         new_AGEMA_signal_4082, new_AGEMA_signal_4086, new_AGEMA_signal_4090,
         new_AGEMA_signal_4094, new_AGEMA_signal_4098, new_AGEMA_signal_4102,
         new_AGEMA_signal_4106, new_AGEMA_signal_4110, new_AGEMA_signal_4114,
         new_AGEMA_signal_4118, new_AGEMA_signal_4122, new_AGEMA_signal_4126,
         new_AGEMA_signal_4130, new_AGEMA_signal_4134, new_AGEMA_signal_4138,
         new_AGEMA_signal_4142, new_AGEMA_signal_4146, new_AGEMA_signal_4150,
         new_AGEMA_signal_4154, new_AGEMA_signal_4158, new_AGEMA_signal_4162,
         new_AGEMA_signal_4166, new_AGEMA_signal_4170, new_AGEMA_signal_4174,
         new_AGEMA_signal_4178, new_AGEMA_signal_4182, new_AGEMA_signal_4186,
         new_AGEMA_signal_4190, new_AGEMA_signal_4194, new_AGEMA_signal_4198,
         new_AGEMA_signal_4202, new_AGEMA_signal_4206, new_AGEMA_signal_4210,
         new_AGEMA_signal_4214, new_AGEMA_signal_4218, new_AGEMA_signal_4222,
         new_AGEMA_signal_4226, new_AGEMA_signal_4230, new_AGEMA_signal_4234,
         new_AGEMA_signal_4238, new_AGEMA_signal_4242, new_AGEMA_signal_4246,
         new_AGEMA_signal_4250, new_AGEMA_signal_4254, new_AGEMA_signal_4258,
         new_AGEMA_signal_4262, new_AGEMA_signal_4266, new_AGEMA_signal_4270,
         new_AGEMA_signal_4274, new_AGEMA_signal_4278, new_AGEMA_signal_4282,
         new_AGEMA_signal_4286, new_AGEMA_signal_4290, new_AGEMA_signal_4294,
         new_AGEMA_signal_4298, new_AGEMA_signal_4302, new_AGEMA_signal_4306,
         new_AGEMA_signal_4310, new_AGEMA_signal_4314, new_AGEMA_signal_4318,
         new_AGEMA_signal_4322, new_AGEMA_signal_4326, new_AGEMA_signal_4330,
         new_AGEMA_signal_4334, new_AGEMA_signal_4338, new_AGEMA_signal_4342,
         new_AGEMA_signal_4344, new_AGEMA_signal_4346, new_AGEMA_signal_4354,
         new_AGEMA_signal_4356, new_AGEMA_signal_4358, new_AGEMA_signal_4360,
         new_AGEMA_signal_4364, new_AGEMA_signal_4368, new_AGEMA_signal_4378,
         new_AGEMA_signal_4380, new_AGEMA_signal_4382, new_AGEMA_signal_4390,
         new_AGEMA_signal_4392, new_AGEMA_signal_4394, new_AGEMA_signal_4396,
         new_AGEMA_signal_4400, new_AGEMA_signal_4404, new_AGEMA_signal_4414,
         new_AGEMA_signal_4416, new_AGEMA_signal_4418, new_AGEMA_signal_4426,
         new_AGEMA_signal_4428, new_AGEMA_signal_4430, new_AGEMA_signal_4432,
         new_AGEMA_signal_4436, new_AGEMA_signal_4440, new_AGEMA_signal_4450,
         new_AGEMA_signal_4452, new_AGEMA_signal_4454, new_AGEMA_signal_4462,
         new_AGEMA_signal_4464, new_AGEMA_signal_4466, new_AGEMA_signal_4468,
         new_AGEMA_signal_4472, new_AGEMA_signal_4476, new_AGEMA_signal_4486,
         new_AGEMA_signal_4488, new_AGEMA_signal_4490, new_AGEMA_signal_4498,
         new_AGEMA_signal_4500, new_AGEMA_signal_4502, new_AGEMA_signal_4504,
         new_AGEMA_signal_4508, new_AGEMA_signal_4512, new_AGEMA_signal_4522,
         new_AGEMA_signal_4524, new_AGEMA_signal_4526, new_AGEMA_signal_4534,
         new_AGEMA_signal_4536, new_AGEMA_signal_4538, new_AGEMA_signal_4540,
         new_AGEMA_signal_4544, new_AGEMA_signal_4548, new_AGEMA_signal_4558,
         new_AGEMA_signal_4560, new_AGEMA_signal_4562, new_AGEMA_signal_4570,
         new_AGEMA_signal_4572, new_AGEMA_signal_4574, new_AGEMA_signal_4576,
         new_AGEMA_signal_4580, new_AGEMA_signal_4584, new_AGEMA_signal_4594,
         new_AGEMA_signal_4596, new_AGEMA_signal_4598, new_AGEMA_signal_4606,
         new_AGEMA_signal_4608, new_AGEMA_signal_4610, new_AGEMA_signal_4612,
         new_AGEMA_signal_4616, new_AGEMA_signal_4620, new_AGEMA_signal_4630,
         new_AGEMA_signal_4632, new_AGEMA_signal_4634, new_AGEMA_signal_4642,
         new_AGEMA_signal_4644, new_AGEMA_signal_4646, new_AGEMA_signal_4648,
         new_AGEMA_signal_4652, new_AGEMA_signal_4656, new_AGEMA_signal_4666,
         new_AGEMA_signal_4668, new_AGEMA_signal_4670, new_AGEMA_signal_4678,
         new_AGEMA_signal_4680, new_AGEMA_signal_4682, new_AGEMA_signal_4684,
         new_AGEMA_signal_4688, new_AGEMA_signal_4692, new_AGEMA_signal_4702,
         new_AGEMA_signal_4704, new_AGEMA_signal_4706, new_AGEMA_signal_4714,
         new_AGEMA_signal_4716, new_AGEMA_signal_4718, new_AGEMA_signal_4720,
         new_AGEMA_signal_4724, new_AGEMA_signal_4728, new_AGEMA_signal_4738,
         new_AGEMA_signal_4740, new_AGEMA_signal_4742, new_AGEMA_signal_4750,
         new_AGEMA_signal_4752, new_AGEMA_signal_4754, new_AGEMA_signal_4756,
         new_AGEMA_signal_4760, new_AGEMA_signal_4764, new_AGEMA_signal_4774,
         new_AGEMA_signal_4776, new_AGEMA_signal_4778, new_AGEMA_signal_4786,
         new_AGEMA_signal_4788, new_AGEMA_signal_4790, new_AGEMA_signal_4792,
         new_AGEMA_signal_4796, new_AGEMA_signal_4800, new_AGEMA_signal_4810,
         new_AGEMA_signal_4812, new_AGEMA_signal_4814, new_AGEMA_signal_4822,
         new_AGEMA_signal_4824, new_AGEMA_signal_4826, new_AGEMA_signal_4828,
         new_AGEMA_signal_4832, new_AGEMA_signal_4836, new_AGEMA_signal_4846,
         new_AGEMA_signal_4848, new_AGEMA_signal_4850, new_AGEMA_signal_4858,
         new_AGEMA_signal_4860, new_AGEMA_signal_4862, new_AGEMA_signal_4864,
         new_AGEMA_signal_4868, new_AGEMA_signal_4872, new_AGEMA_signal_4882,
         new_AGEMA_signal_4884, new_AGEMA_signal_4886, new_AGEMA_signal_4894,
         new_AGEMA_signal_4896, new_AGEMA_signal_4898, new_AGEMA_signal_4900,
         new_AGEMA_signal_4904, new_AGEMA_signal_4908, new_AGEMA_signal_4918,
         new_AGEMA_signal_4922, new_AGEMA_signal_4926, new_AGEMA_signal_4930,
         new_AGEMA_signal_4934, new_AGEMA_signal_4938, new_AGEMA_signal_4942,
         new_AGEMA_signal_4946, new_AGEMA_signal_4950, new_AGEMA_signal_4954,
         new_AGEMA_signal_4958, new_AGEMA_signal_4962, new_AGEMA_signal_4966,
         new_AGEMA_signal_4970, new_AGEMA_signal_4974, new_AGEMA_signal_4978,
         new_AGEMA_signal_4982, new_AGEMA_signal_4986, new_AGEMA_signal_4990,
         new_AGEMA_signal_4994, new_AGEMA_signal_4998, new_AGEMA_signal_5002,
         new_AGEMA_signal_5006, new_AGEMA_signal_5010, new_AGEMA_signal_5014,
         new_AGEMA_signal_5018, new_AGEMA_signal_5022, new_AGEMA_signal_5026,
         new_AGEMA_signal_5030, new_AGEMA_signal_5034, new_AGEMA_signal_5038,
         new_AGEMA_signal_5042, new_AGEMA_signal_5046, new_AGEMA_signal_5050,
         new_AGEMA_signal_5054, new_AGEMA_signal_5058, new_AGEMA_signal_5062,
         new_AGEMA_signal_5066, new_AGEMA_signal_5070, new_AGEMA_signal_5074,
         new_AGEMA_signal_5078, new_AGEMA_signal_5082, new_AGEMA_signal_5086,
         new_AGEMA_signal_5090, new_AGEMA_signal_5094, new_AGEMA_signal_5098,
         new_AGEMA_signal_5102, new_AGEMA_signal_5106, new_AGEMA_signal_5110,
         new_AGEMA_signal_5114, new_AGEMA_signal_5118, new_AGEMA_signal_5122,
         new_AGEMA_signal_5318, new_AGEMA_signal_5322, new_AGEMA_signal_5326,
         new_AGEMA_signal_5330, new_AGEMA_signal_5334, new_AGEMA_signal_5338,
         new_AGEMA_signal_5342, new_AGEMA_signal_5346, new_AGEMA_signal_5350,
         new_AGEMA_signal_5354, new_AGEMA_signal_5358, new_AGEMA_signal_5362,
         new_AGEMA_signal_5366, new_AGEMA_signal_5370, new_AGEMA_signal_5374,
         new_AGEMA_signal_5378, new_AGEMA_signal_5382, new_AGEMA_signal_5386,
         new_AGEMA_signal_5390, new_AGEMA_signal_5394, new_AGEMA_signal_5398,
         new_AGEMA_signal_5402, new_AGEMA_signal_5406, new_AGEMA_signal_5410,
         new_AGEMA_signal_5414, new_AGEMA_signal_5418, new_AGEMA_signal_5422,
         new_AGEMA_signal_5426, new_AGEMA_signal_5430, new_AGEMA_signal_5434,
         new_AGEMA_signal_5438, new_AGEMA_signal_5442, new_AGEMA_signal_5446,
         new_AGEMA_signal_5450, new_AGEMA_signal_5454, new_AGEMA_signal_5458,
         new_AGEMA_signal_5462, new_AGEMA_signal_5466, new_AGEMA_signal_5470,
         new_AGEMA_signal_5474, new_AGEMA_signal_5478, new_AGEMA_signal_5482,
         new_AGEMA_signal_5486, new_AGEMA_signal_5490, new_AGEMA_signal_5494,
         new_AGEMA_signal_5498, new_AGEMA_signal_5502, new_AGEMA_signal_5506,
         new_AGEMA_signal_5510, new_AGEMA_signal_5514, new_AGEMA_signal_5518,
         new_AGEMA_signal_5522, new_AGEMA_signal_5526, new_AGEMA_signal_5530,
         new_AGEMA_signal_5534, new_AGEMA_signal_5538, new_AGEMA_signal_5542,
         new_AGEMA_signal_5546, new_AGEMA_signal_5550, new_AGEMA_signal_5554,
         new_AGEMA_signal_5558, new_AGEMA_signal_5562, new_AGEMA_signal_5566,
         new_AGEMA_signal_5570, new_AGEMA_signal_5574, new_AGEMA_signal_5578,
         new_AGEMA_signal_5582, new_AGEMA_signal_5586, new_AGEMA_signal_5590,
         new_AGEMA_signal_5594, new_AGEMA_signal_5598, new_AGEMA_signal_5602,
         new_AGEMA_signal_5606, new_AGEMA_signal_5610, new_AGEMA_signal_5614,
         new_AGEMA_signal_5618, new_AGEMA_signal_5622, new_AGEMA_signal_5626,
         new_AGEMA_signal_5630, new_AGEMA_signal_5634, new_AGEMA_signal_5638,
         new_AGEMA_signal_5642, new_AGEMA_signal_5646, new_AGEMA_signal_5650,
         new_AGEMA_signal_5654, new_AGEMA_signal_5658, new_AGEMA_signal_5662,
         new_AGEMA_signal_5666, new_AGEMA_signal_5670, new_AGEMA_signal_5674,
         new_AGEMA_signal_5678, new_AGEMA_signal_5682, new_AGEMA_signal_5686,
         new_AGEMA_signal_5690, new_AGEMA_signal_5694, new_AGEMA_signal_5698,
         new_AGEMA_signal_5702, new_AGEMA_signal_5706, new_AGEMA_signal_5710,
         new_AGEMA_signal_5714, new_AGEMA_signal_5718, new_AGEMA_signal_5722,
         new_AGEMA_signal_5726, new_AGEMA_signal_5730, new_AGEMA_signal_5734,
         new_AGEMA_signal_5738, new_AGEMA_signal_5742, new_AGEMA_signal_5746,
         new_AGEMA_signal_5750, new_AGEMA_signal_5754, new_AGEMA_signal_5758,
         new_AGEMA_signal_5762, new_AGEMA_signal_5766, new_AGEMA_signal_5770,
         new_AGEMA_signal_5774, new_AGEMA_signal_5778, new_AGEMA_signal_5782,
         new_AGEMA_signal_5786, new_AGEMA_signal_5790, new_AGEMA_signal_5794,
         new_AGEMA_signal_5798, new_AGEMA_signal_5802, new_AGEMA_signal_5806,
         new_AGEMA_signal_5810, new_AGEMA_signal_5814, new_AGEMA_signal_5818,
         new_AGEMA_signal_5822, new_AGEMA_signal_5826, new_AGEMA_signal_5830,
         new_AGEMA_signal_5834, new_AGEMA_signal_5838, new_AGEMA_signal_5842,
         new_AGEMA_signal_5846, new_AGEMA_signal_5850, new_AGEMA_signal_5854,
         new_AGEMA_signal_5858, new_AGEMA_signal_5862, new_AGEMA_signal_5866,
         new_AGEMA_signal_5870, new_AGEMA_signal_5874, new_AGEMA_signal_5878,
         new_AGEMA_signal_5882, new_AGEMA_signal_5886, new_AGEMA_signal_5890,
         new_AGEMA_signal_5894, new_AGEMA_signal_5898, new_AGEMA_signal_5902,
         new_AGEMA_signal_5906, new_AGEMA_signal_5910, new_AGEMA_signal_5914,
         new_AGEMA_signal_5918, new_AGEMA_signal_5922, new_AGEMA_signal_5926,
         new_AGEMA_signal_5930, new_AGEMA_signal_5934, new_AGEMA_signal_5938,
         new_AGEMA_signal_5942, new_AGEMA_signal_5946, new_AGEMA_signal_5950,
         new_AGEMA_signal_5954, new_AGEMA_signal_5958, new_AGEMA_signal_5962,
         new_AGEMA_signal_5966, new_AGEMA_signal_5970, new_AGEMA_signal_5974,
         new_AGEMA_signal_5978, new_AGEMA_signal_5982, new_AGEMA_signal_5986,
         new_AGEMA_signal_5990, new_AGEMA_signal_5994, new_AGEMA_signal_5998,
         new_AGEMA_signal_6002, new_AGEMA_signal_6006, new_AGEMA_signal_6010,
         new_AGEMA_signal_6014, new_AGEMA_signal_6018, new_AGEMA_signal_6022,
         new_AGEMA_signal_6026, new_AGEMA_signal_6030, new_AGEMA_signal_6034,
         new_AGEMA_signal_6038, new_AGEMA_signal_6042, new_AGEMA_signal_6046,
         new_AGEMA_signal_6050, new_AGEMA_signal_6054, new_AGEMA_signal_6058,
         new_AGEMA_signal_6062, new_AGEMA_signal_6066, new_AGEMA_signal_6070,
         new_AGEMA_signal_6074, new_AGEMA_signal_6078, new_AGEMA_signal_6082,
         new_AGEMA_signal_6086, new_AGEMA_signal_6090, new_AGEMA_signal_6094,
         new_AGEMA_signal_6098, new_AGEMA_signal_6102, new_AGEMA_signal_6106,
         new_AGEMA_signal_3279, new_AGEMA_signal_2681, new_AGEMA_signal_2680,
         new_AGEMA_signal_3285, new_AGEMA_signal_3283, new_AGEMA_signal_3281,
         new_AGEMA_signal_2667, new_AGEMA_signal_2666, new_AGEMA_signal_2801,
         new_AGEMA_signal_2800, new_AGEMA_signal_3291, new_AGEMA_signal_3289,
         new_AGEMA_signal_3287, new_AGEMA_signal_2787, new_AGEMA_signal_2786,
         new_AGEMA_signal_2685, new_AGEMA_signal_2684, new_AGEMA_signal_3297,
         new_AGEMA_signal_3295, new_AGEMA_signal_3293, new_AGEMA_signal_2671,
         new_AGEMA_signal_2670, new_AGEMA_signal_2805, new_AGEMA_signal_2804,
         new_AGEMA_signal_3303, new_AGEMA_signal_3301, new_AGEMA_signal_3299,
         new_AGEMA_signal_2791, new_AGEMA_signal_2790, new_AGEMA_signal_2689,
         new_AGEMA_signal_2688, new_AGEMA_signal_3309, new_AGEMA_signal_3307,
         new_AGEMA_signal_3305, new_AGEMA_signal_2675, new_AGEMA_signal_2674,
         new_AGEMA_signal_2809, new_AGEMA_signal_2808, new_AGEMA_signal_3315,
         new_AGEMA_signal_3313, new_AGEMA_signal_3311, new_AGEMA_signal_2795,
         new_AGEMA_signal_2794, new_AGEMA_signal_2921, new_AGEMA_signal_2920,
         new_AGEMA_signal_3321, new_AGEMA_signal_3319, new_AGEMA_signal_3317,
         new_AGEMA_signal_2903, new_AGEMA_signal_2902, new_AGEMA_signal_3007,
         new_AGEMA_signal_3006, new_AGEMA_signal_3327, new_AGEMA_signal_3325,
         new_AGEMA_signal_3323, new_AGEMA_signal_2991, new_AGEMA_signal_2990,
         new_AGEMA_signal_2693, new_AGEMA_signal_2692, new_AGEMA_signal_3333,
         new_AGEMA_signal_3331, new_AGEMA_signal_3329, new_AGEMA_signal_2655,
         new_AGEMA_signal_2654, new_AGEMA_signal_2813, new_AGEMA_signal_2812,
         new_AGEMA_signal_3339, new_AGEMA_signal_3337, new_AGEMA_signal_3335,
         new_AGEMA_signal_2773, new_AGEMA_signal_2772, new_AGEMA_signal_2697,
         new_AGEMA_signal_2696, new_AGEMA_signal_3345, new_AGEMA_signal_3343,
         new_AGEMA_signal_3341, new_AGEMA_signal_2659, new_AGEMA_signal_2658,
         new_AGEMA_signal_2817, new_AGEMA_signal_2816, new_AGEMA_signal_3351,
         new_AGEMA_signal_3349, new_AGEMA_signal_3347, new_AGEMA_signal_2777,
         new_AGEMA_signal_2776, new_AGEMA_signal_2933, new_AGEMA_signal_2932,
         new_AGEMA_signal_3357, new_AGEMA_signal_3355, new_AGEMA_signal_3353,
         new_AGEMA_signal_2883, new_AGEMA_signal_2882, new_AGEMA_signal_3019,
         new_AGEMA_signal_3018, new_AGEMA_signal_3363, new_AGEMA_signal_3361,
         new_AGEMA_signal_3359, new_AGEMA_signal_2979, new_AGEMA_signal_2978,
         new_AGEMA_signal_2701, new_AGEMA_signal_2700, new_AGEMA_signal_3369,
         new_AGEMA_signal_3367, new_AGEMA_signal_3365, new_AGEMA_signal_2663,
         new_AGEMA_signal_2662, new_AGEMA_signal_2821, new_AGEMA_signal_2820,
         new_AGEMA_signal_3375, new_AGEMA_signal_3373, new_AGEMA_signal_3371,
         new_AGEMA_signal_2783, new_AGEMA_signal_2782, new_AGEMA_signal_2479,
         new_AGEMA_signal_2478, new_AGEMA_signal_3381, new_AGEMA_signal_3379,
         new_AGEMA_signal_3377, new_AGEMA_signal_2457, new_AGEMA_signal_2456,
         new_AGEMA_signal_2585, new_AGEMA_signal_2584, new_AGEMA_signal_3387,
         new_AGEMA_signal_3385, new_AGEMA_signal_3383, new_AGEMA_signal_2545,
         new_AGEMA_signal_2544, new_AGEMA_signal_2483, new_AGEMA_signal_2482,
         new_AGEMA_signal_3393, new_AGEMA_signal_3391, new_AGEMA_signal_3389,
         new_AGEMA_signal_2461, new_AGEMA_signal_2460, new_AGEMA_signal_2589,
         new_AGEMA_signal_2588, new_AGEMA_signal_3399, new_AGEMA_signal_3397,
         new_AGEMA_signal_3395, new_AGEMA_signal_2549, new_AGEMA_signal_2548,
         new_AGEMA_signal_2487, new_AGEMA_signal_2486, new_AGEMA_signal_3405,
         new_AGEMA_signal_3403, new_AGEMA_signal_3401, new_AGEMA_signal_2465,
         new_AGEMA_signal_2464, new_AGEMA_signal_2593, new_AGEMA_signal_2592,
         new_AGEMA_signal_3411, new_AGEMA_signal_3409, new_AGEMA_signal_3407,
         new_AGEMA_signal_2553, new_AGEMA_signal_2552, new_AGEMA_signal_2717,
         new_AGEMA_signal_2716, new_AGEMA_signal_3417, new_AGEMA_signal_3415,
         new_AGEMA_signal_3413, new_AGEMA_signal_2633, new_AGEMA_signal_2632,
         new_AGEMA_signal_2837, new_AGEMA_signal_2836, new_AGEMA_signal_3423,
         new_AGEMA_signal_3421, new_AGEMA_signal_3419, new_AGEMA_signal_2753,
         new_AGEMA_signal_2752, new_AGEMA_signal_2721, new_AGEMA_signal_2720,
         new_AGEMA_signal_3429, new_AGEMA_signal_3427, new_AGEMA_signal_3425,
         new_AGEMA_signal_2639, new_AGEMA_signal_2638, new_AGEMA_signal_2841,
         new_AGEMA_signal_2840, new_AGEMA_signal_3435, new_AGEMA_signal_3433,
         new_AGEMA_signal_3431, new_AGEMA_signal_2757, new_AGEMA_signal_2756,
         new_AGEMA_signal_2725, new_AGEMA_signal_2724, new_AGEMA_signal_3441,
         new_AGEMA_signal_3439, new_AGEMA_signal_3437, new_AGEMA_signal_2643,
         new_AGEMA_signal_2642, new_AGEMA_signal_2845, new_AGEMA_signal_2844,
         new_AGEMA_signal_3447, new_AGEMA_signal_3445, new_AGEMA_signal_3443,
         new_AGEMA_signal_2763, new_AGEMA_signal_2762, new_AGEMA_signal_2729,
         new_AGEMA_signal_2728, new_AGEMA_signal_3453, new_AGEMA_signal_3451,
         new_AGEMA_signal_3449, new_AGEMA_signal_2649, new_AGEMA_signal_2648,
         new_AGEMA_signal_2849, new_AGEMA_signal_2848, new_AGEMA_signal_3459,
         new_AGEMA_signal_3457, new_AGEMA_signal_3455, new_AGEMA_signal_2767,
         new_AGEMA_signal_2766, new_AGEMA_signal_2957, new_AGEMA_signal_2956,
         new_AGEMA_signal_3465, new_AGEMA_signal_3463, new_AGEMA_signal_3461,
         new_AGEMA_signal_2871, new_AGEMA_signal_2870, new_AGEMA_signal_3043,
         new_AGEMA_signal_3042, new_AGEMA_signal_3471, new_AGEMA_signal_3469,
         new_AGEMA_signal_3467, new_AGEMA_signal_2971, new_AGEMA_signal_2970,
         new_AGEMA_signal_2285, new_AGEMA_signal_2284,
         SubCellInst_SboxInst_0_YY_1_, new_AGEMA_signal_2157,
         new_AGEMA_signal_2156, SubCellInst_SboxInst_0_YY_0_,
         new_AGEMA_signal_1933, new_AGEMA_signal_1932,
         SubCellInst_SboxInst_0_T0, new_AGEMA_signal_2029,
         new_AGEMA_signal_2028, SubCellInst_SboxInst_0_Q2,
         new_AGEMA_signal_3477, new_AGEMA_signal_3475, new_AGEMA_signal_3473,
         new_AGEMA_signal_1935, new_AGEMA_signal_1934,
         SubCellInst_SboxInst_0_T2, new_AGEMA_signal_2031,
         new_AGEMA_signal_2030, SubCellInst_SboxInst_0_Q7,
         new_AGEMA_signal_3483, new_AGEMA_signal_3481, new_AGEMA_signal_3479,
         new_AGEMA_signal_2033, new_AGEMA_signal_2032,
         SubCellInst_SboxInst_0_L3, new_AGEMA_signal_3489,
         new_AGEMA_signal_3487, new_AGEMA_signal_3485, new_AGEMA_signal_3495,
         new_AGEMA_signal_3493, new_AGEMA_signal_3491, new_AGEMA_signal_2289,
         new_AGEMA_signal_2288, SubCellInst_SboxInst_1_YY_1_,
         new_AGEMA_signal_2165, new_AGEMA_signal_2164,
         SubCellInst_SboxInst_1_YY_0_, new_AGEMA_signal_1939,
         new_AGEMA_signal_1938, SubCellInst_SboxInst_1_T0,
         new_AGEMA_signal_2037, new_AGEMA_signal_2036,
         SubCellInst_SboxInst_1_Q2, new_AGEMA_signal_3501,
         new_AGEMA_signal_3499, new_AGEMA_signal_3497, new_AGEMA_signal_1941,
         new_AGEMA_signal_1940, SubCellInst_SboxInst_1_T2,
         new_AGEMA_signal_2039, new_AGEMA_signal_2038,
         SubCellInst_SboxInst_1_Q7, new_AGEMA_signal_3507,
         new_AGEMA_signal_3505, new_AGEMA_signal_3503, new_AGEMA_signal_2041,
         new_AGEMA_signal_2040, SubCellInst_SboxInst_1_L3,
         new_AGEMA_signal_3513, new_AGEMA_signal_3511, new_AGEMA_signal_3509,
         new_AGEMA_signal_3519, new_AGEMA_signal_3517, new_AGEMA_signal_3515,
         new_AGEMA_signal_2293, new_AGEMA_signal_2292,
         SubCellInst_SboxInst_2_YY_1_, new_AGEMA_signal_2173,
         new_AGEMA_signal_2172, SubCellInst_SboxInst_2_YY_0_,
         new_AGEMA_signal_1945, new_AGEMA_signal_1944,
         SubCellInst_SboxInst_2_T0, new_AGEMA_signal_2045,
         new_AGEMA_signal_2044, SubCellInst_SboxInst_2_Q2,
         new_AGEMA_signal_3525, new_AGEMA_signal_3523, new_AGEMA_signal_3521,
         new_AGEMA_signal_1947, new_AGEMA_signal_1946,
         SubCellInst_SboxInst_2_T2, new_AGEMA_signal_2047,
         new_AGEMA_signal_2046, SubCellInst_SboxInst_2_Q7,
         new_AGEMA_signal_3531, new_AGEMA_signal_3529, new_AGEMA_signal_3527,
         new_AGEMA_signal_2049, new_AGEMA_signal_2048,
         SubCellInst_SboxInst_2_L3, new_AGEMA_signal_3537,
         new_AGEMA_signal_3535, new_AGEMA_signal_3533, new_AGEMA_signal_3543,
         new_AGEMA_signal_3541, new_AGEMA_signal_3539, new_AGEMA_signal_2297,
         new_AGEMA_signal_2296, SubCellInst_SboxInst_3_YY_1_,
         new_AGEMA_signal_2181, new_AGEMA_signal_2180,
         SubCellInst_SboxInst_3_YY_0_, new_AGEMA_signal_1951,
         new_AGEMA_signal_1950, SubCellInst_SboxInst_3_T0,
         new_AGEMA_signal_2053, new_AGEMA_signal_2052,
         SubCellInst_SboxInst_3_Q2, new_AGEMA_signal_3549,
         new_AGEMA_signal_3547, new_AGEMA_signal_3545, new_AGEMA_signal_1953,
         new_AGEMA_signal_1952, SubCellInst_SboxInst_3_T2,
         new_AGEMA_signal_2055, new_AGEMA_signal_2054,
         SubCellInst_SboxInst_3_Q7, new_AGEMA_signal_3555,
         new_AGEMA_signal_3553, new_AGEMA_signal_3551, new_AGEMA_signal_2057,
         new_AGEMA_signal_2056, SubCellInst_SboxInst_3_L3,
         new_AGEMA_signal_3561, new_AGEMA_signal_3559, new_AGEMA_signal_3557,
         new_AGEMA_signal_3567, new_AGEMA_signal_3565, new_AGEMA_signal_3563,
         new_AGEMA_signal_2301, new_AGEMA_signal_2300,
         SubCellInst_SboxInst_4_YY_1_, new_AGEMA_signal_2189,
         new_AGEMA_signal_2188, SubCellInst_SboxInst_4_YY_0_,
         new_AGEMA_signal_1957, new_AGEMA_signal_1956,
         SubCellInst_SboxInst_4_T0, new_AGEMA_signal_2061,
         new_AGEMA_signal_2060, SubCellInst_SboxInst_4_Q2,
         new_AGEMA_signal_3573, new_AGEMA_signal_3571, new_AGEMA_signal_3569,
         new_AGEMA_signal_1959, new_AGEMA_signal_1958,
         SubCellInst_SboxInst_4_T2, new_AGEMA_signal_2063,
         new_AGEMA_signal_2062, SubCellInst_SboxInst_4_Q7,
         new_AGEMA_signal_3579, new_AGEMA_signal_3577, new_AGEMA_signal_3575,
         new_AGEMA_signal_2065, new_AGEMA_signal_2064,
         SubCellInst_SboxInst_4_L3, new_AGEMA_signal_3585,
         new_AGEMA_signal_3583, new_AGEMA_signal_3581, new_AGEMA_signal_3591,
         new_AGEMA_signal_3589, new_AGEMA_signal_3587, new_AGEMA_signal_2305,
         new_AGEMA_signal_2304, SubCellInst_SboxInst_5_YY_1_,
         new_AGEMA_signal_2197, new_AGEMA_signal_2196,
         SubCellInst_SboxInst_5_YY_0_, new_AGEMA_signal_1963,
         new_AGEMA_signal_1962, SubCellInst_SboxInst_5_T0,
         new_AGEMA_signal_2069, new_AGEMA_signal_2068,
         SubCellInst_SboxInst_5_Q2, new_AGEMA_signal_3597,
         new_AGEMA_signal_3595, new_AGEMA_signal_3593, new_AGEMA_signal_1965,
         new_AGEMA_signal_1964, SubCellInst_SboxInst_5_T2,
         new_AGEMA_signal_2071, new_AGEMA_signal_2070,
         SubCellInst_SboxInst_5_Q7, new_AGEMA_signal_3603,
         new_AGEMA_signal_3601, new_AGEMA_signal_3599, new_AGEMA_signal_2073,
         new_AGEMA_signal_2072, SubCellInst_SboxInst_5_L3,
         new_AGEMA_signal_3609, new_AGEMA_signal_3607, new_AGEMA_signal_3605,
         new_AGEMA_signal_3615, new_AGEMA_signal_3613, new_AGEMA_signal_3611,
         new_AGEMA_signal_2309, new_AGEMA_signal_2308,
         SubCellInst_SboxInst_6_YY_1_, new_AGEMA_signal_2205,
         new_AGEMA_signal_2204, SubCellInst_SboxInst_6_YY_0_,
         new_AGEMA_signal_1969, new_AGEMA_signal_1968,
         SubCellInst_SboxInst_6_T0, new_AGEMA_signal_2077,
         new_AGEMA_signal_2076, SubCellInst_SboxInst_6_Q2,
         new_AGEMA_signal_3621, new_AGEMA_signal_3619, new_AGEMA_signal_3617,
         new_AGEMA_signal_1971, new_AGEMA_signal_1970,
         SubCellInst_SboxInst_6_T2, new_AGEMA_signal_2079,
         new_AGEMA_signal_2078, SubCellInst_SboxInst_6_Q7,
         new_AGEMA_signal_3627, new_AGEMA_signal_3625, new_AGEMA_signal_3623,
         new_AGEMA_signal_2081, new_AGEMA_signal_2080,
         SubCellInst_SboxInst_6_L3, new_AGEMA_signal_3633,
         new_AGEMA_signal_3631, new_AGEMA_signal_3629, new_AGEMA_signal_3639,
         new_AGEMA_signal_3637, new_AGEMA_signal_3635, new_AGEMA_signal_2313,
         new_AGEMA_signal_2312, SubCellInst_SboxInst_7_YY_1_,
         new_AGEMA_signal_2213, new_AGEMA_signal_2212,
         SubCellInst_SboxInst_7_YY_0_, new_AGEMA_signal_1975,
         new_AGEMA_signal_1974, SubCellInst_SboxInst_7_T0,
         new_AGEMA_signal_2085, new_AGEMA_signal_2084,
         SubCellInst_SboxInst_7_Q2, new_AGEMA_signal_3645,
         new_AGEMA_signal_3643, new_AGEMA_signal_3641, new_AGEMA_signal_1977,
         new_AGEMA_signal_1976, SubCellInst_SboxInst_7_T2,
         new_AGEMA_signal_2087, new_AGEMA_signal_2086,
         SubCellInst_SboxInst_7_Q7, new_AGEMA_signal_3651,
         new_AGEMA_signal_3649, new_AGEMA_signal_3647, new_AGEMA_signal_2089,
         new_AGEMA_signal_2088, SubCellInst_SboxInst_7_L3,
         new_AGEMA_signal_3657, new_AGEMA_signal_3655, new_AGEMA_signal_3653,
         new_AGEMA_signal_3663, new_AGEMA_signal_3661, new_AGEMA_signal_3659,
         new_AGEMA_signal_2317, new_AGEMA_signal_2316,
         SubCellInst_SboxInst_8_YY_1_, new_AGEMA_signal_2221,
         new_AGEMA_signal_2220, SubCellInst_SboxInst_8_YY_0_,
         new_AGEMA_signal_1981, new_AGEMA_signal_1980,
         SubCellInst_SboxInst_8_T0, new_AGEMA_signal_2093,
         new_AGEMA_signal_2092, SubCellInst_SboxInst_8_Q2,
         new_AGEMA_signal_3669, new_AGEMA_signal_3667, new_AGEMA_signal_3665,
         new_AGEMA_signal_1983, new_AGEMA_signal_1982,
         SubCellInst_SboxInst_8_T2, new_AGEMA_signal_2095,
         new_AGEMA_signal_2094, SubCellInst_SboxInst_8_Q7,
         new_AGEMA_signal_3675, new_AGEMA_signal_3673, new_AGEMA_signal_3671,
         new_AGEMA_signal_2097, new_AGEMA_signal_2096,
         SubCellInst_SboxInst_8_L3, new_AGEMA_signal_3681,
         new_AGEMA_signal_3679, new_AGEMA_signal_3677, new_AGEMA_signal_3687,
         new_AGEMA_signal_3685, new_AGEMA_signal_3683, new_AGEMA_signal_2321,
         new_AGEMA_signal_2320, SubCellInst_SboxInst_9_YY_1_,
         new_AGEMA_signal_2229, new_AGEMA_signal_2228,
         SubCellInst_SboxInst_9_YY_0_, new_AGEMA_signal_1987,
         new_AGEMA_signal_1986, SubCellInst_SboxInst_9_T0,
         new_AGEMA_signal_2101, new_AGEMA_signal_2100,
         SubCellInst_SboxInst_9_Q2, new_AGEMA_signal_3693,
         new_AGEMA_signal_3691, new_AGEMA_signal_3689, new_AGEMA_signal_1989,
         new_AGEMA_signal_1988, SubCellInst_SboxInst_9_T2,
         new_AGEMA_signal_2103, new_AGEMA_signal_2102,
         SubCellInst_SboxInst_9_Q7, new_AGEMA_signal_3699,
         new_AGEMA_signal_3697, new_AGEMA_signal_3695, new_AGEMA_signal_2105,
         new_AGEMA_signal_2104, SubCellInst_SboxInst_9_L3,
         new_AGEMA_signal_3705, new_AGEMA_signal_3703, new_AGEMA_signal_3701,
         new_AGEMA_signal_3711, new_AGEMA_signal_3709, new_AGEMA_signal_3707,
         new_AGEMA_signal_2325, new_AGEMA_signal_2324,
         SubCellInst_SboxInst_10_YY_1_, new_AGEMA_signal_2237,
         new_AGEMA_signal_2236, SubCellInst_SboxInst_10_YY_0_,
         new_AGEMA_signal_1993, new_AGEMA_signal_1992,
         SubCellInst_SboxInst_10_T0, new_AGEMA_signal_2109,
         new_AGEMA_signal_2108, SubCellInst_SboxInst_10_Q2,
         new_AGEMA_signal_3717, new_AGEMA_signal_3715, new_AGEMA_signal_3713,
         new_AGEMA_signal_1995, new_AGEMA_signal_1994,
         SubCellInst_SboxInst_10_T2, new_AGEMA_signal_2111,
         new_AGEMA_signal_2110, SubCellInst_SboxInst_10_Q7,
         new_AGEMA_signal_3723, new_AGEMA_signal_3721, new_AGEMA_signal_3719,
         new_AGEMA_signal_2113, new_AGEMA_signal_2112,
         SubCellInst_SboxInst_10_L3, new_AGEMA_signal_3729,
         new_AGEMA_signal_3727, new_AGEMA_signal_3725, new_AGEMA_signal_3735,
         new_AGEMA_signal_3733, new_AGEMA_signal_3731, SubCellOutput_47,
         SubCellOutput_46, SubCellOutput_45, SubCellOutput_44,
         SubCellOutput_29, new_AGEMA_signal_2329, new_AGEMA_signal_2328,
         SubCellInst_SboxInst_11_YY_1_, new_AGEMA_signal_2245,
         new_AGEMA_signal_2244, SubCellInst_SboxInst_11_YY_0_,
         new_AGEMA_signal_1999, new_AGEMA_signal_1998,
         SubCellInst_SboxInst_11_T0, new_AGEMA_signal_2117,
         new_AGEMA_signal_2116, SubCellInst_SboxInst_11_Q2,
         new_AGEMA_signal_3741, new_AGEMA_signal_3739, new_AGEMA_signal_3737,
         new_AGEMA_signal_2001, new_AGEMA_signal_2000,
         SubCellInst_SboxInst_11_T2, new_AGEMA_signal_2119,
         new_AGEMA_signal_2118, SubCellInst_SboxInst_11_Q7,
         new_AGEMA_signal_3747, new_AGEMA_signal_3745, new_AGEMA_signal_3743,
         new_AGEMA_signal_2121, new_AGEMA_signal_2120,
         SubCellInst_SboxInst_11_L3, new_AGEMA_signal_3753,
         new_AGEMA_signal_3751, new_AGEMA_signal_3749, new_AGEMA_signal_3759,
         new_AGEMA_signal_3757, new_AGEMA_signal_3755, new_AGEMA_signal_2333,
         new_AGEMA_signal_2332, SubCellInst_SboxInst_12_YY_1_,
         new_AGEMA_signal_2253, new_AGEMA_signal_2252,
         SubCellInst_SboxInst_12_YY_0_, new_AGEMA_signal_2005,
         new_AGEMA_signal_2004, SubCellInst_SboxInst_12_T0,
         new_AGEMA_signal_2125, new_AGEMA_signal_2124,
         SubCellInst_SboxInst_12_Q2, new_AGEMA_signal_3765,
         new_AGEMA_signal_3763, new_AGEMA_signal_3761, new_AGEMA_signal_2007,
         new_AGEMA_signal_2006, SubCellInst_SboxInst_12_T2,
         new_AGEMA_signal_2127, new_AGEMA_signal_2126,
         SubCellInst_SboxInst_12_Q7, new_AGEMA_signal_3771,
         new_AGEMA_signal_3769, new_AGEMA_signal_3767, new_AGEMA_signal_2129,
         new_AGEMA_signal_2128, SubCellInst_SboxInst_12_L3,
         new_AGEMA_signal_3777, new_AGEMA_signal_3775, new_AGEMA_signal_3773,
         new_AGEMA_signal_3783, new_AGEMA_signal_3781, new_AGEMA_signal_3779,
         new_AGEMA_signal_2337, new_AGEMA_signal_2336,
         SubCellInst_SboxInst_13_YY_1_, new_AGEMA_signal_2261,
         new_AGEMA_signal_2260, SubCellInst_SboxInst_13_YY_0_,
         new_AGEMA_signal_2011, new_AGEMA_signal_2010,
         SubCellInst_SboxInst_13_T0, new_AGEMA_signal_2133,
         new_AGEMA_signal_2132, SubCellInst_SboxInst_13_Q2,
         new_AGEMA_signal_3789, new_AGEMA_signal_3787, new_AGEMA_signal_3785,
         new_AGEMA_signal_2013, new_AGEMA_signal_2012,
         SubCellInst_SboxInst_13_T2, new_AGEMA_signal_2135,
         new_AGEMA_signal_2134, SubCellInst_SboxInst_13_Q7,
         new_AGEMA_signal_3795, new_AGEMA_signal_3793, new_AGEMA_signal_3791,
         new_AGEMA_signal_2137, new_AGEMA_signal_2136,
         SubCellInst_SboxInst_13_L3, new_AGEMA_signal_3801,
         new_AGEMA_signal_3799, new_AGEMA_signal_3797, new_AGEMA_signal_3807,
         new_AGEMA_signal_3805, new_AGEMA_signal_3803, new_AGEMA_signal_2341,
         new_AGEMA_signal_2340, SubCellInst_SboxInst_14_YY_1_,
         new_AGEMA_signal_2269, new_AGEMA_signal_2268,
         SubCellInst_SboxInst_14_YY_0_, new_AGEMA_signal_2017,
         new_AGEMA_signal_2016, SubCellInst_SboxInst_14_T0,
         new_AGEMA_signal_2141, new_AGEMA_signal_2140,
         SubCellInst_SboxInst_14_Q2, new_AGEMA_signal_3813,
         new_AGEMA_signal_3811, new_AGEMA_signal_3809, new_AGEMA_signal_2019,
         new_AGEMA_signal_2018, SubCellInst_SboxInst_14_T2,
         new_AGEMA_signal_2143, new_AGEMA_signal_2142,
         SubCellInst_SboxInst_14_Q7, new_AGEMA_signal_3819,
         new_AGEMA_signal_3817, new_AGEMA_signal_3815, new_AGEMA_signal_2145,
         new_AGEMA_signal_2144, SubCellInst_SboxInst_14_L3,
         new_AGEMA_signal_3825, new_AGEMA_signal_3823, new_AGEMA_signal_3821,
         new_AGEMA_signal_3831, new_AGEMA_signal_3829, new_AGEMA_signal_3827,
         new_AGEMA_signal_2345, new_AGEMA_signal_2344,
         SubCellInst_SboxInst_15_YY_1_, new_AGEMA_signal_2277,
         new_AGEMA_signal_2276, SubCellInst_SboxInst_15_YY_0_,
         new_AGEMA_signal_2023, new_AGEMA_signal_2022,
         SubCellInst_SboxInst_15_T0, new_AGEMA_signal_2149,
         new_AGEMA_signal_2148, SubCellInst_SboxInst_15_Q2,
         new_AGEMA_signal_3837, new_AGEMA_signal_3835, new_AGEMA_signal_3833,
         new_AGEMA_signal_2025, new_AGEMA_signal_2024,
         SubCellInst_SboxInst_15_T2, new_AGEMA_signal_2151,
         new_AGEMA_signal_2150, SubCellInst_SboxInst_15_Q7,
         new_AGEMA_signal_3843, new_AGEMA_signal_3841, new_AGEMA_signal_3839,
         new_AGEMA_signal_2153, new_AGEMA_signal_2152,
         SubCellInst_SboxInst_15_L3, new_AGEMA_signal_3849,
         new_AGEMA_signal_3847, new_AGEMA_signal_3845, new_AGEMA_signal_3855,
         new_AGEMA_signal_3853, new_AGEMA_signal_3851, new_AGEMA_signal_2437,
         new_AGEMA_signal_2436, new_AGEMA_signal_3857, new_AGEMA_signal_2349,
         new_AGEMA_signal_2348, AddConstXOR_AddConstXOR_XORInst_0_2_n1,
         new_AGEMA_signal_2523, new_AGEMA_signal_2522, new_AGEMA_signal_3859,
         new_AGEMA_signal_2439, new_AGEMA_signal_2438,
         AddConstXOR_AddConstXOR_XORInst_0_3_n1, new_AGEMA_signal_2441,
         new_AGEMA_signal_2440, new_AGEMA_signal_2351, new_AGEMA_signal_2350,
         AddConstXOR_AddConstXOR_XORInst_1_2_n1, new_AGEMA_signal_2527,
         new_AGEMA_signal_2526, new_AGEMA_signal_2443, new_AGEMA_signal_2442,
         AddConstXOR_AddConstXOR_XORInst_1_3_n1, new_AGEMA_signal_2445,
         new_AGEMA_signal_2444, new_AGEMA_signal_3865, new_AGEMA_signal_3863,
         new_AGEMA_signal_3861, new_AGEMA_signal_2353, new_AGEMA_signal_2352,
         AddRoundTweakeyXOR_XORInst_0_2_n1, new_AGEMA_signal_2531,
         new_AGEMA_signal_2530, new_AGEMA_signal_3871, new_AGEMA_signal_3869,
         new_AGEMA_signal_3867, new_AGEMA_signal_2447, new_AGEMA_signal_2446,
         AddRoundTweakeyXOR_XORInst_0_3_n1, new_AGEMA_signal_2449,
         new_AGEMA_signal_2448, new_AGEMA_signal_3877, new_AGEMA_signal_3875,
         new_AGEMA_signal_3873, new_AGEMA_signal_2355, new_AGEMA_signal_2354,
         AddRoundTweakeyXOR_XORInst_1_2_n1, new_AGEMA_signal_2535,
         new_AGEMA_signal_2534, new_AGEMA_signal_3883, new_AGEMA_signal_3881,
         new_AGEMA_signal_3879, new_AGEMA_signal_2451, new_AGEMA_signal_2450,
         AddRoundTweakeyXOR_XORInst_1_3_n1, new_AGEMA_signal_2453,
         new_AGEMA_signal_2452, new_AGEMA_signal_3889, new_AGEMA_signal_3887,
         new_AGEMA_signal_3885, new_AGEMA_signal_2357, new_AGEMA_signal_2356,
         AddRoundTweakeyXOR_XORInst_2_2_n1, new_AGEMA_signal_2539,
         new_AGEMA_signal_2538, new_AGEMA_signal_3895, new_AGEMA_signal_3893,
         new_AGEMA_signal_3891, new_AGEMA_signal_2455, new_AGEMA_signal_2454,
         AddRoundTweakeyXOR_XORInst_2_3_n1, new_AGEMA_signal_2617,
         new_AGEMA_signal_2616, new_AGEMA_signal_3901, new_AGEMA_signal_3899,
         new_AGEMA_signal_3897, new_AGEMA_signal_2541, new_AGEMA_signal_2540,
         AddRoundTweakeyXOR_XORInst_3_2_n1, new_AGEMA_signal_2743,
         new_AGEMA_signal_2742, new_AGEMA_signal_3907, new_AGEMA_signal_3905,
         new_AGEMA_signal_3903, new_AGEMA_signal_2619, new_AGEMA_signal_2618,
         AddRoundTweakeyXOR_XORInst_3_3_n1, new_AGEMA_signal_3913,
         new_AGEMA_signal_3911, new_AGEMA_signal_3909, new_AGEMA_signal_2359,
         new_AGEMA_signal_2358, AddRoundTweakeyXOR_XORInst_4_2_n1,
         new_AGEMA_signal_3919, new_AGEMA_signal_3917, new_AGEMA_signal_3915,
         new_AGEMA_signal_2459, new_AGEMA_signal_2458,
         AddRoundTweakeyXOR_XORInst_4_3_n1, new_AGEMA_signal_3925,
         new_AGEMA_signal_3923, new_AGEMA_signal_3921, new_AGEMA_signal_2361,
         new_AGEMA_signal_2360, AddRoundTweakeyXOR_XORInst_5_2_n1,
         new_AGEMA_signal_3931, new_AGEMA_signal_3929, new_AGEMA_signal_3927,
         new_AGEMA_signal_2463, new_AGEMA_signal_2462,
         AddRoundTweakeyXOR_XORInst_5_3_n1, new_AGEMA_signal_3937,
         new_AGEMA_signal_3935, new_AGEMA_signal_3933, new_AGEMA_signal_2363,
         new_AGEMA_signal_2362, AddRoundTweakeyXOR_XORInst_6_2_n1,
         new_AGEMA_signal_3943, new_AGEMA_signal_3941, new_AGEMA_signal_3939,
         new_AGEMA_signal_2467, new_AGEMA_signal_2466,
         AddRoundTweakeyXOR_XORInst_6_3_n1, new_AGEMA_signal_3949,
         new_AGEMA_signal_3947, new_AGEMA_signal_3945, new_AGEMA_signal_2555,
         new_AGEMA_signal_2554, AddRoundTweakeyXOR_XORInst_7_2_n1,
         new_AGEMA_signal_3955, new_AGEMA_signal_3953, new_AGEMA_signal_3951,
         new_AGEMA_signal_2635, new_AGEMA_signal_2634,
         AddRoundTweakeyXOR_XORInst_7_3_n1, new_AGEMA_signal_2365,
         new_AGEMA_signal_2364, MCInst_MCR0_XORInst_0_2_n1,
         new_AGEMA_signal_2559, new_AGEMA_signal_2558,
         MCInst_MCR0_XORInst_0_2_n2, new_AGEMA_signal_2469,
         new_AGEMA_signal_2468, MCInst_MCR0_XORInst_0_3_n1,
         new_AGEMA_signal_2641, new_AGEMA_signal_2640,
         MCInst_MCR0_XORInst_0_3_n2, new_AGEMA_signal_2367,
         new_AGEMA_signal_2366, MCInst_MCR0_XORInst_1_2_n1,
         new_AGEMA_signal_2563, new_AGEMA_signal_2562,
         MCInst_MCR0_XORInst_1_2_n2, new_AGEMA_signal_2471,
         new_AGEMA_signal_2470, MCInst_MCR0_XORInst_1_3_n1,
         new_AGEMA_signal_2645, new_AGEMA_signal_2644,
         MCInst_MCR0_XORInst_1_3_n2, new_AGEMA_signal_2369,
         new_AGEMA_signal_2368, MCInst_MCR0_XORInst_2_2_n1,
         new_AGEMA_signal_2567, new_AGEMA_signal_2566,
         MCInst_MCR0_XORInst_2_2_n2, new_AGEMA_signal_2473,
         new_AGEMA_signal_2472, MCInst_MCR0_XORInst_2_3_n1,
         new_AGEMA_signal_2651, new_AGEMA_signal_2650,
         MCInst_MCR0_XORInst_2_3_n2, new_AGEMA_signal_2371,
         new_AGEMA_signal_2370, MCInst_MCR0_XORInst_3_2_n1,
         new_AGEMA_signal_2769, new_AGEMA_signal_2768,
         MCInst_MCR0_XORInst_3_2_n2, new_AGEMA_signal_2475,
         new_AGEMA_signal_2474, MCInst_MCR0_XORInst_3_3_n1,
         new_AGEMA_signal_2873, new_AGEMA_signal_2872,
         MCInst_MCR0_XORInst_3_3_n2, new_AGEMA_signal_2571,
         new_AGEMA_signal_2570, MCInst_MCR2_XORInst_0_2_n1,
         new_AGEMA_signal_2657, new_AGEMA_signal_2656,
         MCInst_MCR2_XORInst_0_3_n1, new_AGEMA_signal_2573,
         new_AGEMA_signal_2572, MCInst_MCR2_XORInst_1_2_n1,
         new_AGEMA_signal_2661, new_AGEMA_signal_2660,
         MCInst_MCR2_XORInst_1_3_n1, new_AGEMA_signal_2779,
         new_AGEMA_signal_2778, MCInst_MCR2_XORInst_2_2_n1,
         new_AGEMA_signal_2885, new_AGEMA_signal_2884,
         MCInst_MCR2_XORInst_2_3_n1, new_AGEMA_signal_2575,
         new_AGEMA_signal_2574, MCInst_MCR2_XORInst_3_2_n1,
         new_AGEMA_signal_2665, new_AGEMA_signal_2664,
         MCInst_MCR2_XORInst_3_3_n1, new_AGEMA_signal_2577,
         new_AGEMA_signal_2576, MCInst_MCR3_XORInst_0_2_n1,
         new_AGEMA_signal_2669, new_AGEMA_signal_2668,
         MCInst_MCR3_XORInst_0_3_n1, new_AGEMA_signal_2579,
         new_AGEMA_signal_2578, MCInst_MCR3_XORInst_1_2_n1,
         new_AGEMA_signal_2673, new_AGEMA_signal_2672,
         MCInst_MCR3_XORInst_1_3_n1, new_AGEMA_signal_2581,
         new_AGEMA_signal_2580, MCInst_MCR3_XORInst_2_2_n1,
         new_AGEMA_signal_2677, new_AGEMA_signal_2676,
         MCInst_MCR3_XORInst_2_3_n1, new_AGEMA_signal_2797,
         new_AGEMA_signal_2796, MCInst_MCR3_XORInst_3_2_n1,
         new_AGEMA_signal_2905, new_AGEMA_signal_2904,
         MCInst_MCR3_XORInst_3_3_n1, new_AGEMA_signal_3959,
         new_AGEMA_signal_3963, new_AGEMA_signal_3967, new_AGEMA_signal_3971,
         new_AGEMA_signal_3975, new_AGEMA_signal_3979, new_AGEMA_signal_3983,
         new_AGEMA_signal_3987, new_AGEMA_signal_3991, new_AGEMA_signal_3995,
         new_AGEMA_signal_3999, new_AGEMA_signal_4003, new_AGEMA_signal_4007,
         new_AGEMA_signal_4011, new_AGEMA_signal_4015, new_AGEMA_signal_4019,
         new_AGEMA_signal_4023, new_AGEMA_signal_4027, new_AGEMA_signal_4031,
         new_AGEMA_signal_4035, new_AGEMA_signal_4039, new_AGEMA_signal_4043,
         new_AGEMA_signal_4047, new_AGEMA_signal_4051, new_AGEMA_signal_4055,
         new_AGEMA_signal_4059, new_AGEMA_signal_4063, new_AGEMA_signal_4067,
         new_AGEMA_signal_4071, new_AGEMA_signal_4075, new_AGEMA_signal_4079,
         new_AGEMA_signal_4083, new_AGEMA_signal_4087, new_AGEMA_signal_4091,
         new_AGEMA_signal_4095, new_AGEMA_signal_4099, new_AGEMA_signal_4103,
         new_AGEMA_signal_4107, new_AGEMA_signal_4111, new_AGEMA_signal_4115,
         new_AGEMA_signal_4119, new_AGEMA_signal_4123, new_AGEMA_signal_4127,
         new_AGEMA_signal_4131, new_AGEMA_signal_4135, new_AGEMA_signal_4139,
         new_AGEMA_signal_4143, new_AGEMA_signal_4147, new_AGEMA_signal_4151,
         new_AGEMA_signal_4155, new_AGEMA_signal_4159, new_AGEMA_signal_4163,
         new_AGEMA_signal_4167, new_AGEMA_signal_4171, new_AGEMA_signal_4175,
         new_AGEMA_signal_4179, new_AGEMA_signal_4183, new_AGEMA_signal_4187,
         new_AGEMA_signal_4191, new_AGEMA_signal_4195, new_AGEMA_signal_4199,
         new_AGEMA_signal_4203, new_AGEMA_signal_4207, new_AGEMA_signal_4211,
         new_AGEMA_signal_4215, new_AGEMA_signal_4219, new_AGEMA_signal_4223,
         new_AGEMA_signal_4227, new_AGEMA_signal_4231, new_AGEMA_signal_4235,
         new_AGEMA_signal_4239, new_AGEMA_signal_4243, new_AGEMA_signal_4247,
         new_AGEMA_signal_4251, new_AGEMA_signal_4255, new_AGEMA_signal_4259,
         new_AGEMA_signal_4263, new_AGEMA_signal_4267, new_AGEMA_signal_4271,
         new_AGEMA_signal_4275, new_AGEMA_signal_4279, new_AGEMA_signal_4283,
         new_AGEMA_signal_4287, new_AGEMA_signal_4291, new_AGEMA_signal_4295,
         new_AGEMA_signal_4299, new_AGEMA_signal_4303, new_AGEMA_signal_4307,
         new_AGEMA_signal_4311, new_AGEMA_signal_4315, new_AGEMA_signal_4319,
         new_AGEMA_signal_4323, new_AGEMA_signal_4327, new_AGEMA_signal_4331,
         new_AGEMA_signal_4335, new_AGEMA_signal_4339, new_AGEMA_signal_4343,
         new_AGEMA_signal_4345, new_AGEMA_signal_4347, new_AGEMA_signal_4355,
         new_AGEMA_signal_4357, new_AGEMA_signal_4359, new_AGEMA_signal_4361,
         new_AGEMA_signal_4365, new_AGEMA_signal_4369, new_AGEMA_signal_4379,
         new_AGEMA_signal_4381, new_AGEMA_signal_4383, new_AGEMA_signal_4391,
         new_AGEMA_signal_4393, new_AGEMA_signal_4395, new_AGEMA_signal_4397,
         new_AGEMA_signal_4401, new_AGEMA_signal_4405, new_AGEMA_signal_4415,
         new_AGEMA_signal_4417, new_AGEMA_signal_4419, new_AGEMA_signal_4427,
         new_AGEMA_signal_4429, new_AGEMA_signal_4431, new_AGEMA_signal_4433,
         new_AGEMA_signal_4437, new_AGEMA_signal_4441, new_AGEMA_signal_4451,
         new_AGEMA_signal_4453, new_AGEMA_signal_4455, new_AGEMA_signal_4463,
         new_AGEMA_signal_4465, new_AGEMA_signal_4467, new_AGEMA_signal_4469,
         new_AGEMA_signal_4473, new_AGEMA_signal_4477, new_AGEMA_signal_4487,
         new_AGEMA_signal_4489, new_AGEMA_signal_4491, new_AGEMA_signal_4499,
         new_AGEMA_signal_4501, new_AGEMA_signal_4503, new_AGEMA_signal_4505,
         new_AGEMA_signal_4509, new_AGEMA_signal_4513, new_AGEMA_signal_4523,
         new_AGEMA_signal_4525, new_AGEMA_signal_4527, new_AGEMA_signal_4535,
         new_AGEMA_signal_4537, new_AGEMA_signal_4539, new_AGEMA_signal_4541,
         new_AGEMA_signal_4545, new_AGEMA_signal_4549, new_AGEMA_signal_4559,
         new_AGEMA_signal_4561, new_AGEMA_signal_4563, new_AGEMA_signal_4571,
         new_AGEMA_signal_4573, new_AGEMA_signal_4575, new_AGEMA_signal_4577,
         new_AGEMA_signal_4581, new_AGEMA_signal_4585, new_AGEMA_signal_4595,
         new_AGEMA_signal_4597, new_AGEMA_signal_4599, new_AGEMA_signal_4607,
         new_AGEMA_signal_4609, new_AGEMA_signal_4611, new_AGEMA_signal_4613,
         new_AGEMA_signal_4617, new_AGEMA_signal_4621, new_AGEMA_signal_4631,
         new_AGEMA_signal_4633, new_AGEMA_signal_4635, new_AGEMA_signal_4643,
         new_AGEMA_signal_4645, new_AGEMA_signal_4647, new_AGEMA_signal_4649,
         new_AGEMA_signal_4653, new_AGEMA_signal_4657, new_AGEMA_signal_4667,
         new_AGEMA_signal_4669, new_AGEMA_signal_4671, new_AGEMA_signal_4679,
         new_AGEMA_signal_4681, new_AGEMA_signal_4683, new_AGEMA_signal_4685,
         new_AGEMA_signal_4689, new_AGEMA_signal_4693, new_AGEMA_signal_4703,
         new_AGEMA_signal_4705, new_AGEMA_signal_4707, new_AGEMA_signal_4715,
         new_AGEMA_signal_4717, new_AGEMA_signal_4719, new_AGEMA_signal_4721,
         new_AGEMA_signal_4725, new_AGEMA_signal_4729, new_AGEMA_signal_4739,
         new_AGEMA_signal_4741, new_AGEMA_signal_4743, new_AGEMA_signal_4751,
         new_AGEMA_signal_4753, new_AGEMA_signal_4755, new_AGEMA_signal_4757,
         new_AGEMA_signal_4761, new_AGEMA_signal_4765, new_AGEMA_signal_4775,
         new_AGEMA_signal_4777, new_AGEMA_signal_4779, new_AGEMA_signal_4787,
         new_AGEMA_signal_4789, new_AGEMA_signal_4791, new_AGEMA_signal_4793,
         new_AGEMA_signal_4797, new_AGEMA_signal_4801, new_AGEMA_signal_4811,
         new_AGEMA_signal_4813, new_AGEMA_signal_4815, new_AGEMA_signal_4823,
         new_AGEMA_signal_4825, new_AGEMA_signal_4827, new_AGEMA_signal_4829,
         new_AGEMA_signal_4833, new_AGEMA_signal_4837, new_AGEMA_signal_4847,
         new_AGEMA_signal_4849, new_AGEMA_signal_4851, new_AGEMA_signal_4859,
         new_AGEMA_signal_4861, new_AGEMA_signal_4863, new_AGEMA_signal_4865,
         new_AGEMA_signal_4869, new_AGEMA_signal_4873, new_AGEMA_signal_4883,
         new_AGEMA_signal_4885, new_AGEMA_signal_4887, new_AGEMA_signal_4895,
         new_AGEMA_signal_4897, new_AGEMA_signal_4899, new_AGEMA_signal_4901,
         new_AGEMA_signal_4905, new_AGEMA_signal_4909, new_AGEMA_signal_4919,
         new_AGEMA_signal_4923, new_AGEMA_signal_4927, new_AGEMA_signal_4931,
         new_AGEMA_signal_4935, new_AGEMA_signal_4939, new_AGEMA_signal_4943,
         new_AGEMA_signal_4947, new_AGEMA_signal_4951, new_AGEMA_signal_4955,
         new_AGEMA_signal_4959, new_AGEMA_signal_4963, new_AGEMA_signal_4967,
         new_AGEMA_signal_4971, new_AGEMA_signal_4975, new_AGEMA_signal_4979,
         new_AGEMA_signal_4983, new_AGEMA_signal_4987, new_AGEMA_signal_4991,
         new_AGEMA_signal_4995, new_AGEMA_signal_4999, new_AGEMA_signal_5003,
         new_AGEMA_signal_5007, new_AGEMA_signal_5011, new_AGEMA_signal_5015,
         new_AGEMA_signal_5019, new_AGEMA_signal_5023, new_AGEMA_signal_5027,
         new_AGEMA_signal_5031, new_AGEMA_signal_5035, new_AGEMA_signal_5039,
         new_AGEMA_signal_5043, new_AGEMA_signal_5047, new_AGEMA_signal_5051,
         new_AGEMA_signal_5055, new_AGEMA_signal_5059, new_AGEMA_signal_5063,
         new_AGEMA_signal_5067, new_AGEMA_signal_5071, new_AGEMA_signal_5075,
         new_AGEMA_signal_5079, new_AGEMA_signal_5083, new_AGEMA_signal_5087,
         new_AGEMA_signal_5091, new_AGEMA_signal_5095, new_AGEMA_signal_5099,
         new_AGEMA_signal_5103, new_AGEMA_signal_5107, new_AGEMA_signal_5111,
         new_AGEMA_signal_5115, new_AGEMA_signal_5119, new_AGEMA_signal_5123,
         new_AGEMA_signal_5319, new_AGEMA_signal_5323, new_AGEMA_signal_5327,
         new_AGEMA_signal_5331, new_AGEMA_signal_5335, new_AGEMA_signal_5339,
         new_AGEMA_signal_5343, new_AGEMA_signal_5347, new_AGEMA_signal_5351,
         new_AGEMA_signal_5355, new_AGEMA_signal_5359, new_AGEMA_signal_5363,
         new_AGEMA_signal_5367, new_AGEMA_signal_5371, new_AGEMA_signal_5375,
         new_AGEMA_signal_5379, new_AGEMA_signal_5383, new_AGEMA_signal_5387,
         new_AGEMA_signal_5391, new_AGEMA_signal_5395, new_AGEMA_signal_5399,
         new_AGEMA_signal_5403, new_AGEMA_signal_5407, new_AGEMA_signal_5411,
         new_AGEMA_signal_5415, new_AGEMA_signal_5419, new_AGEMA_signal_5423,
         new_AGEMA_signal_5427, new_AGEMA_signal_5431, new_AGEMA_signal_5435,
         new_AGEMA_signal_5439, new_AGEMA_signal_5443, new_AGEMA_signal_5447,
         new_AGEMA_signal_5451, new_AGEMA_signal_5455, new_AGEMA_signal_5459,
         new_AGEMA_signal_5463, new_AGEMA_signal_5467, new_AGEMA_signal_5471,
         new_AGEMA_signal_5475, new_AGEMA_signal_5479, new_AGEMA_signal_5483,
         new_AGEMA_signal_5487, new_AGEMA_signal_5491, new_AGEMA_signal_5495,
         new_AGEMA_signal_5499, new_AGEMA_signal_5503, new_AGEMA_signal_5507,
         new_AGEMA_signal_5511, new_AGEMA_signal_5515, new_AGEMA_signal_5519,
         new_AGEMA_signal_5523, new_AGEMA_signal_5527, new_AGEMA_signal_5531,
         new_AGEMA_signal_5535, new_AGEMA_signal_5539, new_AGEMA_signal_5543,
         new_AGEMA_signal_5547, new_AGEMA_signal_5551, new_AGEMA_signal_5555,
         new_AGEMA_signal_5559, new_AGEMA_signal_5563, new_AGEMA_signal_5567,
         new_AGEMA_signal_5571, new_AGEMA_signal_5575, new_AGEMA_signal_5579,
         new_AGEMA_signal_5583, new_AGEMA_signal_5587, new_AGEMA_signal_5591,
         new_AGEMA_signal_5595, new_AGEMA_signal_5599, new_AGEMA_signal_5603,
         new_AGEMA_signal_5607, new_AGEMA_signal_5611, new_AGEMA_signal_5615,
         new_AGEMA_signal_5619, new_AGEMA_signal_5623, new_AGEMA_signal_5627,
         new_AGEMA_signal_5631, new_AGEMA_signal_5635, new_AGEMA_signal_5639,
         new_AGEMA_signal_5643, new_AGEMA_signal_5647, new_AGEMA_signal_5651,
         new_AGEMA_signal_5655, new_AGEMA_signal_5659, new_AGEMA_signal_5663,
         new_AGEMA_signal_5667, new_AGEMA_signal_5671, new_AGEMA_signal_5675,
         new_AGEMA_signal_5679, new_AGEMA_signal_5683, new_AGEMA_signal_5687,
         new_AGEMA_signal_5691, new_AGEMA_signal_5695, new_AGEMA_signal_5699,
         new_AGEMA_signal_5703, new_AGEMA_signal_5707, new_AGEMA_signal_5711,
         new_AGEMA_signal_5715, new_AGEMA_signal_5719, new_AGEMA_signal_5723,
         new_AGEMA_signal_5727, new_AGEMA_signal_5731, new_AGEMA_signal_5735,
         new_AGEMA_signal_5739, new_AGEMA_signal_5743, new_AGEMA_signal_5747,
         new_AGEMA_signal_5751, new_AGEMA_signal_5755, new_AGEMA_signal_5759,
         new_AGEMA_signal_5763, new_AGEMA_signal_5767, new_AGEMA_signal_5771,
         new_AGEMA_signal_5775, new_AGEMA_signal_5779, new_AGEMA_signal_5783,
         new_AGEMA_signal_5787, new_AGEMA_signal_5791, new_AGEMA_signal_5795,
         new_AGEMA_signal_5799, new_AGEMA_signal_5803, new_AGEMA_signal_5807,
         new_AGEMA_signal_5811, new_AGEMA_signal_5815, new_AGEMA_signal_5819,
         new_AGEMA_signal_5823, new_AGEMA_signal_5827, new_AGEMA_signal_5831,
         new_AGEMA_signal_5835, new_AGEMA_signal_5839, new_AGEMA_signal_5843,
         new_AGEMA_signal_5847, new_AGEMA_signal_5851, new_AGEMA_signal_5855,
         new_AGEMA_signal_5859, new_AGEMA_signal_5863, new_AGEMA_signal_5867,
         new_AGEMA_signal_5871, new_AGEMA_signal_5875, new_AGEMA_signal_5879,
         new_AGEMA_signal_5883, new_AGEMA_signal_5887, new_AGEMA_signal_5891,
         new_AGEMA_signal_5895, new_AGEMA_signal_5899, new_AGEMA_signal_5903,
         new_AGEMA_signal_5907, new_AGEMA_signal_5911, new_AGEMA_signal_5915,
         new_AGEMA_signal_5919, new_AGEMA_signal_5923, new_AGEMA_signal_5927,
         new_AGEMA_signal_5931, new_AGEMA_signal_5935, new_AGEMA_signal_5939,
         new_AGEMA_signal_5943, new_AGEMA_signal_5947, new_AGEMA_signal_5951,
         new_AGEMA_signal_5955, new_AGEMA_signal_5959, new_AGEMA_signal_5963,
         new_AGEMA_signal_5967, new_AGEMA_signal_5971, new_AGEMA_signal_5975,
         new_AGEMA_signal_5979, new_AGEMA_signal_5983, new_AGEMA_signal_5987,
         new_AGEMA_signal_5991, new_AGEMA_signal_5995, new_AGEMA_signal_5999,
         new_AGEMA_signal_6003, new_AGEMA_signal_6007, new_AGEMA_signal_6011,
         new_AGEMA_signal_6015, new_AGEMA_signal_6019, new_AGEMA_signal_6023,
         new_AGEMA_signal_6027, new_AGEMA_signal_6031, new_AGEMA_signal_6035,
         new_AGEMA_signal_6039, new_AGEMA_signal_6043, new_AGEMA_signal_6047,
         new_AGEMA_signal_6051, new_AGEMA_signal_6055, new_AGEMA_signal_6059,
         new_AGEMA_signal_6063, new_AGEMA_signal_6067, new_AGEMA_signal_6071,
         new_AGEMA_signal_6075, new_AGEMA_signal_6079, new_AGEMA_signal_6083,
         new_AGEMA_signal_6087, new_AGEMA_signal_6091, new_AGEMA_signal_6095,
         new_AGEMA_signal_6099, new_AGEMA_signal_6103, new_AGEMA_signal_6107,
         new_AGEMA_signal_3956, new_AGEMA_signal_3960, new_AGEMA_signal_3964,
         new_AGEMA_signal_3968, new_AGEMA_signal_3972, new_AGEMA_signal_3976,
         new_AGEMA_signal_3980, new_AGEMA_signal_3984, new_AGEMA_signal_3988,
         new_AGEMA_signal_3992, new_AGEMA_signal_3996, new_AGEMA_signal_4000,
         new_AGEMA_signal_4004, new_AGEMA_signal_4008, new_AGEMA_signal_4012,
         new_AGEMA_signal_4016, new_AGEMA_signal_4020, new_AGEMA_signal_4024,
         new_AGEMA_signal_4028, new_AGEMA_signal_4032, new_AGEMA_signal_4036,
         new_AGEMA_signal_4040, new_AGEMA_signal_4044, new_AGEMA_signal_4048,
         new_AGEMA_signal_4052, new_AGEMA_signal_4056, new_AGEMA_signal_4060,
         new_AGEMA_signal_4064, new_AGEMA_signal_4068, new_AGEMA_signal_4072,
         new_AGEMA_signal_4076, new_AGEMA_signal_4080, new_AGEMA_signal_4084,
         new_AGEMA_signal_4088, new_AGEMA_signal_4092, new_AGEMA_signal_4096,
         new_AGEMA_signal_4100, new_AGEMA_signal_4104, new_AGEMA_signal_4108,
         new_AGEMA_signal_4112, new_AGEMA_signal_4116, new_AGEMA_signal_4120,
         new_AGEMA_signal_4124, new_AGEMA_signal_4128, new_AGEMA_signal_4132,
         new_AGEMA_signal_4136, new_AGEMA_signal_4140, new_AGEMA_signal_4144,
         new_AGEMA_signal_4148, new_AGEMA_signal_4152, new_AGEMA_signal_4156,
         new_AGEMA_signal_4160, new_AGEMA_signal_4164, new_AGEMA_signal_4168,
         new_AGEMA_signal_4172, new_AGEMA_signal_4176, new_AGEMA_signal_4180,
         new_AGEMA_signal_4184, new_AGEMA_signal_4188, new_AGEMA_signal_4192,
         new_AGEMA_signal_4196, new_AGEMA_signal_4200, new_AGEMA_signal_4204,
         new_AGEMA_signal_4208, new_AGEMA_signal_4212, new_AGEMA_signal_4216,
         new_AGEMA_signal_4220, new_AGEMA_signal_4224, new_AGEMA_signal_4228,
         new_AGEMA_signal_4232, new_AGEMA_signal_4236, new_AGEMA_signal_4240,
         new_AGEMA_signal_4244, new_AGEMA_signal_4248, new_AGEMA_signal_4252,
         new_AGEMA_signal_4256, new_AGEMA_signal_4260, new_AGEMA_signal_4264,
         new_AGEMA_signal_4268, new_AGEMA_signal_4272, new_AGEMA_signal_4276,
         new_AGEMA_signal_4280, new_AGEMA_signal_4284, new_AGEMA_signal_4288,
         new_AGEMA_signal_4292, new_AGEMA_signal_4296, new_AGEMA_signal_4300,
         new_AGEMA_signal_4304, new_AGEMA_signal_4308, new_AGEMA_signal_4312,
         new_AGEMA_signal_4316, new_AGEMA_signal_4320, new_AGEMA_signal_4324,
         new_AGEMA_signal_4328, new_AGEMA_signal_4332, new_AGEMA_signal_4336,
         new_AGEMA_signal_4340, new_AGEMA_signal_4348, new_AGEMA_signal_4350,
         new_AGEMA_signal_4352, new_AGEMA_signal_4362, new_AGEMA_signal_4366,
         new_AGEMA_signal_4370, new_AGEMA_signal_4372, new_AGEMA_signal_4374,
         new_AGEMA_signal_4376, new_AGEMA_signal_4384, new_AGEMA_signal_4386,
         new_AGEMA_signal_4388, new_AGEMA_signal_4398, new_AGEMA_signal_4402,
         new_AGEMA_signal_4406, new_AGEMA_signal_4408, new_AGEMA_signal_4410,
         new_AGEMA_signal_4412, new_AGEMA_signal_4420, new_AGEMA_signal_4422,
         new_AGEMA_signal_4424, new_AGEMA_signal_4434, new_AGEMA_signal_4438,
         new_AGEMA_signal_4442, new_AGEMA_signal_4444, new_AGEMA_signal_4446,
         new_AGEMA_signal_4448, new_AGEMA_signal_4456, new_AGEMA_signal_4458,
         new_AGEMA_signal_4460, new_AGEMA_signal_4470, new_AGEMA_signal_4474,
         new_AGEMA_signal_4478, new_AGEMA_signal_4480, new_AGEMA_signal_4482,
         new_AGEMA_signal_4484, new_AGEMA_signal_4492, new_AGEMA_signal_4494,
         new_AGEMA_signal_4496, new_AGEMA_signal_4506, new_AGEMA_signal_4510,
         new_AGEMA_signal_4514, new_AGEMA_signal_4516, new_AGEMA_signal_4518,
         new_AGEMA_signal_4520, new_AGEMA_signal_4528, new_AGEMA_signal_4530,
         new_AGEMA_signal_4532, new_AGEMA_signal_4542, new_AGEMA_signal_4546,
         new_AGEMA_signal_4550, new_AGEMA_signal_4552, new_AGEMA_signal_4554,
         new_AGEMA_signal_4556, new_AGEMA_signal_4564, new_AGEMA_signal_4566,
         new_AGEMA_signal_4568, new_AGEMA_signal_4578, new_AGEMA_signal_4582,
         new_AGEMA_signal_4586, new_AGEMA_signal_4588, new_AGEMA_signal_4590,
         new_AGEMA_signal_4592, new_AGEMA_signal_4600, new_AGEMA_signal_4602,
         new_AGEMA_signal_4604, new_AGEMA_signal_4614, new_AGEMA_signal_4618,
         new_AGEMA_signal_4622, new_AGEMA_signal_4624, new_AGEMA_signal_4626,
         new_AGEMA_signal_4628, new_AGEMA_signal_4636, new_AGEMA_signal_4638,
         new_AGEMA_signal_4640, new_AGEMA_signal_4650, new_AGEMA_signal_4654,
         new_AGEMA_signal_4658, new_AGEMA_signal_4660, new_AGEMA_signal_4662,
         new_AGEMA_signal_4664, new_AGEMA_signal_4672, new_AGEMA_signal_4674,
         new_AGEMA_signal_4676, new_AGEMA_signal_4686, new_AGEMA_signal_4690,
         new_AGEMA_signal_4694, new_AGEMA_signal_4696, new_AGEMA_signal_4698,
         new_AGEMA_signal_4700, new_AGEMA_signal_4708, new_AGEMA_signal_4710,
         new_AGEMA_signal_4712, new_AGEMA_signal_4722, new_AGEMA_signal_4726,
         new_AGEMA_signal_4730, new_AGEMA_signal_4732, new_AGEMA_signal_4734,
         new_AGEMA_signal_4736, new_AGEMA_signal_4744, new_AGEMA_signal_4746,
         new_AGEMA_signal_4748, new_AGEMA_signal_4758, new_AGEMA_signal_4762,
         new_AGEMA_signal_4766, new_AGEMA_signal_4768, new_AGEMA_signal_4770,
         new_AGEMA_signal_4772, new_AGEMA_signal_4780, new_AGEMA_signal_4782,
         new_AGEMA_signal_4784, new_AGEMA_signal_4794, new_AGEMA_signal_4798,
         new_AGEMA_signal_4802, new_AGEMA_signal_4804, new_AGEMA_signal_4806,
         new_AGEMA_signal_4808, new_AGEMA_signal_4816, new_AGEMA_signal_4818,
         new_AGEMA_signal_4820, new_AGEMA_signal_4830, new_AGEMA_signal_4834,
         new_AGEMA_signal_4838, new_AGEMA_signal_4840, new_AGEMA_signal_4842,
         new_AGEMA_signal_4844, new_AGEMA_signal_4852, new_AGEMA_signal_4854,
         new_AGEMA_signal_4856, new_AGEMA_signal_4866, new_AGEMA_signal_4870,
         new_AGEMA_signal_4874, new_AGEMA_signal_4876, new_AGEMA_signal_4878,
         new_AGEMA_signal_4880, new_AGEMA_signal_4888, new_AGEMA_signal_4890,
         new_AGEMA_signal_4892, new_AGEMA_signal_4902, new_AGEMA_signal_4906,
         new_AGEMA_signal_4910, new_AGEMA_signal_4912, new_AGEMA_signal_4914,
         new_AGEMA_signal_4916, new_AGEMA_signal_4920, new_AGEMA_signal_4924,
         new_AGEMA_signal_4928, new_AGEMA_signal_4932, new_AGEMA_signal_4936,
         new_AGEMA_signal_4940, new_AGEMA_signal_4944, new_AGEMA_signal_4948,
         new_AGEMA_signal_4952, new_AGEMA_signal_4956, new_AGEMA_signal_4960,
         new_AGEMA_signal_4964, new_AGEMA_signal_4968, new_AGEMA_signal_4972,
         new_AGEMA_signal_4976, new_AGEMA_signal_4980, new_AGEMA_signal_4984,
         new_AGEMA_signal_4988, new_AGEMA_signal_4992, new_AGEMA_signal_4996,
         new_AGEMA_signal_5000, new_AGEMA_signal_5004, new_AGEMA_signal_5008,
         new_AGEMA_signal_5012, new_AGEMA_signal_5016, new_AGEMA_signal_5020,
         new_AGEMA_signal_5024, new_AGEMA_signal_5028, new_AGEMA_signal_5032,
         new_AGEMA_signal_5036, new_AGEMA_signal_5040, new_AGEMA_signal_5044,
         new_AGEMA_signal_5048, new_AGEMA_signal_5052, new_AGEMA_signal_5056,
         new_AGEMA_signal_5060, new_AGEMA_signal_5064, new_AGEMA_signal_5068,
         new_AGEMA_signal_5072, new_AGEMA_signal_5076, new_AGEMA_signal_5080,
         new_AGEMA_signal_5084, new_AGEMA_signal_5088, new_AGEMA_signal_5092,
         new_AGEMA_signal_5096, new_AGEMA_signal_5100, new_AGEMA_signal_5104,
         new_AGEMA_signal_5108, new_AGEMA_signal_5112, new_AGEMA_signal_5116,
         new_AGEMA_signal_5120, new_AGEMA_signal_5124, new_AGEMA_signal_5126,
         new_AGEMA_signal_5128, new_AGEMA_signal_5130, new_AGEMA_signal_5132,
         new_AGEMA_signal_5134, new_AGEMA_signal_5136, new_AGEMA_signal_5138,
         new_AGEMA_signal_5140, new_AGEMA_signal_5142, new_AGEMA_signal_5144,
         new_AGEMA_signal_5146, new_AGEMA_signal_5148, new_AGEMA_signal_5150,
         new_AGEMA_signal_5152, new_AGEMA_signal_5154, new_AGEMA_signal_5156,
         new_AGEMA_signal_5158, new_AGEMA_signal_5160, new_AGEMA_signal_5162,
         new_AGEMA_signal_5164, new_AGEMA_signal_5166, new_AGEMA_signal_5168,
         new_AGEMA_signal_5170, new_AGEMA_signal_5172, new_AGEMA_signal_5174,
         new_AGEMA_signal_5176, new_AGEMA_signal_5178, new_AGEMA_signal_5180,
         new_AGEMA_signal_5182, new_AGEMA_signal_5184, new_AGEMA_signal_5186,
         new_AGEMA_signal_5188, new_AGEMA_signal_5190, new_AGEMA_signal_5192,
         new_AGEMA_signal_5194, new_AGEMA_signal_5196, new_AGEMA_signal_5198,
         new_AGEMA_signal_5200, new_AGEMA_signal_5202, new_AGEMA_signal_5204,
         new_AGEMA_signal_5206, new_AGEMA_signal_5208, new_AGEMA_signal_5210,
         new_AGEMA_signal_5212, new_AGEMA_signal_5214, new_AGEMA_signal_5216,
         new_AGEMA_signal_5218, new_AGEMA_signal_5220, new_AGEMA_signal_5222,
         new_AGEMA_signal_5224, new_AGEMA_signal_5226, new_AGEMA_signal_5228,
         new_AGEMA_signal_5230, new_AGEMA_signal_5232, new_AGEMA_signal_5234,
         new_AGEMA_signal_5236, new_AGEMA_signal_5238, new_AGEMA_signal_5240,
         new_AGEMA_signal_5242, new_AGEMA_signal_5244, new_AGEMA_signal_5246,
         new_AGEMA_signal_5248, new_AGEMA_signal_5250, new_AGEMA_signal_5252,
         new_AGEMA_signal_5254, new_AGEMA_signal_5256, new_AGEMA_signal_5258,
         new_AGEMA_signal_5260, new_AGEMA_signal_5262, new_AGEMA_signal_5264,
         new_AGEMA_signal_5266, new_AGEMA_signal_5268, new_AGEMA_signal_5270,
         new_AGEMA_signal_5272, new_AGEMA_signal_5274, new_AGEMA_signal_5276,
         new_AGEMA_signal_5278, new_AGEMA_signal_5280, new_AGEMA_signal_5282,
         new_AGEMA_signal_5284, new_AGEMA_signal_5286, new_AGEMA_signal_5288,
         new_AGEMA_signal_5290, new_AGEMA_signal_5292, new_AGEMA_signal_5294,
         new_AGEMA_signal_5296, new_AGEMA_signal_5298, new_AGEMA_signal_5300,
         new_AGEMA_signal_5302, new_AGEMA_signal_5304, new_AGEMA_signal_5306,
         new_AGEMA_signal_5308, new_AGEMA_signal_5310, new_AGEMA_signal_5312,
         new_AGEMA_signal_5314, new_AGEMA_signal_5316, new_AGEMA_signal_5320,
         new_AGEMA_signal_5324, new_AGEMA_signal_5328, new_AGEMA_signal_5332,
         new_AGEMA_signal_5336, new_AGEMA_signal_5340, new_AGEMA_signal_5344,
         new_AGEMA_signal_5348, new_AGEMA_signal_5352, new_AGEMA_signal_5356,
         new_AGEMA_signal_5360, new_AGEMA_signal_5364, new_AGEMA_signal_5368,
         new_AGEMA_signal_5372, new_AGEMA_signal_5376, new_AGEMA_signal_5380,
         new_AGEMA_signal_5384, new_AGEMA_signal_5388, new_AGEMA_signal_5392,
         new_AGEMA_signal_5396, new_AGEMA_signal_5400, new_AGEMA_signal_5404,
         new_AGEMA_signal_5408, new_AGEMA_signal_5412, new_AGEMA_signal_5416,
         new_AGEMA_signal_5420, new_AGEMA_signal_5424, new_AGEMA_signal_5428,
         new_AGEMA_signal_5432, new_AGEMA_signal_5436, new_AGEMA_signal_5440,
         new_AGEMA_signal_5444, new_AGEMA_signal_5448, new_AGEMA_signal_5452,
         new_AGEMA_signal_5456, new_AGEMA_signal_5460, new_AGEMA_signal_5464,
         new_AGEMA_signal_5468, new_AGEMA_signal_5472, new_AGEMA_signal_5476,
         new_AGEMA_signal_5480, new_AGEMA_signal_5484, new_AGEMA_signal_5488,
         new_AGEMA_signal_5492, new_AGEMA_signal_5496, new_AGEMA_signal_5500,
         new_AGEMA_signal_5504, new_AGEMA_signal_5508, new_AGEMA_signal_5512,
         new_AGEMA_signal_5516, new_AGEMA_signal_5520, new_AGEMA_signal_5524,
         new_AGEMA_signal_5528, new_AGEMA_signal_5532, new_AGEMA_signal_5536,
         new_AGEMA_signal_5540, new_AGEMA_signal_5544, new_AGEMA_signal_5548,
         new_AGEMA_signal_5552, new_AGEMA_signal_5556, new_AGEMA_signal_5560,
         new_AGEMA_signal_5564, new_AGEMA_signal_5568, new_AGEMA_signal_5572,
         new_AGEMA_signal_5576, new_AGEMA_signal_5580, new_AGEMA_signal_5584,
         new_AGEMA_signal_5588, new_AGEMA_signal_5592, new_AGEMA_signal_5596,
         new_AGEMA_signal_5600, new_AGEMA_signal_5604, new_AGEMA_signal_5608,
         new_AGEMA_signal_5612, new_AGEMA_signal_5616, new_AGEMA_signal_5620,
         new_AGEMA_signal_5624, new_AGEMA_signal_5628, new_AGEMA_signal_5632,
         new_AGEMA_signal_5636, new_AGEMA_signal_5640, new_AGEMA_signal_5644,
         new_AGEMA_signal_5648, new_AGEMA_signal_5652, new_AGEMA_signal_5656,
         new_AGEMA_signal_5660, new_AGEMA_signal_5664, new_AGEMA_signal_5668,
         new_AGEMA_signal_5672, new_AGEMA_signal_5676, new_AGEMA_signal_5680,
         new_AGEMA_signal_5684, new_AGEMA_signal_5688, new_AGEMA_signal_5692,
         new_AGEMA_signal_5696, new_AGEMA_signal_5700, new_AGEMA_signal_5704,
         new_AGEMA_signal_5708, new_AGEMA_signal_5712, new_AGEMA_signal_5716,
         new_AGEMA_signal_5720, new_AGEMA_signal_5724, new_AGEMA_signal_5728,
         new_AGEMA_signal_5732, new_AGEMA_signal_5736, new_AGEMA_signal_5740,
         new_AGEMA_signal_5744, new_AGEMA_signal_5748, new_AGEMA_signal_5752,
         new_AGEMA_signal_5756, new_AGEMA_signal_5760, new_AGEMA_signal_5764,
         new_AGEMA_signal_5768, new_AGEMA_signal_5772, new_AGEMA_signal_5776,
         new_AGEMA_signal_5780, new_AGEMA_signal_5784, new_AGEMA_signal_5788,
         new_AGEMA_signal_5792, new_AGEMA_signal_5796, new_AGEMA_signal_5800,
         new_AGEMA_signal_5804, new_AGEMA_signal_5808, new_AGEMA_signal_5812,
         new_AGEMA_signal_5816, new_AGEMA_signal_5820, new_AGEMA_signal_5824,
         new_AGEMA_signal_5828, new_AGEMA_signal_5832, new_AGEMA_signal_5836,
         new_AGEMA_signal_5840, new_AGEMA_signal_5844, new_AGEMA_signal_5848,
         new_AGEMA_signal_5852, new_AGEMA_signal_5856, new_AGEMA_signal_5860,
         new_AGEMA_signal_5864, new_AGEMA_signal_5868, new_AGEMA_signal_5872,
         new_AGEMA_signal_5876, new_AGEMA_signal_5880, new_AGEMA_signal_5884,
         new_AGEMA_signal_5888, new_AGEMA_signal_5892, new_AGEMA_signal_5896,
         new_AGEMA_signal_5900, new_AGEMA_signal_5904, new_AGEMA_signal_5908,
         new_AGEMA_signal_5912, new_AGEMA_signal_5916, new_AGEMA_signal_5920,
         new_AGEMA_signal_5924, new_AGEMA_signal_5928, new_AGEMA_signal_5932,
         new_AGEMA_signal_5936, new_AGEMA_signal_5940, new_AGEMA_signal_5944,
         new_AGEMA_signal_5948, new_AGEMA_signal_5952, new_AGEMA_signal_5956,
         new_AGEMA_signal_5960, new_AGEMA_signal_5964, new_AGEMA_signal_5968,
         new_AGEMA_signal_5972, new_AGEMA_signal_5976, new_AGEMA_signal_5980,
         new_AGEMA_signal_5984, new_AGEMA_signal_5988, new_AGEMA_signal_5992,
         new_AGEMA_signal_5996, new_AGEMA_signal_6000, new_AGEMA_signal_6004,
         new_AGEMA_signal_6008, new_AGEMA_signal_6012, new_AGEMA_signal_6016,
         new_AGEMA_signal_6020, new_AGEMA_signal_6024, new_AGEMA_signal_6028,
         new_AGEMA_signal_6032, new_AGEMA_signal_6036, new_AGEMA_signal_6040,
         new_AGEMA_signal_6044, new_AGEMA_signal_6048, new_AGEMA_signal_6052,
         new_AGEMA_signal_6056, new_AGEMA_signal_6060, new_AGEMA_signal_6064,
         new_AGEMA_signal_6068, new_AGEMA_signal_6072, new_AGEMA_signal_6076,
         new_AGEMA_signal_6080, new_AGEMA_signal_6084, new_AGEMA_signal_6088,
         new_AGEMA_signal_6092, new_AGEMA_signal_6096, new_AGEMA_signal_6100,
         new_AGEMA_signal_6104, new_AGEMA_signal_6108, new_AGEMA_signal_3957,
         new_AGEMA_signal_2909, new_AGEMA_signal_2908, new_AGEMA_signal_3969,
         new_AGEMA_signal_3965, new_AGEMA_signal_3961, new_AGEMA_signal_2891,
         new_AGEMA_signal_2890, new_AGEMA_signal_2995, new_AGEMA_signal_2994,
         new_AGEMA_signal_3981, new_AGEMA_signal_3977, new_AGEMA_signal_3973,
         new_AGEMA_signal_2983, new_AGEMA_signal_2982, new_AGEMA_signal_2913,
         new_AGEMA_signal_2912, new_AGEMA_signal_3993, new_AGEMA_signal_3989,
         new_AGEMA_signal_3985, new_AGEMA_signal_2895, new_AGEMA_signal_2894,
         new_AGEMA_signal_2999, new_AGEMA_signal_2998, new_AGEMA_signal_4005,
         new_AGEMA_signal_4001, new_AGEMA_signal_3997, new_AGEMA_signal_2985,
         new_AGEMA_signal_2984, new_AGEMA_signal_2917, new_AGEMA_signal_2916,
         new_AGEMA_signal_4017, new_AGEMA_signal_4013, new_AGEMA_signal_4009,
         new_AGEMA_signal_2899, new_AGEMA_signal_2898, new_AGEMA_signal_3003,
         new_AGEMA_signal_3002, new_AGEMA_signal_4029, new_AGEMA_signal_4025,
         new_AGEMA_signal_4021, new_AGEMA_signal_2987, new_AGEMA_signal_2986,
         new_AGEMA_signal_3059, new_AGEMA_signal_3058, new_AGEMA_signal_4041,
         new_AGEMA_signal_4037, new_AGEMA_signal_4033, new_AGEMA_signal_3053,
         new_AGEMA_signal_3052, new_AGEMA_signal_3077, new_AGEMA_signal_3076,
         new_AGEMA_signal_4053, new_AGEMA_signal_4049, new_AGEMA_signal_4045,
         new_AGEMA_signal_3073, new_AGEMA_signal_3072, new_AGEMA_signal_2925,
         new_AGEMA_signal_2924, new_AGEMA_signal_4065, new_AGEMA_signal_4061,
         new_AGEMA_signal_4057, new_AGEMA_signal_2875, new_AGEMA_signal_2874,
         new_AGEMA_signal_3011, new_AGEMA_signal_3010, new_AGEMA_signal_4077,
         new_AGEMA_signal_4073, new_AGEMA_signal_4069, new_AGEMA_signal_2973,
         new_AGEMA_signal_2972, new_AGEMA_signal_2929, new_AGEMA_signal_2928,
         new_AGEMA_signal_4089, new_AGEMA_signal_4085, new_AGEMA_signal_4081,
         new_AGEMA_signal_2879, new_AGEMA_signal_2878, new_AGEMA_signal_3015,
         new_AGEMA_signal_3014, new_AGEMA_signal_4101, new_AGEMA_signal_4097,
         new_AGEMA_signal_4093, new_AGEMA_signal_2975, new_AGEMA_signal_2974,
         new_AGEMA_signal_3063, new_AGEMA_signal_3062, new_AGEMA_signal_4113,
         new_AGEMA_signal_4109, new_AGEMA_signal_4105, new_AGEMA_signal_3049,
         new_AGEMA_signal_3048, new_AGEMA_signal_3081, new_AGEMA_signal_3080,
         new_AGEMA_signal_4125, new_AGEMA_signal_4121, new_AGEMA_signal_4117,
         new_AGEMA_signal_3071, new_AGEMA_signal_3070, new_AGEMA_signal_2937,
         new_AGEMA_signal_2936, new_AGEMA_signal_4137, new_AGEMA_signal_4133,
         new_AGEMA_signal_4129, new_AGEMA_signal_2887, new_AGEMA_signal_2886,
         new_AGEMA_signal_3023, new_AGEMA_signal_3022, new_AGEMA_signal_4149,
         new_AGEMA_signal_4145, new_AGEMA_signal_4141, new_AGEMA_signal_2981,
         new_AGEMA_signal_2980, new_AGEMA_signal_2705, new_AGEMA_signal_2704,
         new_AGEMA_signal_4161, new_AGEMA_signal_4157, new_AGEMA_signal_4153,
         new_AGEMA_signal_2621, new_AGEMA_signal_2620, new_AGEMA_signal_2825,
         new_AGEMA_signal_2824, new_AGEMA_signal_4173, new_AGEMA_signal_4169,
         new_AGEMA_signal_4165, new_AGEMA_signal_2745, new_AGEMA_signal_2744,
         new_AGEMA_signal_2709, new_AGEMA_signal_2708, new_AGEMA_signal_4185,
         new_AGEMA_signal_4181, new_AGEMA_signal_4177, new_AGEMA_signal_2625,
         new_AGEMA_signal_2624, new_AGEMA_signal_2829, new_AGEMA_signal_2828,
         new_AGEMA_signal_4197, new_AGEMA_signal_4193, new_AGEMA_signal_4189,
         new_AGEMA_signal_2747, new_AGEMA_signal_2746, new_AGEMA_signal_2713,
         new_AGEMA_signal_2712, new_AGEMA_signal_4209, new_AGEMA_signal_4205,
         new_AGEMA_signal_4201, new_AGEMA_signal_2629, new_AGEMA_signal_2628,
         new_AGEMA_signal_2833, new_AGEMA_signal_2832, new_AGEMA_signal_4221,
         new_AGEMA_signal_4217, new_AGEMA_signal_4213, new_AGEMA_signal_2749,
         new_AGEMA_signal_2748, new_AGEMA_signal_2941, new_AGEMA_signal_2940,
         new_AGEMA_signal_4233, new_AGEMA_signal_4229, new_AGEMA_signal_4225,
         new_AGEMA_signal_2855, new_AGEMA_signal_2854, new_AGEMA_signal_3027,
         new_AGEMA_signal_3026, new_AGEMA_signal_4245, new_AGEMA_signal_4241,
         new_AGEMA_signal_4237, new_AGEMA_signal_2961, new_AGEMA_signal_2960,
         new_AGEMA_signal_2945, new_AGEMA_signal_2944, new_AGEMA_signal_4257,
         new_AGEMA_signal_4253, new_AGEMA_signal_4249, new_AGEMA_signal_2859,
         new_AGEMA_signal_2858, new_AGEMA_signal_3031, new_AGEMA_signal_3030,
         new_AGEMA_signal_4269, new_AGEMA_signal_4265, new_AGEMA_signal_4261,
         new_AGEMA_signal_2963, new_AGEMA_signal_2962, new_AGEMA_signal_2949,
         new_AGEMA_signal_2948, new_AGEMA_signal_4281, new_AGEMA_signal_4277,
         new_AGEMA_signal_4273, new_AGEMA_signal_2863, new_AGEMA_signal_2862,
         new_AGEMA_signal_3035, new_AGEMA_signal_3034, new_AGEMA_signal_4293,
         new_AGEMA_signal_4289, new_AGEMA_signal_4285, new_AGEMA_signal_2965,
         new_AGEMA_signal_2964, new_AGEMA_signal_2953, new_AGEMA_signal_2952,
         new_AGEMA_signal_4305, new_AGEMA_signal_4301, new_AGEMA_signal_4297,
         new_AGEMA_signal_2867, new_AGEMA_signal_2866, new_AGEMA_signal_3039,
         new_AGEMA_signal_3038, new_AGEMA_signal_4317, new_AGEMA_signal_4313,
         new_AGEMA_signal_4309, new_AGEMA_signal_2967, new_AGEMA_signal_2966,
         new_AGEMA_signal_3067, new_AGEMA_signal_3066, new_AGEMA_signal_4329,
         new_AGEMA_signal_4325, new_AGEMA_signal_4321, new_AGEMA_signal_3045,
         new_AGEMA_signal_3044, new_AGEMA_signal_3085, new_AGEMA_signal_3084,
         new_AGEMA_signal_4341, new_AGEMA_signal_4337, new_AGEMA_signal_4333,
         new_AGEMA_signal_3069, new_AGEMA_signal_3068, new_AGEMA_signal_2159,
         new_AGEMA_signal_2158, SubCellInst_SboxInst_0_T1,
         new_AGEMA_signal_2287, new_AGEMA_signal_2286,
         SubCellInst_SboxInst_0_L0, new_AGEMA_signal_4353,
         new_AGEMA_signal_4351, new_AGEMA_signal_4349, new_AGEMA_signal_2161,
         new_AGEMA_signal_2160, SubCellInst_SboxInst_0_T3,
         new_AGEMA_signal_2373, new_AGEMA_signal_2372,
         SubCellInst_SboxInst_0_YY_3, new_AGEMA_signal_4371,
         new_AGEMA_signal_4367, new_AGEMA_signal_4363, new_AGEMA_signal_2375,
         new_AGEMA_signal_2374, new_AGEMA_signal_2489, new_AGEMA_signal_2488,
         new_AGEMA_signal_4377, new_AGEMA_signal_4375, new_AGEMA_signal_4373,
         new_AGEMA_signal_2167, new_AGEMA_signal_2166,
         SubCellInst_SboxInst_1_T1, new_AGEMA_signal_2291,
         new_AGEMA_signal_2290, SubCellInst_SboxInst_1_L0,
         new_AGEMA_signal_4389, new_AGEMA_signal_4387, new_AGEMA_signal_4385,
         new_AGEMA_signal_2169, new_AGEMA_signal_2168,
         SubCellInst_SboxInst_1_T3, new_AGEMA_signal_2377,
         new_AGEMA_signal_2376, SubCellInst_SboxInst_1_YY_3,
         new_AGEMA_signal_4407, new_AGEMA_signal_4403, new_AGEMA_signal_4399,
         new_AGEMA_signal_2379, new_AGEMA_signal_2378, new_AGEMA_signal_2491,
         new_AGEMA_signal_2490, new_AGEMA_signal_4413, new_AGEMA_signal_4411,
         new_AGEMA_signal_4409, new_AGEMA_signal_2175, new_AGEMA_signal_2174,
         SubCellInst_SboxInst_2_T1, new_AGEMA_signal_2295,
         new_AGEMA_signal_2294, SubCellInst_SboxInst_2_L0,
         new_AGEMA_signal_4425, new_AGEMA_signal_4423, new_AGEMA_signal_4421,
         new_AGEMA_signal_2177, new_AGEMA_signal_2176,
         SubCellInst_SboxInst_2_T3, new_AGEMA_signal_2381,
         new_AGEMA_signal_2380, SubCellInst_SboxInst_2_YY_3,
         new_AGEMA_signal_4443, new_AGEMA_signal_4439, new_AGEMA_signal_4435,
         new_AGEMA_signal_2383, new_AGEMA_signal_2382, new_AGEMA_signal_2493,
         new_AGEMA_signal_2492, new_AGEMA_signal_4449, new_AGEMA_signal_4447,
         new_AGEMA_signal_4445, new_AGEMA_signal_2183, new_AGEMA_signal_2182,
         SubCellInst_SboxInst_3_T1, new_AGEMA_signal_2299,
         new_AGEMA_signal_2298, SubCellInst_SboxInst_3_L0,
         new_AGEMA_signal_4461, new_AGEMA_signal_4459, new_AGEMA_signal_4457,
         new_AGEMA_signal_2185, new_AGEMA_signal_2184,
         SubCellInst_SboxInst_3_T3, new_AGEMA_signal_2385,
         new_AGEMA_signal_2384, SubCellInst_SboxInst_3_YY_3,
         new_AGEMA_signal_4479, new_AGEMA_signal_4475, new_AGEMA_signal_4471,
         new_AGEMA_signal_2387, new_AGEMA_signal_2386, new_AGEMA_signal_2495,
         new_AGEMA_signal_2494, new_AGEMA_signal_4485, new_AGEMA_signal_4483,
         new_AGEMA_signal_4481, new_AGEMA_signal_2191, new_AGEMA_signal_2190,
         SubCellInst_SboxInst_4_T1, new_AGEMA_signal_2303,
         new_AGEMA_signal_2302, SubCellInst_SboxInst_4_L0,
         new_AGEMA_signal_4497, new_AGEMA_signal_4495, new_AGEMA_signal_4493,
         new_AGEMA_signal_2193, new_AGEMA_signal_2192,
         SubCellInst_SboxInst_4_T3, new_AGEMA_signal_2389,
         new_AGEMA_signal_2388, SubCellInst_SboxInst_4_YY_3,
         new_AGEMA_signal_4515, new_AGEMA_signal_4511, new_AGEMA_signal_4507,
         new_AGEMA_signal_2391, new_AGEMA_signal_2390, new_AGEMA_signal_2497,
         new_AGEMA_signal_2496, new_AGEMA_signal_4521, new_AGEMA_signal_4519,
         new_AGEMA_signal_4517, new_AGEMA_signal_2199, new_AGEMA_signal_2198,
         SubCellInst_SboxInst_5_T1, new_AGEMA_signal_2307,
         new_AGEMA_signal_2306, SubCellInst_SboxInst_5_L0,
         new_AGEMA_signal_4533, new_AGEMA_signal_4531, new_AGEMA_signal_4529,
         new_AGEMA_signal_2201, new_AGEMA_signal_2200,
         SubCellInst_SboxInst_5_T3, new_AGEMA_signal_2393,
         new_AGEMA_signal_2392, SubCellInst_SboxInst_5_YY_3,
         new_AGEMA_signal_4551, new_AGEMA_signal_4547, new_AGEMA_signal_4543,
         new_AGEMA_signal_2395, new_AGEMA_signal_2394, new_AGEMA_signal_2499,
         new_AGEMA_signal_2498, new_AGEMA_signal_4557, new_AGEMA_signal_4555,
         new_AGEMA_signal_4553, new_AGEMA_signal_2207, new_AGEMA_signal_2206,
         SubCellInst_SboxInst_6_T1, new_AGEMA_signal_2311,
         new_AGEMA_signal_2310, SubCellInst_SboxInst_6_L0,
         new_AGEMA_signal_4569, new_AGEMA_signal_4567, new_AGEMA_signal_4565,
         new_AGEMA_signal_2209, new_AGEMA_signal_2208,
         SubCellInst_SboxInst_6_T3, new_AGEMA_signal_2397,
         new_AGEMA_signal_2396, SubCellInst_SboxInst_6_YY_3,
         new_AGEMA_signal_4587, new_AGEMA_signal_4583, new_AGEMA_signal_4579,
         new_AGEMA_signal_2399, new_AGEMA_signal_2398, new_AGEMA_signal_2501,
         new_AGEMA_signal_2500, new_AGEMA_signal_4593, new_AGEMA_signal_4591,
         new_AGEMA_signal_4589, new_AGEMA_signal_2215, new_AGEMA_signal_2214,
         SubCellInst_SboxInst_7_T1, new_AGEMA_signal_2315,
         new_AGEMA_signal_2314, SubCellInst_SboxInst_7_L0,
         new_AGEMA_signal_4605, new_AGEMA_signal_4603, new_AGEMA_signal_4601,
         new_AGEMA_signal_2217, new_AGEMA_signal_2216,
         SubCellInst_SboxInst_7_T3, new_AGEMA_signal_2401,
         new_AGEMA_signal_2400, SubCellInst_SboxInst_7_YY_3,
         new_AGEMA_signal_4623, new_AGEMA_signal_4619, new_AGEMA_signal_4615,
         new_AGEMA_signal_2403, new_AGEMA_signal_2402, new_AGEMA_signal_4629,
         new_AGEMA_signal_4627, new_AGEMA_signal_4625, new_AGEMA_signal_2223,
         new_AGEMA_signal_2222, SubCellInst_SboxInst_8_T1,
         new_AGEMA_signal_2319, new_AGEMA_signal_2318,
         SubCellInst_SboxInst_8_L0, new_AGEMA_signal_4641,
         new_AGEMA_signal_4639, new_AGEMA_signal_4637, new_AGEMA_signal_2225,
         new_AGEMA_signal_2224, SubCellInst_SboxInst_8_T3,
         new_AGEMA_signal_2405, new_AGEMA_signal_2404,
         SubCellInst_SboxInst_8_YY_3, new_AGEMA_signal_4659,
         new_AGEMA_signal_4655, new_AGEMA_signal_4651, new_AGEMA_signal_2407,
         new_AGEMA_signal_2406, new_AGEMA_signal_2505, new_AGEMA_signal_2504,
         new_AGEMA_signal_4665, new_AGEMA_signal_4663, new_AGEMA_signal_4661,
         new_AGEMA_signal_2231, new_AGEMA_signal_2230,
         SubCellInst_SboxInst_9_T1, new_AGEMA_signal_2323,
         new_AGEMA_signal_2322, SubCellInst_SboxInst_9_L0,
         new_AGEMA_signal_4677, new_AGEMA_signal_4675, new_AGEMA_signal_4673,
         new_AGEMA_signal_2233, new_AGEMA_signal_2232,
         SubCellInst_SboxInst_9_T3, new_AGEMA_signal_2409,
         new_AGEMA_signal_2408, SubCellInst_SboxInst_9_YY_3,
         new_AGEMA_signal_4695, new_AGEMA_signal_4691, new_AGEMA_signal_4687,
         new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2507,
         new_AGEMA_signal_2506, new_AGEMA_signal_4701, new_AGEMA_signal_4699,
         new_AGEMA_signal_4697, new_AGEMA_signal_2239, new_AGEMA_signal_2238,
         SubCellInst_SboxInst_10_T1, new_AGEMA_signal_2327,
         new_AGEMA_signal_2326, SubCellInst_SboxInst_10_L0,
         new_AGEMA_signal_4713, new_AGEMA_signal_4711, new_AGEMA_signal_4709,
         new_AGEMA_signal_2241, new_AGEMA_signal_2240,
         SubCellInst_SboxInst_10_T3, new_AGEMA_signal_2413,
         new_AGEMA_signal_2412, SubCellInst_SboxInst_10_YY_3,
         new_AGEMA_signal_4731, new_AGEMA_signal_4727, new_AGEMA_signal_4723,
         new_AGEMA_signal_2415, new_AGEMA_signal_2414, new_AGEMA_signal_2509,
         new_AGEMA_signal_2508, new_AGEMA_signal_4737, new_AGEMA_signal_4735,
         new_AGEMA_signal_4733, new_AGEMA_signal_2247, new_AGEMA_signal_2246,
         SubCellInst_SboxInst_11_T1, new_AGEMA_signal_2331,
         new_AGEMA_signal_2330, SubCellInst_SboxInst_11_L0,
         new_AGEMA_signal_4749, new_AGEMA_signal_4747, new_AGEMA_signal_4745,
         new_AGEMA_signal_2249, new_AGEMA_signal_2248,
         SubCellInst_SboxInst_11_T3, new_AGEMA_signal_2417,
         new_AGEMA_signal_2416, SubCellInst_SboxInst_11_YY_3,
         new_AGEMA_signal_4767, new_AGEMA_signal_4763, new_AGEMA_signal_4759,
         new_AGEMA_signal_2419, new_AGEMA_signal_2418, new_AGEMA_signal_2511,
         new_AGEMA_signal_2510, new_AGEMA_signal_4773, new_AGEMA_signal_4771,
         new_AGEMA_signal_4769, new_AGEMA_signal_2255, new_AGEMA_signal_2254,
         SubCellInst_SboxInst_12_T1, new_AGEMA_signal_2335,
         new_AGEMA_signal_2334, SubCellInst_SboxInst_12_L0,
         new_AGEMA_signal_4785, new_AGEMA_signal_4783, new_AGEMA_signal_4781,
         new_AGEMA_signal_2257, new_AGEMA_signal_2256,
         SubCellInst_SboxInst_12_T3, new_AGEMA_signal_2421,
         new_AGEMA_signal_2420, SubCellInst_SboxInst_12_YY_3,
         new_AGEMA_signal_4803, new_AGEMA_signal_4799, new_AGEMA_signal_4795,
         new_AGEMA_signal_2423, new_AGEMA_signal_2422, new_AGEMA_signal_2513,
         new_AGEMA_signal_2512, new_AGEMA_signal_4809, new_AGEMA_signal_4807,
         new_AGEMA_signal_4805, new_AGEMA_signal_2263, new_AGEMA_signal_2262,
         SubCellInst_SboxInst_13_T1, new_AGEMA_signal_2339,
         new_AGEMA_signal_2338, SubCellInst_SboxInst_13_L0,
         new_AGEMA_signal_4821, new_AGEMA_signal_4819, new_AGEMA_signal_4817,
         new_AGEMA_signal_2265, new_AGEMA_signal_2264,
         SubCellInst_SboxInst_13_T3, new_AGEMA_signal_2425,
         new_AGEMA_signal_2424, SubCellInst_SboxInst_13_YY_3,
         new_AGEMA_signal_4839, new_AGEMA_signal_4835, new_AGEMA_signal_4831,
         new_AGEMA_signal_2427, new_AGEMA_signal_2426, new_AGEMA_signal_2515,
         new_AGEMA_signal_2514, new_AGEMA_signal_4845, new_AGEMA_signal_4843,
         new_AGEMA_signal_4841, new_AGEMA_signal_2271, new_AGEMA_signal_2270,
         SubCellInst_SboxInst_14_T1, new_AGEMA_signal_2343,
         new_AGEMA_signal_2342, SubCellInst_SboxInst_14_L0,
         new_AGEMA_signal_4857, new_AGEMA_signal_4855, new_AGEMA_signal_4853,
         new_AGEMA_signal_2273, new_AGEMA_signal_2272,
         SubCellInst_SboxInst_14_T3, new_AGEMA_signal_2429,
         new_AGEMA_signal_2428, SubCellInst_SboxInst_14_YY_3,
         new_AGEMA_signal_4875, new_AGEMA_signal_4871, new_AGEMA_signal_4867,
         new_AGEMA_signal_2431, new_AGEMA_signal_2430, new_AGEMA_signal_2517,
         new_AGEMA_signal_2516, new_AGEMA_signal_4881, new_AGEMA_signal_4879,
         new_AGEMA_signal_4877, new_AGEMA_signal_2279, new_AGEMA_signal_2278,
         SubCellInst_SboxInst_15_T1, new_AGEMA_signal_2347,
         new_AGEMA_signal_2346, SubCellInst_SboxInst_15_L0,
         new_AGEMA_signal_4893, new_AGEMA_signal_4891, new_AGEMA_signal_4889,
         new_AGEMA_signal_2281, new_AGEMA_signal_2280,
         SubCellInst_SboxInst_15_T3, new_AGEMA_signal_2433,
         new_AGEMA_signal_2432, SubCellInst_SboxInst_15_YY_3,
         new_AGEMA_signal_4911, new_AGEMA_signal_4907, new_AGEMA_signal_4903,
         new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2519,
         new_AGEMA_signal_2518, new_AGEMA_signal_4917, new_AGEMA_signal_4915,
         new_AGEMA_signal_4913, new_AGEMA_signal_2595, new_AGEMA_signal_2594,
         new_AGEMA_signal_2597, new_AGEMA_signal_2596, new_AGEMA_signal_4921,
         new_AGEMA_signal_2521, new_AGEMA_signal_2520,
         AddConstXOR_AddConstXOR_XORInst_0_0_n1, new_AGEMA_signal_2731,
         new_AGEMA_signal_2730, new_AGEMA_signal_4925, new_AGEMA_signal_2599,
         new_AGEMA_signal_2598, AddConstXOR_AddConstXOR_XORInst_0_1_n1,
         new_AGEMA_signal_2601, new_AGEMA_signal_2600, new_AGEMA_signal_4929,
         new_AGEMA_signal_2525, new_AGEMA_signal_2524,
         AddConstXOR_AddConstXOR_XORInst_1_0_n1, new_AGEMA_signal_2733,
         new_AGEMA_signal_2732, new_AGEMA_signal_4933, new_AGEMA_signal_2603,
         new_AGEMA_signal_2602, AddConstXOR_AddConstXOR_XORInst_1_1_n1,
         new_AGEMA_signal_2605, new_AGEMA_signal_2604, new_AGEMA_signal_4945,
         new_AGEMA_signal_4941, new_AGEMA_signal_4937, new_AGEMA_signal_2529,
         new_AGEMA_signal_2528, AddRoundTweakeyXOR_XORInst_0_0_n1,
         new_AGEMA_signal_2735, new_AGEMA_signal_2734, new_AGEMA_signal_4957,
         new_AGEMA_signal_4953, new_AGEMA_signal_4949, new_AGEMA_signal_2607,
         new_AGEMA_signal_2606, AddRoundTweakeyXOR_XORInst_0_1_n1,
         new_AGEMA_signal_2609, new_AGEMA_signal_2608, new_AGEMA_signal_4969,
         new_AGEMA_signal_4965, new_AGEMA_signal_4961, new_AGEMA_signal_2533,
         new_AGEMA_signal_2532, AddRoundTweakeyXOR_XORInst_1_0_n1,
         new_AGEMA_signal_2737, new_AGEMA_signal_2736, new_AGEMA_signal_4981,
         new_AGEMA_signal_4977, new_AGEMA_signal_4973, new_AGEMA_signal_2611,
         new_AGEMA_signal_2610, AddRoundTweakeyXOR_XORInst_1_1_n1,
         new_AGEMA_signal_2613, new_AGEMA_signal_2612, new_AGEMA_signal_4993,
         new_AGEMA_signal_4989, new_AGEMA_signal_4985, new_AGEMA_signal_2537,
         new_AGEMA_signal_2536, AddRoundTweakeyXOR_XORInst_2_0_n1,
         new_AGEMA_signal_2739, new_AGEMA_signal_2738, new_AGEMA_signal_5005,
         new_AGEMA_signal_5001, new_AGEMA_signal_4997, new_AGEMA_signal_2615,
         new_AGEMA_signal_2614, AddRoundTweakeyXOR_XORInst_2_1_n1,
         new_AGEMA_signal_2851, new_AGEMA_signal_2850, new_AGEMA_signal_5017,
         new_AGEMA_signal_5013, new_AGEMA_signal_5009, new_AGEMA_signal_2741,
         new_AGEMA_signal_2740, AddRoundTweakeyXOR_XORInst_3_0_n1,
         new_AGEMA_signal_2959, new_AGEMA_signal_2958, new_AGEMA_signal_5029,
         new_AGEMA_signal_5025, new_AGEMA_signal_5021, new_AGEMA_signal_2853,
         new_AGEMA_signal_2852, AddRoundTweakeyXOR_XORInst_3_1_n1,
         new_AGEMA_signal_5041, new_AGEMA_signal_5037, new_AGEMA_signal_5033,
         new_AGEMA_signal_2543, new_AGEMA_signal_2542,
         AddRoundTweakeyXOR_XORInst_4_0_n1, new_AGEMA_signal_5053,
         new_AGEMA_signal_5049, new_AGEMA_signal_5045, new_AGEMA_signal_2623,
         new_AGEMA_signal_2622, AddRoundTweakeyXOR_XORInst_4_1_n1,
         new_AGEMA_signal_5065, new_AGEMA_signal_5061, new_AGEMA_signal_5057,
         new_AGEMA_signal_2547, new_AGEMA_signal_2546,
         AddRoundTweakeyXOR_XORInst_5_0_n1, new_AGEMA_signal_5077,
         new_AGEMA_signal_5073, new_AGEMA_signal_5069, new_AGEMA_signal_2627,
         new_AGEMA_signal_2626, AddRoundTweakeyXOR_XORInst_5_1_n1,
         new_AGEMA_signal_5089, new_AGEMA_signal_5085, new_AGEMA_signal_5081,
         new_AGEMA_signal_2551, new_AGEMA_signal_2550,
         AddRoundTweakeyXOR_XORInst_6_0_n1, new_AGEMA_signal_5101,
         new_AGEMA_signal_5097, new_AGEMA_signal_5093, new_AGEMA_signal_2631,
         new_AGEMA_signal_2630, AddRoundTweakeyXOR_XORInst_6_1_n1,
         new_AGEMA_signal_5113, new_AGEMA_signal_5109, new_AGEMA_signal_5105,
         new_AGEMA_signal_2751, new_AGEMA_signal_2750,
         AddRoundTweakeyXOR_XORInst_7_0_n1, new_AGEMA_signal_5125,
         new_AGEMA_signal_5121, new_AGEMA_signal_5117, new_AGEMA_signal_2857,
         new_AGEMA_signal_2856, AddRoundTweakeyXOR_XORInst_7_1_n1,
         new_AGEMA_signal_2557, new_AGEMA_signal_2556,
         MCInst_MCR0_XORInst_0_0_n1, new_AGEMA_signal_2755,
         new_AGEMA_signal_2754, MCInst_MCR0_XORInst_0_0_n2,
         new_AGEMA_signal_2637, new_AGEMA_signal_2636,
         MCInst_MCR0_XORInst_0_1_n1, new_AGEMA_signal_2861,
         new_AGEMA_signal_2860, MCInst_MCR0_XORInst_0_1_n2,
         new_AGEMA_signal_2561, new_AGEMA_signal_2560,
         MCInst_MCR0_XORInst_1_0_n1, new_AGEMA_signal_2759,
         new_AGEMA_signal_2758, MCInst_MCR0_XORInst_1_0_n2,
         new_AGEMA_signal_2761, new_AGEMA_signal_2760,
         MCInst_MCR0_XORInst_1_1_n1, new_AGEMA_signal_2865,
         new_AGEMA_signal_2864, MCInst_MCR0_XORInst_1_1_n2,
         new_AGEMA_signal_2565, new_AGEMA_signal_2564,
         MCInst_MCR0_XORInst_2_0_n1, new_AGEMA_signal_2765,
         new_AGEMA_signal_2764, MCInst_MCR0_XORInst_2_0_n2,
         new_AGEMA_signal_2647, new_AGEMA_signal_2646,
         MCInst_MCR0_XORInst_2_1_n1, new_AGEMA_signal_2869,
         new_AGEMA_signal_2868, MCInst_MCR0_XORInst_2_1_n2,
         new_AGEMA_signal_2569, new_AGEMA_signal_2568,
         MCInst_MCR0_XORInst_3_0_n1, new_AGEMA_signal_2969,
         new_AGEMA_signal_2968, MCInst_MCR0_XORInst_3_0_n2,
         new_AGEMA_signal_2653, new_AGEMA_signal_2652,
         MCInst_MCR0_XORInst_3_1_n1, new_AGEMA_signal_3047,
         new_AGEMA_signal_3046, MCInst_MCR0_XORInst_3_1_n2,
         new_AGEMA_signal_2771, new_AGEMA_signal_2770,
         MCInst_MCR2_XORInst_0_0_n1, new_AGEMA_signal_2877,
         new_AGEMA_signal_2876, MCInst_MCR2_XORInst_0_1_n1,
         new_AGEMA_signal_2775, new_AGEMA_signal_2774,
         MCInst_MCR2_XORInst_1_0_n1, new_AGEMA_signal_2881,
         new_AGEMA_signal_2880, MCInst_MCR2_XORInst_1_1_n1,
         new_AGEMA_signal_2977, new_AGEMA_signal_2976,
         MCInst_MCR2_XORInst_2_0_n1, new_AGEMA_signal_3051,
         new_AGEMA_signal_3050, MCInst_MCR2_XORInst_2_1_n1,
         new_AGEMA_signal_2781, new_AGEMA_signal_2780,
         MCInst_MCR2_XORInst_3_0_n1, new_AGEMA_signal_2889,
         new_AGEMA_signal_2888, MCInst_MCR2_XORInst_3_1_n1,
         new_AGEMA_signal_2785, new_AGEMA_signal_2784,
         MCInst_MCR3_XORInst_0_0_n1, new_AGEMA_signal_2893,
         new_AGEMA_signal_2892, MCInst_MCR3_XORInst_0_1_n1,
         new_AGEMA_signal_2789, new_AGEMA_signal_2788,
         MCInst_MCR3_XORInst_1_0_n1, new_AGEMA_signal_2897,
         new_AGEMA_signal_2896, MCInst_MCR3_XORInst_1_1_n1,
         new_AGEMA_signal_2793, new_AGEMA_signal_2792,
         MCInst_MCR3_XORInst_2_0_n1, new_AGEMA_signal_2901,
         new_AGEMA_signal_2900, MCInst_MCR3_XORInst_2_1_n1,
         new_AGEMA_signal_2989, new_AGEMA_signal_2988,
         MCInst_MCR3_XORInst_3_0_n1, new_AGEMA_signal_3055,
         new_AGEMA_signal_3054, MCInst_MCR3_XORInst_3_1_n1,
         new_AGEMA_signal_5127, new_AGEMA_signal_5129, new_AGEMA_signal_5131,
         new_AGEMA_signal_5133, new_AGEMA_signal_5135, new_AGEMA_signal_5137,
         new_AGEMA_signal_5139, new_AGEMA_signal_5141, new_AGEMA_signal_5143,
         new_AGEMA_signal_5145, new_AGEMA_signal_5147, new_AGEMA_signal_5149,
         new_AGEMA_signal_5151, new_AGEMA_signal_5153, new_AGEMA_signal_5155,
         new_AGEMA_signal_5157, new_AGEMA_signal_5159, new_AGEMA_signal_5161,
         new_AGEMA_signal_5163, new_AGEMA_signal_5165, new_AGEMA_signal_5167,
         new_AGEMA_signal_5169, new_AGEMA_signal_5171, new_AGEMA_signal_5173,
         new_AGEMA_signal_5175, new_AGEMA_signal_5177, new_AGEMA_signal_5179,
         new_AGEMA_signal_5181, new_AGEMA_signal_5183, new_AGEMA_signal_5185,
         new_AGEMA_signal_5187, new_AGEMA_signal_5189, new_AGEMA_signal_5191,
         new_AGEMA_signal_5193, new_AGEMA_signal_5195, new_AGEMA_signal_5197,
         new_AGEMA_signal_5199, new_AGEMA_signal_5201, new_AGEMA_signal_5203,
         new_AGEMA_signal_5205, new_AGEMA_signal_5207, new_AGEMA_signal_5209,
         new_AGEMA_signal_5211, new_AGEMA_signal_5213, new_AGEMA_signal_5215,
         new_AGEMA_signal_5217, new_AGEMA_signal_5219, new_AGEMA_signal_5221,
         new_AGEMA_signal_5223, new_AGEMA_signal_5225, new_AGEMA_signal_5227,
         new_AGEMA_signal_5229, new_AGEMA_signal_5231, new_AGEMA_signal_5233,
         new_AGEMA_signal_5235, new_AGEMA_signal_5237, new_AGEMA_signal_5239,
         new_AGEMA_signal_5241, new_AGEMA_signal_5243, new_AGEMA_signal_5245,
         new_AGEMA_signal_5247, new_AGEMA_signal_5249, new_AGEMA_signal_5251,
         new_AGEMA_signal_5253, new_AGEMA_signal_5255, new_AGEMA_signal_5257,
         new_AGEMA_signal_5259, new_AGEMA_signal_5261, new_AGEMA_signal_5263,
         new_AGEMA_signal_5265, new_AGEMA_signal_5267, new_AGEMA_signal_5269,
         new_AGEMA_signal_5271, new_AGEMA_signal_5273, new_AGEMA_signal_5275,
         new_AGEMA_signal_5277, new_AGEMA_signal_5279, new_AGEMA_signal_5281,
         new_AGEMA_signal_5283, new_AGEMA_signal_5285, new_AGEMA_signal_5287,
         new_AGEMA_signal_5289, new_AGEMA_signal_5291, new_AGEMA_signal_5293,
         new_AGEMA_signal_5295, new_AGEMA_signal_5297, new_AGEMA_signal_5299,
         new_AGEMA_signal_5301, new_AGEMA_signal_5303, new_AGEMA_signal_5305,
         new_AGEMA_signal_5307, new_AGEMA_signal_5309, new_AGEMA_signal_5311,
         new_AGEMA_signal_5313, new_AGEMA_signal_5315, new_AGEMA_signal_5317,
         new_AGEMA_signal_5321, new_AGEMA_signal_5325, new_AGEMA_signal_5329,
         new_AGEMA_signal_5333, new_AGEMA_signal_5337, new_AGEMA_signal_5341,
         new_AGEMA_signal_5345, new_AGEMA_signal_5349, new_AGEMA_signal_5353,
         new_AGEMA_signal_5357, new_AGEMA_signal_5361, new_AGEMA_signal_5365,
         new_AGEMA_signal_5369, new_AGEMA_signal_5373, new_AGEMA_signal_5377,
         new_AGEMA_signal_5381, new_AGEMA_signal_5385, new_AGEMA_signal_5389,
         new_AGEMA_signal_5393, new_AGEMA_signal_5397, new_AGEMA_signal_5401,
         new_AGEMA_signal_5405, new_AGEMA_signal_5409, new_AGEMA_signal_5413,
         new_AGEMA_signal_5417, new_AGEMA_signal_5421, new_AGEMA_signal_5425,
         new_AGEMA_signal_5429, new_AGEMA_signal_5433, new_AGEMA_signal_5437,
         new_AGEMA_signal_5441, new_AGEMA_signal_5445, new_AGEMA_signal_5449,
         new_AGEMA_signal_5453, new_AGEMA_signal_5457, new_AGEMA_signal_5461,
         new_AGEMA_signal_5465, new_AGEMA_signal_5469, new_AGEMA_signal_5473,
         new_AGEMA_signal_5477, new_AGEMA_signal_5481, new_AGEMA_signal_5485,
         new_AGEMA_signal_5489, new_AGEMA_signal_5493, new_AGEMA_signal_5497,
         new_AGEMA_signal_5501, new_AGEMA_signal_5505, new_AGEMA_signal_5509,
         new_AGEMA_signal_5513, new_AGEMA_signal_5517, new_AGEMA_signal_5521,
         new_AGEMA_signal_5525, new_AGEMA_signal_5529, new_AGEMA_signal_5533,
         new_AGEMA_signal_5537, new_AGEMA_signal_5541, new_AGEMA_signal_5545,
         new_AGEMA_signal_5549, new_AGEMA_signal_5553, new_AGEMA_signal_5557,
         new_AGEMA_signal_5561, new_AGEMA_signal_5565, new_AGEMA_signal_5569,
         new_AGEMA_signal_5573, new_AGEMA_signal_5577, new_AGEMA_signal_5581,
         new_AGEMA_signal_5585, new_AGEMA_signal_5589, new_AGEMA_signal_5593,
         new_AGEMA_signal_5597, new_AGEMA_signal_5601, new_AGEMA_signal_5605,
         new_AGEMA_signal_5609, new_AGEMA_signal_5613, new_AGEMA_signal_5617,
         new_AGEMA_signal_5621, new_AGEMA_signal_5625, new_AGEMA_signal_5629,
         new_AGEMA_signal_5633, new_AGEMA_signal_5637, new_AGEMA_signal_5641,
         new_AGEMA_signal_5645, new_AGEMA_signal_5649, new_AGEMA_signal_5653,
         new_AGEMA_signal_5657, new_AGEMA_signal_5661, new_AGEMA_signal_5665,
         new_AGEMA_signal_5669, new_AGEMA_signal_5673, new_AGEMA_signal_5677,
         new_AGEMA_signal_5681, new_AGEMA_signal_5685, new_AGEMA_signal_5689,
         new_AGEMA_signal_5693, new_AGEMA_signal_5697, new_AGEMA_signal_5701,
         new_AGEMA_signal_5705, new_AGEMA_signal_5709, new_AGEMA_signal_5713,
         new_AGEMA_signal_5717, new_AGEMA_signal_5721, new_AGEMA_signal_5725,
         new_AGEMA_signal_5729, new_AGEMA_signal_5733, new_AGEMA_signal_5737,
         new_AGEMA_signal_5741, new_AGEMA_signal_5745, new_AGEMA_signal_5749,
         new_AGEMA_signal_5753, new_AGEMA_signal_5757, new_AGEMA_signal_5761,
         new_AGEMA_signal_5765, new_AGEMA_signal_5769, new_AGEMA_signal_5773,
         new_AGEMA_signal_5777, new_AGEMA_signal_5781, new_AGEMA_signal_5785,
         new_AGEMA_signal_5789, new_AGEMA_signal_5793, new_AGEMA_signal_5797,
         new_AGEMA_signal_5801, new_AGEMA_signal_5805, new_AGEMA_signal_5809,
         new_AGEMA_signal_5813, new_AGEMA_signal_5817, new_AGEMA_signal_5821,
         new_AGEMA_signal_5825, new_AGEMA_signal_5829, new_AGEMA_signal_5833,
         new_AGEMA_signal_5837, new_AGEMA_signal_5841, new_AGEMA_signal_5845,
         new_AGEMA_signal_5849, new_AGEMA_signal_5853, new_AGEMA_signal_5857,
         new_AGEMA_signal_5861, new_AGEMA_signal_5865, new_AGEMA_signal_5869,
         new_AGEMA_signal_5873, new_AGEMA_signal_5877, new_AGEMA_signal_5881,
         new_AGEMA_signal_5885, new_AGEMA_signal_5889, new_AGEMA_signal_5893,
         new_AGEMA_signal_5897, new_AGEMA_signal_5901, new_AGEMA_signal_5905,
         new_AGEMA_signal_5909, new_AGEMA_signal_5913, new_AGEMA_signal_5917,
         new_AGEMA_signal_5921, new_AGEMA_signal_5925, new_AGEMA_signal_5929,
         new_AGEMA_signal_5933, new_AGEMA_signal_5937, new_AGEMA_signal_5941,
         new_AGEMA_signal_5945, new_AGEMA_signal_5949, new_AGEMA_signal_5953,
         new_AGEMA_signal_5957, new_AGEMA_signal_5961, new_AGEMA_signal_5965,
         new_AGEMA_signal_5969, new_AGEMA_signal_5973, new_AGEMA_signal_5977,
         new_AGEMA_signal_5981, new_AGEMA_signal_5985, new_AGEMA_signal_5989,
         new_AGEMA_signal_5993, new_AGEMA_signal_5997, new_AGEMA_signal_6001,
         new_AGEMA_signal_6005, new_AGEMA_signal_6009, new_AGEMA_signal_6013,
         new_AGEMA_signal_6017, new_AGEMA_signal_6021, new_AGEMA_signal_6025,
         new_AGEMA_signal_6029, new_AGEMA_signal_6033, new_AGEMA_signal_6037,
         new_AGEMA_signal_6041, new_AGEMA_signal_6045, new_AGEMA_signal_6049,
         new_AGEMA_signal_6053, new_AGEMA_signal_6057, new_AGEMA_signal_6061,
         new_AGEMA_signal_6065, new_AGEMA_signal_6069, new_AGEMA_signal_6073,
         new_AGEMA_signal_6077, new_AGEMA_signal_6081, new_AGEMA_signal_6085,
         new_AGEMA_signal_6089, new_AGEMA_signal_6093, new_AGEMA_signal_6097,
         new_AGEMA_signal_6101, new_AGEMA_signal_6105, new_AGEMA_signal_6109,
         n13, n14, n15, n16, n17, n18, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56,
         SubCellInst_SboxInst_0_AND1_U1_n36,
         SubCellInst_SboxInst_0_AND1_U1_n35,
         SubCellInst_SboxInst_0_AND1_U1_n34,
         SubCellInst_SboxInst_0_AND1_U1_n33,
         SubCellInst_SboxInst_0_AND1_U1_n32,
         SubCellInst_SboxInst_0_AND1_U1_n31,
         SubCellInst_SboxInst_0_AND1_U1_n30,
         SubCellInst_SboxInst_0_AND1_U1_n29,
         SubCellInst_SboxInst_0_AND1_U1_n28,
         SubCellInst_SboxInst_0_AND1_U1_n27,
         SubCellInst_SboxInst_0_AND1_U1_n26,
         SubCellInst_SboxInst_0_AND1_U1_n25,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_0_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_0_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_0_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_0_AND3_U1_n36,
         SubCellInst_SboxInst_0_AND3_U1_n35,
         SubCellInst_SboxInst_0_AND3_U1_n34,
         SubCellInst_SboxInst_0_AND3_U1_n33,
         SubCellInst_SboxInst_0_AND3_U1_n32,
         SubCellInst_SboxInst_0_AND3_U1_n31,
         SubCellInst_SboxInst_0_AND3_U1_n30,
         SubCellInst_SboxInst_0_AND3_U1_n29,
         SubCellInst_SboxInst_0_AND3_U1_n28,
         SubCellInst_SboxInst_0_AND3_U1_n27,
         SubCellInst_SboxInst_0_AND3_U1_n26,
         SubCellInst_SboxInst_0_AND3_U1_n25,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_0_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_0_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_0_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_1_AND1_U1_n36,
         SubCellInst_SboxInst_1_AND1_U1_n35,
         SubCellInst_SboxInst_1_AND1_U1_n34,
         SubCellInst_SboxInst_1_AND1_U1_n33,
         SubCellInst_SboxInst_1_AND1_U1_n32,
         SubCellInst_SboxInst_1_AND1_U1_n31,
         SubCellInst_SboxInst_1_AND1_U1_n30,
         SubCellInst_SboxInst_1_AND1_U1_n29,
         SubCellInst_SboxInst_1_AND1_U1_n28,
         SubCellInst_SboxInst_1_AND1_U1_n27,
         SubCellInst_SboxInst_1_AND1_U1_n26,
         SubCellInst_SboxInst_1_AND1_U1_n25,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_1_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_1_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_1_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_1_AND3_U1_n36,
         SubCellInst_SboxInst_1_AND3_U1_n35,
         SubCellInst_SboxInst_1_AND3_U1_n34,
         SubCellInst_SboxInst_1_AND3_U1_n33,
         SubCellInst_SboxInst_1_AND3_U1_n32,
         SubCellInst_SboxInst_1_AND3_U1_n31,
         SubCellInst_SboxInst_1_AND3_U1_n30,
         SubCellInst_SboxInst_1_AND3_U1_n29,
         SubCellInst_SboxInst_1_AND3_U1_n28,
         SubCellInst_SboxInst_1_AND3_U1_n27,
         SubCellInst_SboxInst_1_AND3_U1_n26,
         SubCellInst_SboxInst_1_AND3_U1_n25,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_1_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_1_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_1_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_2_AND1_U1_n36,
         SubCellInst_SboxInst_2_AND1_U1_n35,
         SubCellInst_SboxInst_2_AND1_U1_n34,
         SubCellInst_SboxInst_2_AND1_U1_n33,
         SubCellInst_SboxInst_2_AND1_U1_n32,
         SubCellInst_SboxInst_2_AND1_U1_n31,
         SubCellInst_SboxInst_2_AND1_U1_n30,
         SubCellInst_SboxInst_2_AND1_U1_n29,
         SubCellInst_SboxInst_2_AND1_U1_n28,
         SubCellInst_SboxInst_2_AND1_U1_n27,
         SubCellInst_SboxInst_2_AND1_U1_n26,
         SubCellInst_SboxInst_2_AND1_U1_n25,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_2_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_2_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_2_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_2_AND3_U1_n36,
         SubCellInst_SboxInst_2_AND3_U1_n35,
         SubCellInst_SboxInst_2_AND3_U1_n34,
         SubCellInst_SboxInst_2_AND3_U1_n33,
         SubCellInst_SboxInst_2_AND3_U1_n32,
         SubCellInst_SboxInst_2_AND3_U1_n31,
         SubCellInst_SboxInst_2_AND3_U1_n30,
         SubCellInst_SboxInst_2_AND3_U1_n29,
         SubCellInst_SboxInst_2_AND3_U1_n28,
         SubCellInst_SboxInst_2_AND3_U1_n27,
         SubCellInst_SboxInst_2_AND3_U1_n26,
         SubCellInst_SboxInst_2_AND3_U1_n25,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_2_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_2_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_2_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_3_AND1_U1_n36,
         SubCellInst_SboxInst_3_AND1_U1_n35,
         SubCellInst_SboxInst_3_AND1_U1_n34,
         SubCellInst_SboxInst_3_AND1_U1_n33,
         SubCellInst_SboxInst_3_AND1_U1_n32,
         SubCellInst_SboxInst_3_AND1_U1_n31,
         SubCellInst_SboxInst_3_AND1_U1_n30,
         SubCellInst_SboxInst_3_AND1_U1_n29,
         SubCellInst_SboxInst_3_AND1_U1_n28,
         SubCellInst_SboxInst_3_AND1_U1_n27,
         SubCellInst_SboxInst_3_AND1_U1_n26,
         SubCellInst_SboxInst_3_AND1_U1_n25,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_3_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_3_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_3_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_3_AND3_U1_n36,
         SubCellInst_SboxInst_3_AND3_U1_n35,
         SubCellInst_SboxInst_3_AND3_U1_n34,
         SubCellInst_SboxInst_3_AND3_U1_n33,
         SubCellInst_SboxInst_3_AND3_U1_n32,
         SubCellInst_SboxInst_3_AND3_U1_n31,
         SubCellInst_SboxInst_3_AND3_U1_n30,
         SubCellInst_SboxInst_3_AND3_U1_n29,
         SubCellInst_SboxInst_3_AND3_U1_n28,
         SubCellInst_SboxInst_3_AND3_U1_n27,
         SubCellInst_SboxInst_3_AND3_U1_n26,
         SubCellInst_SboxInst_3_AND3_U1_n25,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_3_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_3_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_3_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_4_AND1_U1_n36,
         SubCellInst_SboxInst_4_AND1_U1_n35,
         SubCellInst_SboxInst_4_AND1_U1_n34,
         SubCellInst_SboxInst_4_AND1_U1_n33,
         SubCellInst_SboxInst_4_AND1_U1_n32,
         SubCellInst_SboxInst_4_AND1_U1_n31,
         SubCellInst_SboxInst_4_AND1_U1_n30,
         SubCellInst_SboxInst_4_AND1_U1_n29,
         SubCellInst_SboxInst_4_AND1_U1_n28,
         SubCellInst_SboxInst_4_AND1_U1_n27,
         SubCellInst_SboxInst_4_AND1_U1_n26,
         SubCellInst_SboxInst_4_AND1_U1_n25,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_4_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_4_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_4_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_4_AND3_U1_n36,
         SubCellInst_SboxInst_4_AND3_U1_n35,
         SubCellInst_SboxInst_4_AND3_U1_n34,
         SubCellInst_SboxInst_4_AND3_U1_n33,
         SubCellInst_SboxInst_4_AND3_U1_n32,
         SubCellInst_SboxInst_4_AND3_U1_n31,
         SubCellInst_SboxInst_4_AND3_U1_n30,
         SubCellInst_SboxInst_4_AND3_U1_n29,
         SubCellInst_SboxInst_4_AND3_U1_n28,
         SubCellInst_SboxInst_4_AND3_U1_n27,
         SubCellInst_SboxInst_4_AND3_U1_n26,
         SubCellInst_SboxInst_4_AND3_U1_n25,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_4_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_4_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_4_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_5_AND1_U1_n36,
         SubCellInst_SboxInst_5_AND1_U1_n35,
         SubCellInst_SboxInst_5_AND1_U1_n34,
         SubCellInst_SboxInst_5_AND1_U1_n33,
         SubCellInst_SboxInst_5_AND1_U1_n32,
         SubCellInst_SboxInst_5_AND1_U1_n31,
         SubCellInst_SboxInst_5_AND1_U1_n30,
         SubCellInst_SboxInst_5_AND1_U1_n29,
         SubCellInst_SboxInst_5_AND1_U1_n28,
         SubCellInst_SboxInst_5_AND1_U1_n27,
         SubCellInst_SboxInst_5_AND1_U1_n26,
         SubCellInst_SboxInst_5_AND1_U1_n25,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_5_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_5_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_5_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_5_AND3_U1_n36,
         SubCellInst_SboxInst_5_AND3_U1_n35,
         SubCellInst_SboxInst_5_AND3_U1_n34,
         SubCellInst_SboxInst_5_AND3_U1_n33,
         SubCellInst_SboxInst_5_AND3_U1_n32,
         SubCellInst_SboxInst_5_AND3_U1_n31,
         SubCellInst_SboxInst_5_AND3_U1_n30,
         SubCellInst_SboxInst_5_AND3_U1_n29,
         SubCellInst_SboxInst_5_AND3_U1_n28,
         SubCellInst_SboxInst_5_AND3_U1_n27,
         SubCellInst_SboxInst_5_AND3_U1_n26,
         SubCellInst_SboxInst_5_AND3_U1_n25,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_5_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_5_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_5_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_6_AND1_U1_n36,
         SubCellInst_SboxInst_6_AND1_U1_n35,
         SubCellInst_SboxInst_6_AND1_U1_n34,
         SubCellInst_SboxInst_6_AND1_U1_n33,
         SubCellInst_SboxInst_6_AND1_U1_n32,
         SubCellInst_SboxInst_6_AND1_U1_n31,
         SubCellInst_SboxInst_6_AND1_U1_n30,
         SubCellInst_SboxInst_6_AND1_U1_n29,
         SubCellInst_SboxInst_6_AND1_U1_n28,
         SubCellInst_SboxInst_6_AND1_U1_n27,
         SubCellInst_SboxInst_6_AND1_U1_n26,
         SubCellInst_SboxInst_6_AND1_U1_n25,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_6_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_6_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_6_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_6_AND3_U1_n36,
         SubCellInst_SboxInst_6_AND3_U1_n35,
         SubCellInst_SboxInst_6_AND3_U1_n34,
         SubCellInst_SboxInst_6_AND3_U1_n33,
         SubCellInst_SboxInst_6_AND3_U1_n32,
         SubCellInst_SboxInst_6_AND3_U1_n31,
         SubCellInst_SboxInst_6_AND3_U1_n30,
         SubCellInst_SboxInst_6_AND3_U1_n29,
         SubCellInst_SboxInst_6_AND3_U1_n28,
         SubCellInst_SboxInst_6_AND3_U1_n27,
         SubCellInst_SboxInst_6_AND3_U1_n26,
         SubCellInst_SboxInst_6_AND3_U1_n25,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_6_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_6_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_6_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_7_AND1_U1_n36,
         SubCellInst_SboxInst_7_AND1_U1_n35,
         SubCellInst_SboxInst_7_AND1_U1_n34,
         SubCellInst_SboxInst_7_AND1_U1_n33,
         SubCellInst_SboxInst_7_AND1_U1_n32,
         SubCellInst_SboxInst_7_AND1_U1_n31,
         SubCellInst_SboxInst_7_AND1_U1_n30,
         SubCellInst_SboxInst_7_AND1_U1_n29,
         SubCellInst_SboxInst_7_AND1_U1_n28,
         SubCellInst_SboxInst_7_AND1_U1_n27,
         SubCellInst_SboxInst_7_AND1_U1_n26,
         SubCellInst_SboxInst_7_AND1_U1_n25,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_7_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_7_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_7_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_7_AND3_U1_n36,
         SubCellInst_SboxInst_7_AND3_U1_n35,
         SubCellInst_SboxInst_7_AND3_U1_n34,
         SubCellInst_SboxInst_7_AND3_U1_n33,
         SubCellInst_SboxInst_7_AND3_U1_n32,
         SubCellInst_SboxInst_7_AND3_U1_n31,
         SubCellInst_SboxInst_7_AND3_U1_n30,
         SubCellInst_SboxInst_7_AND3_U1_n29,
         SubCellInst_SboxInst_7_AND3_U1_n28,
         SubCellInst_SboxInst_7_AND3_U1_n27,
         SubCellInst_SboxInst_7_AND3_U1_n26,
         SubCellInst_SboxInst_7_AND3_U1_n25,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_7_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_7_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_7_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_8_AND1_U1_n36,
         SubCellInst_SboxInst_8_AND1_U1_n35,
         SubCellInst_SboxInst_8_AND1_U1_n34,
         SubCellInst_SboxInst_8_AND1_U1_n33,
         SubCellInst_SboxInst_8_AND1_U1_n32,
         SubCellInst_SboxInst_8_AND1_U1_n31,
         SubCellInst_SboxInst_8_AND1_U1_n30,
         SubCellInst_SboxInst_8_AND1_U1_n29,
         SubCellInst_SboxInst_8_AND1_U1_n28,
         SubCellInst_SboxInst_8_AND1_U1_n27,
         SubCellInst_SboxInst_8_AND1_U1_n26,
         SubCellInst_SboxInst_8_AND1_U1_n25,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_8_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_8_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_8_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_8_AND3_U1_n36,
         SubCellInst_SboxInst_8_AND3_U1_n35,
         SubCellInst_SboxInst_8_AND3_U1_n34,
         SubCellInst_SboxInst_8_AND3_U1_n33,
         SubCellInst_SboxInst_8_AND3_U1_n32,
         SubCellInst_SboxInst_8_AND3_U1_n31,
         SubCellInst_SboxInst_8_AND3_U1_n30,
         SubCellInst_SboxInst_8_AND3_U1_n29,
         SubCellInst_SboxInst_8_AND3_U1_n28,
         SubCellInst_SboxInst_8_AND3_U1_n27,
         SubCellInst_SboxInst_8_AND3_U1_n26,
         SubCellInst_SboxInst_8_AND3_U1_n25,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_8_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_8_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_8_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_9_AND1_U1_n36,
         SubCellInst_SboxInst_9_AND1_U1_n35,
         SubCellInst_SboxInst_9_AND1_U1_n34,
         SubCellInst_SboxInst_9_AND1_U1_n33,
         SubCellInst_SboxInst_9_AND1_U1_n32,
         SubCellInst_SboxInst_9_AND1_U1_n31,
         SubCellInst_SboxInst_9_AND1_U1_n30,
         SubCellInst_SboxInst_9_AND1_U1_n29,
         SubCellInst_SboxInst_9_AND1_U1_n28,
         SubCellInst_SboxInst_9_AND1_U1_n27,
         SubCellInst_SboxInst_9_AND1_U1_n26,
         SubCellInst_SboxInst_9_AND1_U1_n25,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_9_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_9_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_9_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_9_AND3_U1_n36,
         SubCellInst_SboxInst_9_AND3_U1_n35,
         SubCellInst_SboxInst_9_AND3_U1_n34,
         SubCellInst_SboxInst_9_AND3_U1_n33,
         SubCellInst_SboxInst_9_AND3_U1_n32,
         SubCellInst_SboxInst_9_AND3_U1_n31,
         SubCellInst_SboxInst_9_AND3_U1_n30,
         SubCellInst_SboxInst_9_AND3_U1_n29,
         SubCellInst_SboxInst_9_AND3_U1_n28,
         SubCellInst_SboxInst_9_AND3_U1_n27,
         SubCellInst_SboxInst_9_AND3_U1_n26,
         SubCellInst_SboxInst_9_AND3_U1_n25,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_9_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_9_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_9_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_10_AND1_U1_n36,
         SubCellInst_SboxInst_10_AND1_U1_n35,
         SubCellInst_SboxInst_10_AND1_U1_n34,
         SubCellInst_SboxInst_10_AND1_U1_n33,
         SubCellInst_SboxInst_10_AND1_U1_n32,
         SubCellInst_SboxInst_10_AND1_U1_n31,
         SubCellInst_SboxInst_10_AND1_U1_n30,
         SubCellInst_SboxInst_10_AND1_U1_n29,
         SubCellInst_SboxInst_10_AND1_U1_n28,
         SubCellInst_SboxInst_10_AND1_U1_n27,
         SubCellInst_SboxInst_10_AND1_U1_n26,
         SubCellInst_SboxInst_10_AND1_U1_n25,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_10_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_10_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_10_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_10_AND3_U1_n36,
         SubCellInst_SboxInst_10_AND3_U1_n35,
         SubCellInst_SboxInst_10_AND3_U1_n34,
         SubCellInst_SboxInst_10_AND3_U1_n33,
         SubCellInst_SboxInst_10_AND3_U1_n32,
         SubCellInst_SboxInst_10_AND3_U1_n31,
         SubCellInst_SboxInst_10_AND3_U1_n30,
         SubCellInst_SboxInst_10_AND3_U1_n29,
         SubCellInst_SboxInst_10_AND3_U1_n28,
         SubCellInst_SboxInst_10_AND3_U1_n27,
         SubCellInst_SboxInst_10_AND3_U1_n26,
         SubCellInst_SboxInst_10_AND3_U1_n25,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_10_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_10_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_10_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_11_AND1_U1_n36,
         SubCellInst_SboxInst_11_AND1_U1_n35,
         SubCellInst_SboxInst_11_AND1_U1_n34,
         SubCellInst_SboxInst_11_AND1_U1_n33,
         SubCellInst_SboxInst_11_AND1_U1_n32,
         SubCellInst_SboxInst_11_AND1_U1_n31,
         SubCellInst_SboxInst_11_AND1_U1_n30,
         SubCellInst_SboxInst_11_AND1_U1_n29,
         SubCellInst_SboxInst_11_AND1_U1_n28,
         SubCellInst_SboxInst_11_AND1_U1_n27,
         SubCellInst_SboxInst_11_AND1_U1_n26,
         SubCellInst_SboxInst_11_AND1_U1_n25,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_11_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_11_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_11_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_11_AND3_U1_n36,
         SubCellInst_SboxInst_11_AND3_U1_n35,
         SubCellInst_SboxInst_11_AND3_U1_n34,
         SubCellInst_SboxInst_11_AND3_U1_n33,
         SubCellInst_SboxInst_11_AND3_U1_n32,
         SubCellInst_SboxInst_11_AND3_U1_n31,
         SubCellInst_SboxInst_11_AND3_U1_n30,
         SubCellInst_SboxInst_11_AND3_U1_n29,
         SubCellInst_SboxInst_11_AND3_U1_n28,
         SubCellInst_SboxInst_11_AND3_U1_n27,
         SubCellInst_SboxInst_11_AND3_U1_n26,
         SubCellInst_SboxInst_11_AND3_U1_n25,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_11_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_11_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_11_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_12_AND1_U1_n36,
         SubCellInst_SboxInst_12_AND1_U1_n35,
         SubCellInst_SboxInst_12_AND1_U1_n34,
         SubCellInst_SboxInst_12_AND1_U1_n33,
         SubCellInst_SboxInst_12_AND1_U1_n32,
         SubCellInst_SboxInst_12_AND1_U1_n31,
         SubCellInst_SboxInst_12_AND1_U1_n30,
         SubCellInst_SboxInst_12_AND1_U1_n29,
         SubCellInst_SboxInst_12_AND1_U1_n28,
         SubCellInst_SboxInst_12_AND1_U1_n27,
         SubCellInst_SboxInst_12_AND1_U1_n26,
         SubCellInst_SboxInst_12_AND1_U1_n25,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_12_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_12_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_12_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_12_AND3_U1_n36,
         SubCellInst_SboxInst_12_AND3_U1_n35,
         SubCellInst_SboxInst_12_AND3_U1_n34,
         SubCellInst_SboxInst_12_AND3_U1_n33,
         SubCellInst_SboxInst_12_AND3_U1_n32,
         SubCellInst_SboxInst_12_AND3_U1_n31,
         SubCellInst_SboxInst_12_AND3_U1_n30,
         SubCellInst_SboxInst_12_AND3_U1_n29,
         SubCellInst_SboxInst_12_AND3_U1_n28,
         SubCellInst_SboxInst_12_AND3_U1_n27,
         SubCellInst_SboxInst_12_AND3_U1_n26,
         SubCellInst_SboxInst_12_AND3_U1_n25,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_12_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_12_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_12_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_13_AND1_U1_n36,
         SubCellInst_SboxInst_13_AND1_U1_n35,
         SubCellInst_SboxInst_13_AND1_U1_n34,
         SubCellInst_SboxInst_13_AND1_U1_n33,
         SubCellInst_SboxInst_13_AND1_U1_n32,
         SubCellInst_SboxInst_13_AND1_U1_n31,
         SubCellInst_SboxInst_13_AND1_U1_n30,
         SubCellInst_SboxInst_13_AND1_U1_n29,
         SubCellInst_SboxInst_13_AND1_U1_n28,
         SubCellInst_SboxInst_13_AND1_U1_n27,
         SubCellInst_SboxInst_13_AND1_U1_n26,
         SubCellInst_SboxInst_13_AND1_U1_n25,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_13_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_13_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_13_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_13_AND3_U1_n36,
         SubCellInst_SboxInst_13_AND3_U1_n35,
         SubCellInst_SboxInst_13_AND3_U1_n34,
         SubCellInst_SboxInst_13_AND3_U1_n33,
         SubCellInst_SboxInst_13_AND3_U1_n32,
         SubCellInst_SboxInst_13_AND3_U1_n31,
         SubCellInst_SboxInst_13_AND3_U1_n30,
         SubCellInst_SboxInst_13_AND3_U1_n29,
         SubCellInst_SboxInst_13_AND3_U1_n28,
         SubCellInst_SboxInst_13_AND3_U1_n27,
         SubCellInst_SboxInst_13_AND3_U1_n26,
         SubCellInst_SboxInst_13_AND3_U1_n25,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_13_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_13_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_13_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_14_AND1_U1_n36,
         SubCellInst_SboxInst_14_AND1_U1_n35,
         SubCellInst_SboxInst_14_AND1_U1_n34,
         SubCellInst_SboxInst_14_AND1_U1_n33,
         SubCellInst_SboxInst_14_AND1_U1_n32,
         SubCellInst_SboxInst_14_AND1_U1_n31,
         SubCellInst_SboxInst_14_AND1_U1_n30,
         SubCellInst_SboxInst_14_AND1_U1_n29,
         SubCellInst_SboxInst_14_AND1_U1_n28,
         SubCellInst_SboxInst_14_AND1_U1_n27,
         SubCellInst_SboxInst_14_AND1_U1_n26,
         SubCellInst_SboxInst_14_AND1_U1_n25,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_14_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_14_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_14_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_14_AND3_U1_n36,
         SubCellInst_SboxInst_14_AND3_U1_n35,
         SubCellInst_SboxInst_14_AND3_U1_n34,
         SubCellInst_SboxInst_14_AND3_U1_n33,
         SubCellInst_SboxInst_14_AND3_U1_n32,
         SubCellInst_SboxInst_14_AND3_U1_n31,
         SubCellInst_SboxInst_14_AND3_U1_n30,
         SubCellInst_SboxInst_14_AND3_U1_n29,
         SubCellInst_SboxInst_14_AND3_U1_n28,
         SubCellInst_SboxInst_14_AND3_U1_n27,
         SubCellInst_SboxInst_14_AND3_U1_n26,
         SubCellInst_SboxInst_14_AND3_U1_n25,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_14_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_14_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_14_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_15_AND1_U1_n36,
         SubCellInst_SboxInst_15_AND1_U1_n35,
         SubCellInst_SboxInst_15_AND1_U1_n34,
         SubCellInst_SboxInst_15_AND1_U1_n33,
         SubCellInst_SboxInst_15_AND1_U1_n32,
         SubCellInst_SboxInst_15_AND1_U1_n31,
         SubCellInst_SboxInst_15_AND1_U1_n30,
         SubCellInst_SboxInst_15_AND1_U1_n29,
         SubCellInst_SboxInst_15_AND1_U1_n28,
         SubCellInst_SboxInst_15_AND1_U1_n27,
         SubCellInst_SboxInst_15_AND1_U1_n26,
         SubCellInst_SboxInst_15_AND1_U1_n25,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_0__2_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_1__2_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_2__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_2__1_,
         SubCellInst_SboxInst_15_AND1_U1_a_reg_0_,
         SubCellInst_SboxInst_15_AND1_U1_a_reg_1_,
         SubCellInst_SboxInst_15_AND1_U1_a_reg_2_,
         SubCellInst_SboxInst_15_AND3_U1_n36,
         SubCellInst_SboxInst_15_AND3_U1_n35,
         SubCellInst_SboxInst_15_AND3_U1_n34,
         SubCellInst_SboxInst_15_AND3_U1_n33,
         SubCellInst_SboxInst_15_AND3_U1_n32,
         SubCellInst_SboxInst_15_AND3_U1_n31,
         SubCellInst_SboxInst_15_AND3_U1_n30,
         SubCellInst_SboxInst_15_AND3_U1_n29,
         SubCellInst_SboxInst_15_AND3_U1_n28,
         SubCellInst_SboxInst_15_AND3_U1_n27,
         SubCellInst_SboxInst_15_AND3_U1_n26,
         SubCellInst_SboxInst_15_AND3_U1_n25,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_0__2_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_1__2_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_2__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_2__1_,
         SubCellInst_SboxInst_15_AND3_U1_a_reg_0_,
         SubCellInst_SboxInst_15_AND3_U1_a_reg_1_,
         SubCellInst_SboxInst_15_AND3_U1_a_reg_2_,
         SubCellInst_SboxInst_0_AND2_U1_n36,
         SubCellInst_SboxInst_0_AND2_U1_n35,
         SubCellInst_SboxInst_0_AND2_U1_n34,
         SubCellInst_SboxInst_0_AND2_U1_n33,
         SubCellInst_SboxInst_0_AND2_U1_n32,
         SubCellInst_SboxInst_0_AND2_U1_n31,
         SubCellInst_SboxInst_0_AND2_U1_n30,
         SubCellInst_SboxInst_0_AND2_U1_n29,
         SubCellInst_SboxInst_0_AND2_U1_n28,
         SubCellInst_SboxInst_0_AND2_U1_n27,
         SubCellInst_SboxInst_0_AND2_U1_n26,
         SubCellInst_SboxInst_0_AND2_U1_n25,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_0_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_0_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_0_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_0_AND4_U1_n36,
         SubCellInst_SboxInst_0_AND4_U1_n35,
         SubCellInst_SboxInst_0_AND4_U1_n34,
         SubCellInst_SboxInst_0_AND4_U1_n33,
         SubCellInst_SboxInst_0_AND4_U1_n32,
         SubCellInst_SboxInst_0_AND4_U1_n31,
         SubCellInst_SboxInst_0_AND4_U1_n30,
         SubCellInst_SboxInst_0_AND4_U1_n29,
         SubCellInst_SboxInst_0_AND4_U1_n28,
         SubCellInst_SboxInst_0_AND4_U1_n27,
         SubCellInst_SboxInst_0_AND4_U1_n26,
         SubCellInst_SboxInst_0_AND4_U1_n25,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_0_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_0_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_0_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_1_AND2_U1_n36,
         SubCellInst_SboxInst_1_AND2_U1_n35,
         SubCellInst_SboxInst_1_AND2_U1_n34,
         SubCellInst_SboxInst_1_AND2_U1_n33,
         SubCellInst_SboxInst_1_AND2_U1_n32,
         SubCellInst_SboxInst_1_AND2_U1_n31,
         SubCellInst_SboxInst_1_AND2_U1_n30,
         SubCellInst_SboxInst_1_AND2_U1_n29,
         SubCellInst_SboxInst_1_AND2_U1_n28,
         SubCellInst_SboxInst_1_AND2_U1_n27,
         SubCellInst_SboxInst_1_AND2_U1_n26,
         SubCellInst_SboxInst_1_AND2_U1_n25,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_1_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_1_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_1_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_1_AND4_U1_n36,
         SubCellInst_SboxInst_1_AND4_U1_n35,
         SubCellInst_SboxInst_1_AND4_U1_n34,
         SubCellInst_SboxInst_1_AND4_U1_n33,
         SubCellInst_SboxInst_1_AND4_U1_n32,
         SubCellInst_SboxInst_1_AND4_U1_n31,
         SubCellInst_SboxInst_1_AND4_U1_n30,
         SubCellInst_SboxInst_1_AND4_U1_n29,
         SubCellInst_SboxInst_1_AND4_U1_n28,
         SubCellInst_SboxInst_1_AND4_U1_n27,
         SubCellInst_SboxInst_1_AND4_U1_n26,
         SubCellInst_SboxInst_1_AND4_U1_n25,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_1_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_1_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_1_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_2_AND2_U1_n36,
         SubCellInst_SboxInst_2_AND2_U1_n35,
         SubCellInst_SboxInst_2_AND2_U1_n34,
         SubCellInst_SboxInst_2_AND2_U1_n33,
         SubCellInst_SboxInst_2_AND2_U1_n32,
         SubCellInst_SboxInst_2_AND2_U1_n31,
         SubCellInst_SboxInst_2_AND2_U1_n30,
         SubCellInst_SboxInst_2_AND2_U1_n29,
         SubCellInst_SboxInst_2_AND2_U1_n28,
         SubCellInst_SboxInst_2_AND2_U1_n27,
         SubCellInst_SboxInst_2_AND2_U1_n26,
         SubCellInst_SboxInst_2_AND2_U1_n25,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_2_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_2_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_2_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_2_AND4_U1_n36,
         SubCellInst_SboxInst_2_AND4_U1_n35,
         SubCellInst_SboxInst_2_AND4_U1_n34,
         SubCellInst_SboxInst_2_AND4_U1_n33,
         SubCellInst_SboxInst_2_AND4_U1_n32,
         SubCellInst_SboxInst_2_AND4_U1_n31,
         SubCellInst_SboxInst_2_AND4_U1_n30,
         SubCellInst_SboxInst_2_AND4_U1_n29,
         SubCellInst_SboxInst_2_AND4_U1_n28,
         SubCellInst_SboxInst_2_AND4_U1_n27,
         SubCellInst_SboxInst_2_AND4_U1_n26,
         SubCellInst_SboxInst_2_AND4_U1_n25,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_2_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_2_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_2_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_3_AND2_U1_n36,
         SubCellInst_SboxInst_3_AND2_U1_n35,
         SubCellInst_SboxInst_3_AND2_U1_n34,
         SubCellInst_SboxInst_3_AND2_U1_n33,
         SubCellInst_SboxInst_3_AND2_U1_n32,
         SubCellInst_SboxInst_3_AND2_U1_n31,
         SubCellInst_SboxInst_3_AND2_U1_n30,
         SubCellInst_SboxInst_3_AND2_U1_n29,
         SubCellInst_SboxInst_3_AND2_U1_n28,
         SubCellInst_SboxInst_3_AND2_U1_n27,
         SubCellInst_SboxInst_3_AND2_U1_n26,
         SubCellInst_SboxInst_3_AND2_U1_n25,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_3_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_3_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_3_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_3_AND4_U1_n36,
         SubCellInst_SboxInst_3_AND4_U1_n35,
         SubCellInst_SboxInst_3_AND4_U1_n34,
         SubCellInst_SboxInst_3_AND4_U1_n33,
         SubCellInst_SboxInst_3_AND4_U1_n32,
         SubCellInst_SboxInst_3_AND4_U1_n31,
         SubCellInst_SboxInst_3_AND4_U1_n30,
         SubCellInst_SboxInst_3_AND4_U1_n29,
         SubCellInst_SboxInst_3_AND4_U1_n28,
         SubCellInst_SboxInst_3_AND4_U1_n27,
         SubCellInst_SboxInst_3_AND4_U1_n26,
         SubCellInst_SboxInst_3_AND4_U1_n25,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_3_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_3_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_3_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_4_AND2_U1_n36,
         SubCellInst_SboxInst_4_AND2_U1_n35,
         SubCellInst_SboxInst_4_AND2_U1_n34,
         SubCellInst_SboxInst_4_AND2_U1_n33,
         SubCellInst_SboxInst_4_AND2_U1_n32,
         SubCellInst_SboxInst_4_AND2_U1_n31,
         SubCellInst_SboxInst_4_AND2_U1_n30,
         SubCellInst_SboxInst_4_AND2_U1_n29,
         SubCellInst_SboxInst_4_AND2_U1_n28,
         SubCellInst_SboxInst_4_AND2_U1_n27,
         SubCellInst_SboxInst_4_AND2_U1_n26,
         SubCellInst_SboxInst_4_AND2_U1_n25,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_4_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_4_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_4_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_4_AND4_U1_n36,
         SubCellInst_SboxInst_4_AND4_U1_n35,
         SubCellInst_SboxInst_4_AND4_U1_n34,
         SubCellInst_SboxInst_4_AND4_U1_n33,
         SubCellInst_SboxInst_4_AND4_U1_n32,
         SubCellInst_SboxInst_4_AND4_U1_n31,
         SubCellInst_SboxInst_4_AND4_U1_n30,
         SubCellInst_SboxInst_4_AND4_U1_n29,
         SubCellInst_SboxInst_4_AND4_U1_n28,
         SubCellInst_SboxInst_4_AND4_U1_n27,
         SubCellInst_SboxInst_4_AND4_U1_n26,
         SubCellInst_SboxInst_4_AND4_U1_n25,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_4_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_4_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_4_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_5_AND2_U1_n36,
         SubCellInst_SboxInst_5_AND2_U1_n35,
         SubCellInst_SboxInst_5_AND2_U1_n34,
         SubCellInst_SboxInst_5_AND2_U1_n33,
         SubCellInst_SboxInst_5_AND2_U1_n32,
         SubCellInst_SboxInst_5_AND2_U1_n31,
         SubCellInst_SboxInst_5_AND2_U1_n30,
         SubCellInst_SboxInst_5_AND2_U1_n29,
         SubCellInst_SboxInst_5_AND2_U1_n28,
         SubCellInst_SboxInst_5_AND2_U1_n27,
         SubCellInst_SboxInst_5_AND2_U1_n26,
         SubCellInst_SboxInst_5_AND2_U1_n25,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_5_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_5_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_5_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_5_AND4_U1_n36,
         SubCellInst_SboxInst_5_AND4_U1_n35,
         SubCellInst_SboxInst_5_AND4_U1_n34,
         SubCellInst_SboxInst_5_AND4_U1_n33,
         SubCellInst_SboxInst_5_AND4_U1_n32,
         SubCellInst_SboxInst_5_AND4_U1_n31,
         SubCellInst_SboxInst_5_AND4_U1_n30,
         SubCellInst_SboxInst_5_AND4_U1_n29,
         SubCellInst_SboxInst_5_AND4_U1_n28,
         SubCellInst_SboxInst_5_AND4_U1_n27,
         SubCellInst_SboxInst_5_AND4_U1_n26,
         SubCellInst_SboxInst_5_AND4_U1_n25,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_5_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_5_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_5_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_6_AND2_U1_n36,
         SubCellInst_SboxInst_6_AND2_U1_n35,
         SubCellInst_SboxInst_6_AND2_U1_n34,
         SubCellInst_SboxInst_6_AND2_U1_n33,
         SubCellInst_SboxInst_6_AND2_U1_n32,
         SubCellInst_SboxInst_6_AND2_U1_n31,
         SubCellInst_SboxInst_6_AND2_U1_n30,
         SubCellInst_SboxInst_6_AND2_U1_n29,
         SubCellInst_SboxInst_6_AND2_U1_n28,
         SubCellInst_SboxInst_6_AND2_U1_n27,
         SubCellInst_SboxInst_6_AND2_U1_n26,
         SubCellInst_SboxInst_6_AND2_U1_n25,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_6_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_6_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_6_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_6_AND4_U1_n36,
         SubCellInst_SboxInst_6_AND4_U1_n35,
         SubCellInst_SboxInst_6_AND4_U1_n34,
         SubCellInst_SboxInst_6_AND4_U1_n33,
         SubCellInst_SboxInst_6_AND4_U1_n32,
         SubCellInst_SboxInst_6_AND4_U1_n31,
         SubCellInst_SboxInst_6_AND4_U1_n30,
         SubCellInst_SboxInst_6_AND4_U1_n29,
         SubCellInst_SboxInst_6_AND4_U1_n28,
         SubCellInst_SboxInst_6_AND4_U1_n27,
         SubCellInst_SboxInst_6_AND4_U1_n26,
         SubCellInst_SboxInst_6_AND4_U1_n25,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_6_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_6_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_6_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_7_AND2_U1_n36,
         SubCellInst_SboxInst_7_AND2_U1_n35,
         SubCellInst_SboxInst_7_AND2_U1_n34,
         SubCellInst_SboxInst_7_AND2_U1_n33,
         SubCellInst_SboxInst_7_AND2_U1_n32,
         SubCellInst_SboxInst_7_AND2_U1_n31,
         SubCellInst_SboxInst_7_AND2_U1_n30,
         SubCellInst_SboxInst_7_AND2_U1_n29,
         SubCellInst_SboxInst_7_AND2_U1_n28,
         SubCellInst_SboxInst_7_AND2_U1_n27,
         SubCellInst_SboxInst_7_AND2_U1_n26,
         SubCellInst_SboxInst_7_AND2_U1_n25,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_7_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_7_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_7_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_7_AND4_U1_n36,
         SubCellInst_SboxInst_7_AND4_U1_n35,
         SubCellInst_SboxInst_7_AND4_U1_n34,
         SubCellInst_SboxInst_7_AND4_U1_n33,
         SubCellInst_SboxInst_7_AND4_U1_n32,
         SubCellInst_SboxInst_7_AND4_U1_n31,
         SubCellInst_SboxInst_7_AND4_U1_n30,
         SubCellInst_SboxInst_7_AND4_U1_n29,
         SubCellInst_SboxInst_7_AND4_U1_n28,
         SubCellInst_SboxInst_7_AND4_U1_n27,
         SubCellInst_SboxInst_7_AND4_U1_n26,
         SubCellInst_SboxInst_7_AND4_U1_n25,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_7_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_7_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_7_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_8_AND2_U1_n36,
         SubCellInst_SboxInst_8_AND2_U1_n35,
         SubCellInst_SboxInst_8_AND2_U1_n34,
         SubCellInst_SboxInst_8_AND2_U1_n33,
         SubCellInst_SboxInst_8_AND2_U1_n32,
         SubCellInst_SboxInst_8_AND2_U1_n31,
         SubCellInst_SboxInst_8_AND2_U1_n30,
         SubCellInst_SboxInst_8_AND2_U1_n29,
         SubCellInst_SboxInst_8_AND2_U1_n28,
         SubCellInst_SboxInst_8_AND2_U1_n27,
         SubCellInst_SboxInst_8_AND2_U1_n26,
         SubCellInst_SboxInst_8_AND2_U1_n25,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_8_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_8_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_8_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_8_AND4_U1_n36,
         SubCellInst_SboxInst_8_AND4_U1_n35,
         SubCellInst_SboxInst_8_AND4_U1_n34,
         SubCellInst_SboxInst_8_AND4_U1_n33,
         SubCellInst_SboxInst_8_AND4_U1_n32,
         SubCellInst_SboxInst_8_AND4_U1_n31,
         SubCellInst_SboxInst_8_AND4_U1_n30,
         SubCellInst_SboxInst_8_AND4_U1_n29,
         SubCellInst_SboxInst_8_AND4_U1_n28,
         SubCellInst_SboxInst_8_AND4_U1_n27,
         SubCellInst_SboxInst_8_AND4_U1_n26,
         SubCellInst_SboxInst_8_AND4_U1_n25,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_8_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_8_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_8_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_9_AND2_U1_n36,
         SubCellInst_SboxInst_9_AND2_U1_n35,
         SubCellInst_SboxInst_9_AND2_U1_n34,
         SubCellInst_SboxInst_9_AND2_U1_n33,
         SubCellInst_SboxInst_9_AND2_U1_n32,
         SubCellInst_SboxInst_9_AND2_U1_n31,
         SubCellInst_SboxInst_9_AND2_U1_n30,
         SubCellInst_SboxInst_9_AND2_U1_n29,
         SubCellInst_SboxInst_9_AND2_U1_n28,
         SubCellInst_SboxInst_9_AND2_U1_n27,
         SubCellInst_SboxInst_9_AND2_U1_n26,
         SubCellInst_SboxInst_9_AND2_U1_n25,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_9_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_9_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_9_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_9_AND4_U1_n36,
         SubCellInst_SboxInst_9_AND4_U1_n35,
         SubCellInst_SboxInst_9_AND4_U1_n34,
         SubCellInst_SboxInst_9_AND4_U1_n33,
         SubCellInst_SboxInst_9_AND4_U1_n32,
         SubCellInst_SboxInst_9_AND4_U1_n31,
         SubCellInst_SboxInst_9_AND4_U1_n30,
         SubCellInst_SboxInst_9_AND4_U1_n29,
         SubCellInst_SboxInst_9_AND4_U1_n28,
         SubCellInst_SboxInst_9_AND4_U1_n27,
         SubCellInst_SboxInst_9_AND4_U1_n26,
         SubCellInst_SboxInst_9_AND4_U1_n25,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_9_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_9_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_9_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_10_AND2_U1_n36,
         SubCellInst_SboxInst_10_AND2_U1_n35,
         SubCellInst_SboxInst_10_AND2_U1_n34,
         SubCellInst_SboxInst_10_AND2_U1_n33,
         SubCellInst_SboxInst_10_AND2_U1_n32,
         SubCellInst_SboxInst_10_AND2_U1_n31,
         SubCellInst_SboxInst_10_AND2_U1_n30,
         SubCellInst_SboxInst_10_AND2_U1_n29,
         SubCellInst_SboxInst_10_AND2_U1_n28,
         SubCellInst_SboxInst_10_AND2_U1_n27,
         SubCellInst_SboxInst_10_AND2_U1_n26,
         SubCellInst_SboxInst_10_AND2_U1_n25,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_10_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_10_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_10_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_10_AND4_U1_n36,
         SubCellInst_SboxInst_10_AND4_U1_n35,
         SubCellInst_SboxInst_10_AND4_U1_n34,
         SubCellInst_SboxInst_10_AND4_U1_n33,
         SubCellInst_SboxInst_10_AND4_U1_n32,
         SubCellInst_SboxInst_10_AND4_U1_n31,
         SubCellInst_SboxInst_10_AND4_U1_n30,
         SubCellInst_SboxInst_10_AND4_U1_n29,
         SubCellInst_SboxInst_10_AND4_U1_n28,
         SubCellInst_SboxInst_10_AND4_U1_n27,
         SubCellInst_SboxInst_10_AND4_U1_n26,
         SubCellInst_SboxInst_10_AND4_U1_n25,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_10_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_10_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_10_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_11_AND2_U1_n36,
         SubCellInst_SboxInst_11_AND2_U1_n35,
         SubCellInst_SboxInst_11_AND2_U1_n34,
         SubCellInst_SboxInst_11_AND2_U1_n33,
         SubCellInst_SboxInst_11_AND2_U1_n32,
         SubCellInst_SboxInst_11_AND2_U1_n31,
         SubCellInst_SboxInst_11_AND2_U1_n30,
         SubCellInst_SboxInst_11_AND2_U1_n29,
         SubCellInst_SboxInst_11_AND2_U1_n28,
         SubCellInst_SboxInst_11_AND2_U1_n27,
         SubCellInst_SboxInst_11_AND2_U1_n26,
         SubCellInst_SboxInst_11_AND2_U1_n25,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_11_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_11_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_11_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_11_AND4_U1_n36,
         SubCellInst_SboxInst_11_AND4_U1_n35,
         SubCellInst_SboxInst_11_AND4_U1_n34,
         SubCellInst_SboxInst_11_AND4_U1_n33,
         SubCellInst_SboxInst_11_AND4_U1_n32,
         SubCellInst_SboxInst_11_AND4_U1_n31,
         SubCellInst_SboxInst_11_AND4_U1_n30,
         SubCellInst_SboxInst_11_AND4_U1_n29,
         SubCellInst_SboxInst_11_AND4_U1_n28,
         SubCellInst_SboxInst_11_AND4_U1_n27,
         SubCellInst_SboxInst_11_AND4_U1_n26,
         SubCellInst_SboxInst_11_AND4_U1_n25,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_11_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_11_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_11_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_12_AND2_U1_n36,
         SubCellInst_SboxInst_12_AND2_U1_n35,
         SubCellInst_SboxInst_12_AND2_U1_n34,
         SubCellInst_SboxInst_12_AND2_U1_n33,
         SubCellInst_SboxInst_12_AND2_U1_n32,
         SubCellInst_SboxInst_12_AND2_U1_n31,
         SubCellInst_SboxInst_12_AND2_U1_n30,
         SubCellInst_SboxInst_12_AND2_U1_n29,
         SubCellInst_SboxInst_12_AND2_U1_n28,
         SubCellInst_SboxInst_12_AND2_U1_n27,
         SubCellInst_SboxInst_12_AND2_U1_n26,
         SubCellInst_SboxInst_12_AND2_U1_n25,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_12_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_12_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_12_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_12_AND4_U1_n36,
         SubCellInst_SboxInst_12_AND4_U1_n35,
         SubCellInst_SboxInst_12_AND4_U1_n34,
         SubCellInst_SboxInst_12_AND4_U1_n33,
         SubCellInst_SboxInst_12_AND4_U1_n32,
         SubCellInst_SboxInst_12_AND4_U1_n31,
         SubCellInst_SboxInst_12_AND4_U1_n30,
         SubCellInst_SboxInst_12_AND4_U1_n29,
         SubCellInst_SboxInst_12_AND4_U1_n28,
         SubCellInst_SboxInst_12_AND4_U1_n27,
         SubCellInst_SboxInst_12_AND4_U1_n26,
         SubCellInst_SboxInst_12_AND4_U1_n25,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_12_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_12_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_12_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_13_AND2_U1_n36,
         SubCellInst_SboxInst_13_AND2_U1_n35,
         SubCellInst_SboxInst_13_AND2_U1_n34,
         SubCellInst_SboxInst_13_AND2_U1_n33,
         SubCellInst_SboxInst_13_AND2_U1_n32,
         SubCellInst_SboxInst_13_AND2_U1_n31,
         SubCellInst_SboxInst_13_AND2_U1_n30,
         SubCellInst_SboxInst_13_AND2_U1_n29,
         SubCellInst_SboxInst_13_AND2_U1_n28,
         SubCellInst_SboxInst_13_AND2_U1_n27,
         SubCellInst_SboxInst_13_AND2_U1_n26,
         SubCellInst_SboxInst_13_AND2_U1_n25,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_13_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_13_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_13_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_13_AND4_U1_n36,
         SubCellInst_SboxInst_13_AND4_U1_n35,
         SubCellInst_SboxInst_13_AND4_U1_n34,
         SubCellInst_SboxInst_13_AND4_U1_n33,
         SubCellInst_SboxInst_13_AND4_U1_n32,
         SubCellInst_SboxInst_13_AND4_U1_n31,
         SubCellInst_SboxInst_13_AND4_U1_n30,
         SubCellInst_SboxInst_13_AND4_U1_n29,
         SubCellInst_SboxInst_13_AND4_U1_n28,
         SubCellInst_SboxInst_13_AND4_U1_n27,
         SubCellInst_SboxInst_13_AND4_U1_n26,
         SubCellInst_SboxInst_13_AND4_U1_n25,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_13_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_13_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_13_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_14_AND2_U1_n36,
         SubCellInst_SboxInst_14_AND2_U1_n35,
         SubCellInst_SboxInst_14_AND2_U1_n34,
         SubCellInst_SboxInst_14_AND2_U1_n33,
         SubCellInst_SboxInst_14_AND2_U1_n32,
         SubCellInst_SboxInst_14_AND2_U1_n31,
         SubCellInst_SboxInst_14_AND2_U1_n30,
         SubCellInst_SboxInst_14_AND2_U1_n29,
         SubCellInst_SboxInst_14_AND2_U1_n28,
         SubCellInst_SboxInst_14_AND2_U1_n27,
         SubCellInst_SboxInst_14_AND2_U1_n26,
         SubCellInst_SboxInst_14_AND2_U1_n25,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_14_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_14_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_14_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_14_AND4_U1_n36,
         SubCellInst_SboxInst_14_AND4_U1_n35,
         SubCellInst_SboxInst_14_AND4_U1_n34,
         SubCellInst_SboxInst_14_AND4_U1_n33,
         SubCellInst_SboxInst_14_AND4_U1_n32,
         SubCellInst_SboxInst_14_AND4_U1_n31,
         SubCellInst_SboxInst_14_AND4_U1_n30,
         SubCellInst_SboxInst_14_AND4_U1_n29,
         SubCellInst_SboxInst_14_AND4_U1_n28,
         SubCellInst_SboxInst_14_AND4_U1_n27,
         SubCellInst_SboxInst_14_AND4_U1_n26,
         SubCellInst_SboxInst_14_AND4_U1_n25,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_14_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_14_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_14_AND4_U1_a_reg_2_,
         SubCellInst_SboxInst_15_AND2_U1_n36,
         SubCellInst_SboxInst_15_AND2_U1_n35,
         SubCellInst_SboxInst_15_AND2_U1_n34,
         SubCellInst_SboxInst_15_AND2_U1_n33,
         SubCellInst_SboxInst_15_AND2_U1_n32,
         SubCellInst_SboxInst_15_AND2_U1_n31,
         SubCellInst_SboxInst_15_AND2_U1_n30,
         SubCellInst_SboxInst_15_AND2_U1_n29,
         SubCellInst_SboxInst_15_AND2_U1_n28,
         SubCellInst_SboxInst_15_AND2_U1_n27,
         SubCellInst_SboxInst_15_AND2_U1_n26,
         SubCellInst_SboxInst_15_AND2_U1_n25,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_0__2_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_1__2_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_2__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_2__1_,
         SubCellInst_SboxInst_15_AND2_U1_a_reg_0_,
         SubCellInst_SboxInst_15_AND2_U1_a_reg_1_,
         SubCellInst_SboxInst_15_AND2_U1_a_reg_2_,
         SubCellInst_SboxInst_15_AND4_U1_n36,
         SubCellInst_SboxInst_15_AND4_U1_n35,
         SubCellInst_SboxInst_15_AND4_U1_n34,
         SubCellInst_SboxInst_15_AND4_U1_n33,
         SubCellInst_SboxInst_15_AND4_U1_n32,
         SubCellInst_SboxInst_15_AND4_U1_n31,
         SubCellInst_SboxInst_15_AND4_U1_n30,
         SubCellInst_SboxInst_15_AND4_U1_n29,
         SubCellInst_SboxInst_15_AND4_U1_n28,
         SubCellInst_SboxInst_15_AND4_U1_n27,
         SubCellInst_SboxInst_15_AND4_U1_n26,
         SubCellInst_SboxInst_15_AND4_U1_n25,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_0__2_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_1__2_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_2__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_2__1_,
         SubCellInst_SboxInst_15_AND4_U1_a_reg_0_,
         SubCellInst_SboxInst_15_AND4_U1_a_reg_1_,
         SubCellInst_SboxInst_15_AND4_U1_a_reg_2_;
  wire   [63:0] TweakeyGeneration_StateRegInput;
  wire   [63:0] TweakeyGeneration_key_Feedback;
  wire   [4:1] FSMUpdate;
  wire   [5:0] FSMSelected;
  wire   [5:4] FSM;
  wire   [63:0] StateRegInput;
  wire   [63:0] MCOutput;
  wire   [47:0] ShiftRowsOutput;
  wire   [63:32] AddRoundConstantOutput;
  wire   [63:60] SubCellOutput;
  wire   [2:0] SubCellInst_SboxInst_0_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_0_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_0_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_0_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_0_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_0_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_1_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_1_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_1_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_1_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_1_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_1_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_2_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_2_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_2_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_2_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_2_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_2_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_3_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_3_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_3_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_3_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_3_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_3_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_4_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_4_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_4_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_4_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_4_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_4_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_5_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_5_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_5_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_5_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_5_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_5_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_6_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_6_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_6_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_6_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_6_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_6_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_7_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_7_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_7_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_7_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_7_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_7_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_8_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_8_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_8_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_8_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_8_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_8_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_9_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_9_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_9_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_9_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_9_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_9_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_10_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_10_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_10_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_10_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_10_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_10_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_11_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_11_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_11_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_11_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_11_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_11_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_12_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_12_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_12_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_12_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_12_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_12_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_13_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_13_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_13_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_13_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_13_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_13_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_14_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_14_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_14_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_14_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_14_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_14_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_15_AND1_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_15_AND1_U1_z;
  wire   [2:0] SubCellInst_SboxInst_15_AND1_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_15_AND3_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_15_AND3_U1_z;
  wire   [2:0] SubCellInst_SboxInst_15_AND3_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_0_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_0_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_0_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_0_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_0_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_0_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_1_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_1_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_1_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_1_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_1_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_1_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_2_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_2_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_2_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_2_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_2_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_2_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_3_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_3_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_3_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_3_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_3_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_3_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_4_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_4_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_4_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_4_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_4_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_4_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_5_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_5_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_5_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_5_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_5_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_5_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_6_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_6_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_6_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_6_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_6_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_6_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_7_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_7_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_7_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_7_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_7_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_7_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_8_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_8_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_8_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_8_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_8_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_8_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_9_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_9_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_9_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_9_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_9_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_9_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_10_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_10_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_10_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_10_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_10_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_10_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_11_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_11_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_11_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_11_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_11_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_11_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_12_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_12_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_12_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_12_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_12_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_12_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_13_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_13_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_13_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_13_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_13_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_13_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_14_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_14_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_14_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_14_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_14_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_14_AND4_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_15_AND2_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_15_AND2_U1_z;
  wire   [2:0] SubCellInst_SboxInst_15_AND2_U1_mul;
  wire   [2:0] SubCellInst_SboxInst_15_AND4_U1_mul_s1_out;
  wire   [2:0] SubCellInst_SboxInst_15_AND4_U1_z;
  wire   [2:0] SubCellInst_SboxInst_15_AND4_U1_mul;

  DFF_X1 FSMReg_s_current_state_reg_5__FF_FF ( .D(new_AGEMA_signal_6089), .CK(
        clk), .Q(FSM[5]), .QN(n13) );
  DFF_X1 FSMReg_s_current_state_reg_4__FF_FF ( .D(new_AGEMA_signal_6093), .CK(
        clk), .Q(FSM[4]), .QN(n14) );
  DFF_X1 FSMReg_s_current_state_reg_3__FF_FF ( .D(new_AGEMA_signal_6097), .CK(
        clk), .Q(FSMUpdate[4]), .QN(n16) );
  DFF_X1 FSMReg_s_current_state_reg_2__FF_FF ( .D(new_AGEMA_signal_6101), .CK(
        clk), .Q(FSMUpdate[3]), .QN(n17) );
  DFF_X1 FSMReg_s_current_state_reg_1__FF_FF ( .D(new_AGEMA_signal_6105), .CK(
        clk), .Q(FSM_1), .QN(n15) );
  DFF_X1 FSMReg_s_current_state_reg_0__FF_FF ( .D(new_AGEMA_signal_6109), .CK(
        clk), .Q(FSMUpdate[1]), .QN(n18) );
  BUF_X2 U39 ( .A(new_AGEMA_signal_3279), .Z(n46) );
  BUF_X1 U40 ( .A(new_AGEMA_signal_3957), .Z(n42) );
  BUF_X1 U41 ( .A(new_AGEMA_signal_3957), .Z(n44) );
  BUF_X1 U42 ( .A(new_AGEMA_signal_3957), .Z(n43) );
  BUF_X2 U43 ( .A(new_AGEMA_signal_3279), .Z(n47) );
  BUF_X2 U44 ( .A(new_AGEMA_signal_3279), .Z(n45) );
  BUF_X1 U45 ( .A(new_AGEMA_signal_3957), .Z(n41) );
  BUF_X1 U46 ( .A(new_AGEMA_signal_3957), .Z(n40) );
  INV_X1 U47 ( .A(rst), .ZN(n48) );
  NAND3_X1 U48 ( .A1(n16), .A2(n17), .A3(FSM_1), .ZN(n54) );
  NOR2_X1 U49 ( .A1(n18), .A2(n54), .ZN(n49) );
  OAI21_X1 U50 ( .B1(n13), .B2(n49), .A(n14), .ZN(n50) );
  OAI211_X1 U51 ( .C1(n13), .C2(n14), .A(n48), .B(n50), .ZN(FSMSelected[0]) );
  NOR2_X1 U52 ( .A1(rst), .A2(n18), .ZN(FSMSelected[1]) );
  NOR2_X1 U53 ( .A1(rst), .A2(n16), .ZN(FSMSelected[4]) );
  NOR2_X1 U54 ( .A1(rst), .A2(n17), .ZN(FSMSelected[3]) );
  NOR2_X1 U55 ( .A1(FSMSelected[4]), .A2(FSMSelected[3]), .ZN(n53) );
  NAND2_X1 U56 ( .A1(n14), .A2(FSM[5]), .ZN(n51) );
  OAI21_X1 U57 ( .B1(n18), .B2(n51), .A(n48), .ZN(n52) );
  AOI21_X1 U58 ( .B1(n53), .B2(n52), .A(n15), .ZN(FSMSelected[2]) );
  NAND2_X1 U59 ( .A1(FSMSelected[1]), .A2(FSM[5]), .ZN(n55) );
  OAI22_X1 U60 ( .A1(rst), .A2(n14), .B1(n55), .B2(n54), .ZN(FSMSelected[5])
         );
  NAND4_X1 U61 ( .A1(n15), .A2(n16), .A3(n17), .A4(FSM[5]), .ZN(n56) );
  NOR3_X1 U62 ( .A1(n14), .A2(n18), .A3(n56), .ZN(done) );
  INV_X1 SubCellInst_SboxInst_0_U1_U1 ( .A(Ciphertext_s0[2]), .ZN(
        SubCellInst_SboxInst_0_n3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[2]), 
        .B(Ciphertext_s0[3]), .Z(SubCellInst_SboxInst_0_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[2]), 
        .B(Ciphertext_s1[3]), .Z(new_AGEMA_signal_1170) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[2]), 
        .B(Ciphertext_s2[3]), .Z(new_AGEMA_signal_1171) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[0]), 
        .B(Ciphertext_s0[2]), .Z(SubCellInst_SboxInst_0_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[0]), 
        .B(Ciphertext_s1[2]), .Z(new_AGEMA_signal_1174) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[0]), 
        .B(Ciphertext_s2[2]), .Z(new_AGEMA_signal_1175) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_XX_2_), .Z(SubCellInst_SboxInst_0_Q0) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        new_AGEMA_signal_1174), .Z(new_AGEMA_signal_1742) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[1]), .B(
        new_AGEMA_signal_1175), .Z(new_AGEMA_signal_1743) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_XX_1_), .Z(SubCellInst_SboxInst_0_Q1) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        new_AGEMA_signal_1170), .Z(new_AGEMA_signal_1744) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[1]), .B(
        new_AGEMA_signal_1171), .Z(new_AGEMA_signal_1745) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_n3), .ZN(SubCellInst_SboxInst_0_Q4) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        Ciphertext_s1[2]), .Z(new_AGEMA_signal_1746) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[1]), .B(
        Ciphertext_s2[2]), .Z(new_AGEMA_signal_1747) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_XX_2_), .B(SubCellInst_SboxInst_0_n3), .Z(
        SubCellInst_SboxInst_0_Q6) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1174), 
        .B(Ciphertext_s1[2]), .Z(new_AGEMA_signal_1748) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1175), 
        .B(Ciphertext_s2[2]), .Z(new_AGEMA_signal_1749) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_0_Q1), .B(SubCellInst_SboxInst_0_Q6), .ZN(
        SubCellInst_SboxInst_0_L1) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1744), 
        .B(new_AGEMA_signal_1748), .Z(new_AGEMA_signal_1936) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1745), 
        .B(new_AGEMA_signal_1749), .Z(new_AGEMA_signal_1937) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_n3), .Z(SubCellInst_SboxInst_0_L2) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        Ciphertext_s1[2]), .Z(new_AGEMA_signal_1750) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[1]), .B(
        Ciphertext_s2[2]), .Z(new_AGEMA_signal_1751) );
  INV_X1 SubCellInst_SboxInst_1_U1_U1 ( .A(Ciphertext_s0[6]), .ZN(
        SubCellInst_SboxInst_1_n3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[6]), 
        .B(Ciphertext_s0[7]), .Z(SubCellInst_SboxInst_1_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[6]), 
        .B(Ciphertext_s1[7]), .Z(new_AGEMA_signal_1182) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[6]), 
        .B(Ciphertext_s2[7]), .Z(new_AGEMA_signal_1183) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[4]), 
        .B(Ciphertext_s0[6]), .Z(SubCellInst_SboxInst_1_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[4]), 
        .B(Ciphertext_s1[6]), .Z(new_AGEMA_signal_1186) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[4]), 
        .B(Ciphertext_s2[6]), .Z(new_AGEMA_signal_1187) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_XX_2_), .Z(SubCellInst_SboxInst_1_Q0) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        new_AGEMA_signal_1186), .Z(new_AGEMA_signal_1754) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[5]), .B(
        new_AGEMA_signal_1187), .Z(new_AGEMA_signal_1755) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_XX_1_), .Z(SubCellInst_SboxInst_1_Q1) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        new_AGEMA_signal_1182), .Z(new_AGEMA_signal_1756) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[5]), .B(
        new_AGEMA_signal_1183), .Z(new_AGEMA_signal_1757) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_n3), .ZN(SubCellInst_SboxInst_1_Q4) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        Ciphertext_s1[6]), .Z(new_AGEMA_signal_1758) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[5]), .B(
        Ciphertext_s2[6]), .Z(new_AGEMA_signal_1759) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_XX_2_), .B(SubCellInst_SboxInst_1_n3), .Z(
        SubCellInst_SboxInst_1_Q6) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1186), 
        .B(Ciphertext_s1[6]), .Z(new_AGEMA_signal_1760) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1187), 
        .B(Ciphertext_s2[6]), .Z(new_AGEMA_signal_1761) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_1_Q1), .B(SubCellInst_SboxInst_1_Q6), .ZN(
        SubCellInst_SboxInst_1_L1) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1756), 
        .B(new_AGEMA_signal_1760), .Z(new_AGEMA_signal_1942) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1757), 
        .B(new_AGEMA_signal_1761), .Z(new_AGEMA_signal_1943) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_n3), .Z(SubCellInst_SboxInst_1_L2) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        Ciphertext_s1[6]), .Z(new_AGEMA_signal_1762) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[5]), .B(
        Ciphertext_s2[6]), .Z(new_AGEMA_signal_1763) );
  INV_X1 SubCellInst_SboxInst_2_U1_U1 ( .A(Ciphertext_s0[10]), .ZN(
        SubCellInst_SboxInst_2_n3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[10]), 
        .B(Ciphertext_s0[11]), .Z(SubCellInst_SboxInst_2_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[10]), 
        .B(Ciphertext_s1[11]), .Z(new_AGEMA_signal_1194) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[10]), 
        .B(Ciphertext_s2[11]), .Z(new_AGEMA_signal_1195) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[8]), 
        .B(Ciphertext_s0[10]), .Z(SubCellInst_SboxInst_2_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[8]), 
        .B(Ciphertext_s1[10]), .Z(new_AGEMA_signal_1198) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[8]), 
        .B(Ciphertext_s2[10]), .Z(new_AGEMA_signal_1199) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_XX_2_), .Z(SubCellInst_SboxInst_2_Q0) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        new_AGEMA_signal_1198), .Z(new_AGEMA_signal_1766) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[9]), .B(
        new_AGEMA_signal_1199), .Z(new_AGEMA_signal_1767) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_XX_1_), .Z(SubCellInst_SboxInst_2_Q1) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        new_AGEMA_signal_1194), .Z(new_AGEMA_signal_1768) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[9]), .B(
        new_AGEMA_signal_1195), .Z(new_AGEMA_signal_1769) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_n3), .ZN(SubCellInst_SboxInst_2_Q4) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        Ciphertext_s1[10]), .Z(new_AGEMA_signal_1770) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[9]), .B(
        Ciphertext_s2[10]), .Z(new_AGEMA_signal_1771) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_XX_2_), .B(SubCellInst_SboxInst_2_n3), .Z(
        SubCellInst_SboxInst_2_Q6) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1198), 
        .B(Ciphertext_s1[10]), .Z(new_AGEMA_signal_1772) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1199), 
        .B(Ciphertext_s2[10]), .Z(new_AGEMA_signal_1773) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_2_Q1), .B(SubCellInst_SboxInst_2_Q6), .ZN(
        SubCellInst_SboxInst_2_L1) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1768), 
        .B(new_AGEMA_signal_1772), .Z(new_AGEMA_signal_1948) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1769), 
        .B(new_AGEMA_signal_1773), .Z(new_AGEMA_signal_1949) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_n3), .Z(SubCellInst_SboxInst_2_L2) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        Ciphertext_s1[10]), .Z(new_AGEMA_signal_1774) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[9]), .B(
        Ciphertext_s2[10]), .Z(new_AGEMA_signal_1775) );
  INV_X1 SubCellInst_SboxInst_3_U1_U1 ( .A(Ciphertext_s0[14]), .ZN(
        SubCellInst_SboxInst_3_n3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[14]), 
        .B(Ciphertext_s0[15]), .Z(SubCellInst_SboxInst_3_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[14]), 
        .B(Ciphertext_s1[15]), .Z(new_AGEMA_signal_1206) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[14]), 
        .B(Ciphertext_s2[15]), .Z(new_AGEMA_signal_1207) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[12]), 
        .B(Ciphertext_s0[14]), .Z(SubCellInst_SboxInst_3_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[12]), 
        .B(Ciphertext_s1[14]), .Z(new_AGEMA_signal_1210) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[12]), 
        .B(Ciphertext_s2[14]), .Z(new_AGEMA_signal_1211) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_XX_2_), .Z(SubCellInst_SboxInst_3_Q0) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        new_AGEMA_signal_1210), .Z(new_AGEMA_signal_1778) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[13]), .B(
        new_AGEMA_signal_1211), .Z(new_AGEMA_signal_1779) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_XX_1_), .Z(SubCellInst_SboxInst_3_Q1) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        new_AGEMA_signal_1206), .Z(new_AGEMA_signal_1780) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[13]), .B(
        new_AGEMA_signal_1207), .Z(new_AGEMA_signal_1781) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_n3), .ZN(SubCellInst_SboxInst_3_Q4) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        Ciphertext_s1[14]), .Z(new_AGEMA_signal_1782) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[13]), .B(
        Ciphertext_s2[14]), .Z(new_AGEMA_signal_1783) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_XX_2_), .B(SubCellInst_SboxInst_3_n3), .Z(
        SubCellInst_SboxInst_3_Q6) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1210), 
        .B(Ciphertext_s1[14]), .Z(new_AGEMA_signal_1784) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1211), 
        .B(Ciphertext_s2[14]), .Z(new_AGEMA_signal_1785) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_3_Q1), .B(SubCellInst_SboxInst_3_Q6), .ZN(
        SubCellInst_SboxInst_3_L1) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1780), 
        .B(new_AGEMA_signal_1784), .Z(new_AGEMA_signal_1954) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1781), 
        .B(new_AGEMA_signal_1785), .Z(new_AGEMA_signal_1955) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_n3), .Z(SubCellInst_SboxInst_3_L2) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        Ciphertext_s1[14]), .Z(new_AGEMA_signal_1786) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[13]), .B(
        Ciphertext_s2[14]), .Z(new_AGEMA_signal_1787) );
  INV_X1 SubCellInst_SboxInst_4_U1_U1 ( .A(Ciphertext_s0[18]), .ZN(
        SubCellInst_SboxInst_4_n3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[18]), 
        .B(Ciphertext_s0[19]), .Z(SubCellInst_SboxInst_4_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[18]), 
        .B(Ciphertext_s1[19]), .Z(new_AGEMA_signal_1218) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[18]), 
        .B(Ciphertext_s2[19]), .Z(new_AGEMA_signal_1219) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[16]), 
        .B(Ciphertext_s0[18]), .Z(SubCellInst_SboxInst_4_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[16]), 
        .B(Ciphertext_s1[18]), .Z(new_AGEMA_signal_1222) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[16]), 
        .B(Ciphertext_s2[18]), .Z(new_AGEMA_signal_1223) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_XX_2_), .Z(SubCellInst_SboxInst_4_Q0) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        new_AGEMA_signal_1222), .Z(new_AGEMA_signal_1790) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[17]), .B(
        new_AGEMA_signal_1223), .Z(new_AGEMA_signal_1791) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_XX_1_), .Z(SubCellInst_SboxInst_4_Q1) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        new_AGEMA_signal_1218), .Z(new_AGEMA_signal_1792) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[17]), .B(
        new_AGEMA_signal_1219), .Z(new_AGEMA_signal_1793) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_n3), .ZN(SubCellInst_SboxInst_4_Q4) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        Ciphertext_s1[18]), .Z(new_AGEMA_signal_1794) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[17]), .B(
        Ciphertext_s2[18]), .Z(new_AGEMA_signal_1795) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_XX_2_), .B(SubCellInst_SboxInst_4_n3), .Z(
        SubCellInst_SboxInst_4_Q6) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1222), 
        .B(Ciphertext_s1[18]), .Z(new_AGEMA_signal_1796) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1223), 
        .B(Ciphertext_s2[18]), .Z(new_AGEMA_signal_1797) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_4_Q1), .B(SubCellInst_SboxInst_4_Q6), .ZN(
        SubCellInst_SboxInst_4_L1) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1792), 
        .B(new_AGEMA_signal_1796), .Z(new_AGEMA_signal_1960) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1793), 
        .B(new_AGEMA_signal_1797), .Z(new_AGEMA_signal_1961) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_n3), .Z(SubCellInst_SboxInst_4_L2) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        Ciphertext_s1[18]), .Z(new_AGEMA_signal_1798) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[17]), .B(
        Ciphertext_s2[18]), .Z(new_AGEMA_signal_1799) );
  INV_X1 SubCellInst_SboxInst_5_U1_U1 ( .A(Ciphertext_s0[22]), .ZN(
        SubCellInst_SboxInst_5_n3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[22]), 
        .B(Ciphertext_s0[23]), .Z(SubCellInst_SboxInst_5_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[22]), 
        .B(Ciphertext_s1[23]), .Z(new_AGEMA_signal_1230) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[22]), 
        .B(Ciphertext_s2[23]), .Z(new_AGEMA_signal_1231) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[20]), 
        .B(Ciphertext_s0[22]), .Z(SubCellInst_SboxInst_5_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[20]), 
        .B(Ciphertext_s1[22]), .Z(new_AGEMA_signal_1234) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[20]), 
        .B(Ciphertext_s2[22]), .Z(new_AGEMA_signal_1235) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_XX_2_), .Z(SubCellInst_SboxInst_5_Q0) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        new_AGEMA_signal_1234), .Z(new_AGEMA_signal_1802) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[21]), .B(
        new_AGEMA_signal_1235), .Z(new_AGEMA_signal_1803) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_XX_1_), .Z(SubCellInst_SboxInst_5_Q1) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        new_AGEMA_signal_1230), .Z(new_AGEMA_signal_1804) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[21]), .B(
        new_AGEMA_signal_1231), .Z(new_AGEMA_signal_1805) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_n3), .ZN(SubCellInst_SboxInst_5_Q4) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        Ciphertext_s1[22]), .Z(new_AGEMA_signal_1806) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[21]), .B(
        Ciphertext_s2[22]), .Z(new_AGEMA_signal_1807) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_XX_2_), .B(SubCellInst_SboxInst_5_n3), .Z(
        SubCellInst_SboxInst_5_Q6) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1234), 
        .B(Ciphertext_s1[22]), .Z(new_AGEMA_signal_1808) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1235), 
        .B(Ciphertext_s2[22]), .Z(new_AGEMA_signal_1809) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_5_Q1), .B(SubCellInst_SboxInst_5_Q6), .ZN(
        SubCellInst_SboxInst_5_L1) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1804), 
        .B(new_AGEMA_signal_1808), .Z(new_AGEMA_signal_1966) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1805), 
        .B(new_AGEMA_signal_1809), .Z(new_AGEMA_signal_1967) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_n3), .Z(SubCellInst_SboxInst_5_L2) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        Ciphertext_s1[22]), .Z(new_AGEMA_signal_1810) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[21]), .B(
        Ciphertext_s2[22]), .Z(new_AGEMA_signal_1811) );
  INV_X1 SubCellInst_SboxInst_6_U1_U1 ( .A(Ciphertext_s0[26]), .ZN(
        SubCellInst_SboxInst_6_n3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[26]), 
        .B(Ciphertext_s0[27]), .Z(SubCellInst_SboxInst_6_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[26]), 
        .B(Ciphertext_s1[27]), .Z(new_AGEMA_signal_1242) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[26]), 
        .B(Ciphertext_s2[27]), .Z(new_AGEMA_signal_1243) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[24]), 
        .B(Ciphertext_s0[26]), .Z(SubCellInst_SboxInst_6_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[24]), 
        .B(Ciphertext_s1[26]), .Z(new_AGEMA_signal_1246) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[24]), 
        .B(Ciphertext_s2[26]), .Z(new_AGEMA_signal_1247) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_XX_2_), .Z(SubCellInst_SboxInst_6_Q0) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        new_AGEMA_signal_1246), .Z(new_AGEMA_signal_1814) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[25]), .B(
        new_AGEMA_signal_1247), .Z(new_AGEMA_signal_1815) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_XX_1_), .Z(SubCellInst_SboxInst_6_Q1) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        new_AGEMA_signal_1242), .Z(new_AGEMA_signal_1816) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[25]), .B(
        new_AGEMA_signal_1243), .Z(new_AGEMA_signal_1817) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_n3), .ZN(SubCellInst_SboxInst_6_Q4) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        Ciphertext_s1[26]), .Z(new_AGEMA_signal_1818) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[25]), .B(
        Ciphertext_s2[26]), .Z(new_AGEMA_signal_1819) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_XX_2_), .B(SubCellInst_SboxInst_6_n3), .Z(
        SubCellInst_SboxInst_6_Q6) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1246), 
        .B(Ciphertext_s1[26]), .Z(new_AGEMA_signal_1820) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1247), 
        .B(Ciphertext_s2[26]), .Z(new_AGEMA_signal_1821) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_6_Q1), .B(SubCellInst_SboxInst_6_Q6), .ZN(
        SubCellInst_SboxInst_6_L1) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1816), 
        .B(new_AGEMA_signal_1820), .Z(new_AGEMA_signal_1972) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1817), 
        .B(new_AGEMA_signal_1821), .Z(new_AGEMA_signal_1973) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_n3), .Z(SubCellInst_SboxInst_6_L2) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        Ciphertext_s1[26]), .Z(new_AGEMA_signal_1822) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[25]), .B(
        Ciphertext_s2[26]), .Z(new_AGEMA_signal_1823) );
  INV_X1 SubCellInst_SboxInst_7_U1_U1 ( .A(Ciphertext_s0[30]), .ZN(
        SubCellInst_SboxInst_7_n3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[30]), 
        .B(Ciphertext_s0[31]), .Z(SubCellInst_SboxInst_7_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[30]), 
        .B(Ciphertext_s1[31]), .Z(new_AGEMA_signal_1254) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[30]), 
        .B(Ciphertext_s2[31]), .Z(new_AGEMA_signal_1255) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[28]), 
        .B(Ciphertext_s0[30]), .Z(SubCellInst_SboxInst_7_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[28]), 
        .B(Ciphertext_s1[30]), .Z(new_AGEMA_signal_1258) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[28]), 
        .B(Ciphertext_s2[30]), .Z(new_AGEMA_signal_1259) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_XX_2_), .Z(SubCellInst_SboxInst_7_Q0) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        new_AGEMA_signal_1258), .Z(new_AGEMA_signal_1826) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[29]), .B(
        new_AGEMA_signal_1259), .Z(new_AGEMA_signal_1827) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_XX_1_), .Z(SubCellInst_SboxInst_7_Q1) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        new_AGEMA_signal_1254), .Z(new_AGEMA_signal_1828) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[29]), .B(
        new_AGEMA_signal_1255), .Z(new_AGEMA_signal_1829) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_n3), .ZN(SubCellInst_SboxInst_7_Q4) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        Ciphertext_s1[30]), .Z(new_AGEMA_signal_1830) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[29]), .B(
        Ciphertext_s2[30]), .Z(new_AGEMA_signal_1831) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_XX_2_), .B(SubCellInst_SboxInst_7_n3), .Z(
        SubCellInst_SboxInst_7_Q6) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1258), 
        .B(Ciphertext_s1[30]), .Z(new_AGEMA_signal_1832) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1259), 
        .B(Ciphertext_s2[30]), .Z(new_AGEMA_signal_1833) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_7_Q1), .B(SubCellInst_SboxInst_7_Q6), .ZN(
        SubCellInst_SboxInst_7_L1) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1828), 
        .B(new_AGEMA_signal_1832), .Z(new_AGEMA_signal_1978) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1829), 
        .B(new_AGEMA_signal_1833), .Z(new_AGEMA_signal_1979) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_n3), .Z(SubCellInst_SboxInst_7_L2) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        Ciphertext_s1[30]), .Z(new_AGEMA_signal_1834) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[29]), .B(
        Ciphertext_s2[30]), .Z(new_AGEMA_signal_1835) );
  INV_X1 SubCellInst_SboxInst_8_U1_U1 ( .A(Ciphertext_s0[34]), .ZN(
        SubCellInst_SboxInst_8_n3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[34]), 
        .B(Ciphertext_s0[35]), .Z(SubCellInst_SboxInst_8_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[34]), 
        .B(Ciphertext_s1[35]), .Z(new_AGEMA_signal_1266) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[34]), 
        .B(Ciphertext_s2[35]), .Z(new_AGEMA_signal_1267) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[32]), 
        .B(Ciphertext_s0[34]), .Z(SubCellInst_SboxInst_8_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[32]), 
        .B(Ciphertext_s1[34]), .Z(new_AGEMA_signal_1270) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[32]), 
        .B(Ciphertext_s2[34]), .Z(new_AGEMA_signal_1271) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_XX_2_), .Z(SubCellInst_SboxInst_8_Q0) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        new_AGEMA_signal_1270), .Z(new_AGEMA_signal_1838) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[33]), .B(
        new_AGEMA_signal_1271), .Z(new_AGEMA_signal_1839) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_XX_1_), .Z(SubCellInst_SboxInst_8_Q1) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        new_AGEMA_signal_1266), .Z(new_AGEMA_signal_1840) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[33]), .B(
        new_AGEMA_signal_1267), .Z(new_AGEMA_signal_1841) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_n3), .ZN(SubCellInst_SboxInst_8_Q4) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        Ciphertext_s1[34]), .Z(new_AGEMA_signal_1842) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[33]), .B(
        Ciphertext_s2[34]), .Z(new_AGEMA_signal_1843) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_XX_2_), .B(SubCellInst_SboxInst_8_n3), .Z(
        SubCellInst_SboxInst_8_Q6) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1270), 
        .B(Ciphertext_s1[34]), .Z(new_AGEMA_signal_1844) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1271), 
        .B(Ciphertext_s2[34]), .Z(new_AGEMA_signal_1845) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_8_Q1), .B(SubCellInst_SboxInst_8_Q6), .ZN(
        SubCellInst_SboxInst_8_L1) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1840), 
        .B(new_AGEMA_signal_1844), .Z(new_AGEMA_signal_1984) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1841), 
        .B(new_AGEMA_signal_1845), .Z(new_AGEMA_signal_1985) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_n3), .Z(SubCellInst_SboxInst_8_L2) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        Ciphertext_s1[34]), .Z(new_AGEMA_signal_1846) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[33]), .B(
        Ciphertext_s2[34]), .Z(new_AGEMA_signal_1847) );
  INV_X1 SubCellInst_SboxInst_9_U1_U1 ( .A(Ciphertext_s0[38]), .ZN(
        SubCellInst_SboxInst_9_n3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[38]), 
        .B(Ciphertext_s0[39]), .Z(SubCellInst_SboxInst_9_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[38]), 
        .B(Ciphertext_s1[39]), .Z(new_AGEMA_signal_1278) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[38]), 
        .B(Ciphertext_s2[39]), .Z(new_AGEMA_signal_1279) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[36]), 
        .B(Ciphertext_s0[38]), .Z(SubCellInst_SboxInst_9_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[36]), 
        .B(Ciphertext_s1[38]), .Z(new_AGEMA_signal_1282) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[36]), 
        .B(Ciphertext_s2[38]), .Z(new_AGEMA_signal_1283) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_XX_2_), .Z(SubCellInst_SboxInst_9_Q0) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        new_AGEMA_signal_1282), .Z(new_AGEMA_signal_1850) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[37]), .B(
        new_AGEMA_signal_1283), .Z(new_AGEMA_signal_1851) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_XX_1_), .Z(SubCellInst_SboxInst_9_Q1) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        new_AGEMA_signal_1278), .Z(new_AGEMA_signal_1852) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[37]), .B(
        new_AGEMA_signal_1279), .Z(new_AGEMA_signal_1853) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_n3), .ZN(SubCellInst_SboxInst_9_Q4) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        Ciphertext_s1[38]), .Z(new_AGEMA_signal_1854) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[37]), .B(
        Ciphertext_s2[38]), .Z(new_AGEMA_signal_1855) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_XX_2_), .B(SubCellInst_SboxInst_9_n3), .Z(
        SubCellInst_SboxInst_9_Q6) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1282), 
        .B(Ciphertext_s1[38]), .Z(new_AGEMA_signal_1856) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1283), 
        .B(Ciphertext_s2[38]), .Z(new_AGEMA_signal_1857) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_9_Q1), .B(SubCellInst_SboxInst_9_Q6), .ZN(
        SubCellInst_SboxInst_9_L1) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1852), 
        .B(new_AGEMA_signal_1856), .Z(new_AGEMA_signal_1990) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1853), 
        .B(new_AGEMA_signal_1857), .Z(new_AGEMA_signal_1991) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_n3), .Z(SubCellInst_SboxInst_9_L2) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        Ciphertext_s1[38]), .Z(new_AGEMA_signal_1858) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[37]), .B(
        Ciphertext_s2[38]), .Z(new_AGEMA_signal_1859) );
  INV_X1 SubCellInst_SboxInst_10_U1_U1 ( .A(Ciphertext_s0[42]), .ZN(
        SubCellInst_SboxInst_10_n3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[42]), 
        .B(Ciphertext_s0[43]), .Z(SubCellInst_SboxInst_10_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[42]), 
        .B(Ciphertext_s1[43]), .Z(new_AGEMA_signal_1290) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[42]), 
        .B(Ciphertext_s2[43]), .Z(new_AGEMA_signal_1291) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[40]), 
        .B(Ciphertext_s0[42]), .Z(SubCellInst_SboxInst_10_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[40]), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1294) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[40]), 
        .B(Ciphertext_s2[42]), .Z(new_AGEMA_signal_1295) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_XX_2_), .Z(SubCellInst_SboxInst_10_Q0) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(new_AGEMA_signal_1294), .Z(new_AGEMA_signal_1862) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[41]), 
        .B(new_AGEMA_signal_1295), .Z(new_AGEMA_signal_1863) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_XX_1_), .Z(SubCellInst_SboxInst_10_Q1) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(new_AGEMA_signal_1290), .Z(new_AGEMA_signal_1864) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[41]), 
        .B(new_AGEMA_signal_1291), .Z(new_AGEMA_signal_1865) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_n3), .ZN(SubCellInst_SboxInst_10_Q4) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1866) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[41]), 
        .B(Ciphertext_s2[42]), .Z(new_AGEMA_signal_1867) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_XX_2_), .B(SubCellInst_SboxInst_10_n3), .Z(
        SubCellInst_SboxInst_10_Q6) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1294), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1868) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1295), 
        .B(Ciphertext_s2[42]), .Z(new_AGEMA_signal_1869) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_10_Q1), .B(SubCellInst_SboxInst_10_Q6), .ZN(
        SubCellInst_SboxInst_10_L1) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1864), 
        .B(new_AGEMA_signal_1868), .Z(new_AGEMA_signal_1996) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1865), 
        .B(new_AGEMA_signal_1869), .Z(new_AGEMA_signal_1997) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_n3), .Z(SubCellInst_SboxInst_10_L2) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1870) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[41]), 
        .B(Ciphertext_s2[42]), .Z(new_AGEMA_signal_1871) );
  INV_X1 SubCellInst_SboxInst_11_U1_U1 ( .A(Ciphertext_s0[46]), .ZN(
        SubCellInst_SboxInst_11_n3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[46]), 
        .B(Ciphertext_s0[47]), .Z(SubCellInst_SboxInst_11_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[46]), 
        .B(Ciphertext_s1[47]), .Z(new_AGEMA_signal_1302) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[46]), 
        .B(Ciphertext_s2[47]), .Z(new_AGEMA_signal_1303) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[44]), 
        .B(Ciphertext_s0[46]), .Z(SubCellInst_SboxInst_11_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[44]), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1306) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[44]), 
        .B(Ciphertext_s2[46]), .Z(new_AGEMA_signal_1307) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_XX_2_), .Z(SubCellInst_SboxInst_11_Q0) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(new_AGEMA_signal_1306), .Z(new_AGEMA_signal_1874) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[45]), 
        .B(new_AGEMA_signal_1307), .Z(new_AGEMA_signal_1875) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_XX_1_), .Z(SubCellInst_SboxInst_11_Q1) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(new_AGEMA_signal_1302), .Z(new_AGEMA_signal_1876) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[45]), 
        .B(new_AGEMA_signal_1303), .Z(new_AGEMA_signal_1877) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_n3), .ZN(SubCellInst_SboxInst_11_Q4) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1878) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[45]), 
        .B(Ciphertext_s2[46]), .Z(new_AGEMA_signal_1879) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_XX_2_), .B(SubCellInst_SboxInst_11_n3), .Z(
        SubCellInst_SboxInst_11_Q6) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1306), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1880) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1307), 
        .B(Ciphertext_s2[46]), .Z(new_AGEMA_signal_1881) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_11_Q1), .B(SubCellInst_SboxInst_11_Q6), .ZN(
        SubCellInst_SboxInst_11_L1) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1876), 
        .B(new_AGEMA_signal_1880), .Z(new_AGEMA_signal_2002) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1877), 
        .B(new_AGEMA_signal_1881), .Z(new_AGEMA_signal_2003) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_n3), .Z(SubCellInst_SboxInst_11_L2) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1882) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[45]), 
        .B(Ciphertext_s2[46]), .Z(new_AGEMA_signal_1883) );
  INV_X1 SubCellInst_SboxInst_12_U1_U1 ( .A(Ciphertext_s0[50]), .ZN(
        SubCellInst_SboxInst_12_n3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[50]), 
        .B(Ciphertext_s0[51]), .Z(SubCellInst_SboxInst_12_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[50]), 
        .B(Ciphertext_s1[51]), .Z(new_AGEMA_signal_1314) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[50]), 
        .B(Ciphertext_s2[51]), .Z(new_AGEMA_signal_1315) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[48]), 
        .B(Ciphertext_s0[50]), .Z(SubCellInst_SboxInst_12_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[48]), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1318) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[48]), 
        .B(Ciphertext_s2[50]), .Z(new_AGEMA_signal_1319) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_XX_2_), .Z(SubCellInst_SboxInst_12_Q0) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(new_AGEMA_signal_1318), .Z(new_AGEMA_signal_1886) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[49]), 
        .B(new_AGEMA_signal_1319), .Z(new_AGEMA_signal_1887) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_XX_1_), .Z(SubCellInst_SboxInst_12_Q1) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(new_AGEMA_signal_1314), .Z(new_AGEMA_signal_1888) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[49]), 
        .B(new_AGEMA_signal_1315), .Z(new_AGEMA_signal_1889) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_n3), .ZN(SubCellInst_SboxInst_12_Q4) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1890) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[49]), 
        .B(Ciphertext_s2[50]), .Z(new_AGEMA_signal_1891) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_XX_2_), .B(SubCellInst_SboxInst_12_n3), .Z(
        SubCellInst_SboxInst_12_Q6) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1318), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1892) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1319), 
        .B(Ciphertext_s2[50]), .Z(new_AGEMA_signal_1893) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_12_Q1), .B(SubCellInst_SboxInst_12_Q6), .ZN(
        SubCellInst_SboxInst_12_L1) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1888), 
        .B(new_AGEMA_signal_1892), .Z(new_AGEMA_signal_2008) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1889), 
        .B(new_AGEMA_signal_1893), .Z(new_AGEMA_signal_2009) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_n3), .Z(SubCellInst_SboxInst_12_L2) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1894) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[49]), 
        .B(Ciphertext_s2[50]), .Z(new_AGEMA_signal_1895) );
  INV_X1 SubCellInst_SboxInst_13_U1_U1 ( .A(Ciphertext_s0[54]), .ZN(
        SubCellInst_SboxInst_13_n3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[54]), 
        .B(Ciphertext_s0[55]), .Z(SubCellInst_SboxInst_13_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[54]), 
        .B(Ciphertext_s1[55]), .Z(new_AGEMA_signal_1326) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[54]), 
        .B(Ciphertext_s2[55]), .Z(new_AGEMA_signal_1327) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[52]), 
        .B(Ciphertext_s0[54]), .Z(SubCellInst_SboxInst_13_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[52]), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1330) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[52]), 
        .B(Ciphertext_s2[54]), .Z(new_AGEMA_signal_1331) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_XX_2_), .Z(SubCellInst_SboxInst_13_Q0) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(new_AGEMA_signal_1330), .Z(new_AGEMA_signal_1898) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[53]), 
        .B(new_AGEMA_signal_1331), .Z(new_AGEMA_signal_1899) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_XX_1_), .Z(SubCellInst_SboxInst_13_Q1) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(new_AGEMA_signal_1326), .Z(new_AGEMA_signal_1900) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[53]), 
        .B(new_AGEMA_signal_1327), .Z(new_AGEMA_signal_1901) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_n3), .ZN(SubCellInst_SboxInst_13_Q4) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1902) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[53]), 
        .B(Ciphertext_s2[54]), .Z(new_AGEMA_signal_1903) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_XX_2_), .B(SubCellInst_SboxInst_13_n3), .Z(
        SubCellInst_SboxInst_13_Q6) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1330), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1904) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1331), 
        .B(Ciphertext_s2[54]), .Z(new_AGEMA_signal_1905) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_13_Q1), .B(SubCellInst_SboxInst_13_Q6), .ZN(
        SubCellInst_SboxInst_13_L1) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1900), 
        .B(new_AGEMA_signal_1904), .Z(new_AGEMA_signal_2014) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1901), 
        .B(new_AGEMA_signal_1905), .Z(new_AGEMA_signal_2015) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_n3), .Z(SubCellInst_SboxInst_13_L2) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1906) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[53]), 
        .B(Ciphertext_s2[54]), .Z(new_AGEMA_signal_1907) );
  INV_X1 SubCellInst_SboxInst_14_U1_U1 ( .A(Ciphertext_s0[58]), .ZN(
        SubCellInst_SboxInst_14_n3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[58]), 
        .B(Ciphertext_s0[59]), .Z(SubCellInst_SboxInst_14_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[58]), 
        .B(Ciphertext_s1[59]), .Z(new_AGEMA_signal_1338) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[58]), 
        .B(Ciphertext_s2[59]), .Z(new_AGEMA_signal_1339) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[56]), 
        .B(Ciphertext_s0[58]), .Z(SubCellInst_SboxInst_14_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[56]), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1342) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[56]), 
        .B(Ciphertext_s2[58]), .Z(new_AGEMA_signal_1343) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_XX_2_), .Z(SubCellInst_SboxInst_14_Q0) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(new_AGEMA_signal_1342), .Z(new_AGEMA_signal_1910) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[57]), 
        .B(new_AGEMA_signal_1343), .Z(new_AGEMA_signal_1911) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_XX_1_), .Z(SubCellInst_SboxInst_14_Q1) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(new_AGEMA_signal_1338), .Z(new_AGEMA_signal_1912) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[57]), 
        .B(new_AGEMA_signal_1339), .Z(new_AGEMA_signal_1913) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_n3), .ZN(SubCellInst_SboxInst_14_Q4) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1914) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[57]), 
        .B(Ciphertext_s2[58]), .Z(new_AGEMA_signal_1915) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_XX_2_), .B(SubCellInst_SboxInst_14_n3), .Z(
        SubCellInst_SboxInst_14_Q6) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1342), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1916) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1343), 
        .B(Ciphertext_s2[58]), .Z(new_AGEMA_signal_1917) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_14_Q1), .B(SubCellInst_SboxInst_14_Q6), .ZN(
        SubCellInst_SboxInst_14_L1) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1912), 
        .B(new_AGEMA_signal_1916), .Z(new_AGEMA_signal_2020) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1913), 
        .B(new_AGEMA_signal_1917), .Z(new_AGEMA_signal_2021) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_n3), .Z(SubCellInst_SboxInst_14_L2) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1918) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[57]), 
        .B(Ciphertext_s2[58]), .Z(new_AGEMA_signal_1919) );
  INV_X1 SubCellInst_SboxInst_15_U1_U1 ( .A(Ciphertext_s0[62]), .ZN(
        SubCellInst_SboxInst_15_n3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[62]), 
        .B(Ciphertext_s0[63]), .Z(SubCellInst_SboxInst_15_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[62]), 
        .B(Ciphertext_s1[63]), .Z(new_AGEMA_signal_1350) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i1_U1_Ins_2_U1 ( .A(Ciphertext_s2[62]), 
        .B(Ciphertext_s2[63]), .Z(new_AGEMA_signal_1351) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[60]), 
        .B(Ciphertext_s0[62]), .Z(SubCellInst_SboxInst_15_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[60]), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1354) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i2_U1_Ins_2_U1 ( .A(Ciphertext_s2[60]), 
        .B(Ciphertext_s2[62]), .Z(new_AGEMA_signal_1355) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_XX_2_), .Z(SubCellInst_SboxInst_15_Q0) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(new_AGEMA_signal_1354), .Z(new_AGEMA_signal_1922) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR0_U1_Ins_2_U1 ( .A(Ciphertext_s2[61]), 
        .B(new_AGEMA_signal_1355), .Z(new_AGEMA_signal_1923) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_XX_1_), .Z(SubCellInst_SboxInst_15_Q1) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(new_AGEMA_signal_1350), .Z(new_AGEMA_signal_1924) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR1_U1_Ins_2_U1 ( .A(Ciphertext_s2[61]), 
        .B(new_AGEMA_signal_1351), .Z(new_AGEMA_signal_1925) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_n3), .ZN(SubCellInst_SboxInst_15_Q4) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1926) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR3_U1_Ins_2_U1 ( .A(Ciphertext_s2[61]), 
        .B(Ciphertext_s2[62]), .Z(new_AGEMA_signal_1927) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_XX_2_), .B(SubCellInst_SboxInst_15_n3), .Z(
        SubCellInst_SboxInst_15_Q6) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1354), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1928) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1355), 
        .B(Ciphertext_s2[62]), .Z(new_AGEMA_signal_1929) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_15_Q1), .B(SubCellInst_SboxInst_15_Q6), .ZN(
        SubCellInst_SboxInst_15_L1) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1924), 
        .B(new_AGEMA_signal_1928), .Z(new_AGEMA_signal_2026) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_1925), 
        .B(new_AGEMA_signal_1929), .Z(new_AGEMA_signal_2027) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_n3), .Z(SubCellInst_SboxInst_15_L2) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1930) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR8_U1_Ins_2_U1 ( .A(Ciphertext_s2[61]), 
        .B(Ciphertext_s2[62]), .Z(new_AGEMA_signal_1931) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_0_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[0]), .B(Key_s0[0]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[0]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_0_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1356), .B(Key_s1[0]), .S(rst), .Z(
        new_AGEMA_signal_1360) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_0_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1357), .B(Key_s2[0]), .S(rst), .Z(
        new_AGEMA_signal_1361) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_1_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[1]), .B(Key_s0[1]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[1]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1362), .B(Key_s1[1]), .S(rst), .Z(
        new_AGEMA_signal_1366) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1363), .B(Key_s2[1]), .S(rst), .Z(
        new_AGEMA_signal_1367) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_2_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[2]), .B(Key_s0[2]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[2]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_2_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1368), .B(Key_s1[2]), .S(rst), .Z(
        new_AGEMA_signal_1372) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_2_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1369), .B(Key_s2[2]), .S(rst), .Z(
        new_AGEMA_signal_1373) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_3_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[3]), .B(Key_s0[3]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[3]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_3_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1374), .B(Key_s1[3]), .S(rst), .Z(
        new_AGEMA_signal_1378) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_3_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1375), .B(Key_s2[3]), .S(rst), .Z(
        new_AGEMA_signal_1379) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_4_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[4]), .B(Key_s0[4]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[4]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_4_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1380), .B(Key_s1[4]), .S(rst), .Z(
        new_AGEMA_signal_1384) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_4_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1381), .B(Key_s2[4]), .S(rst), .Z(
        new_AGEMA_signal_1385) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_5_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[5]), .B(Key_s0[5]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[5]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_5_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1386), .B(Key_s1[5]), .S(rst), .Z(
        new_AGEMA_signal_1390) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_5_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1387), .B(Key_s2[5]), .S(rst), .Z(
        new_AGEMA_signal_1391) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_6_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[6]), .B(Key_s0[6]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[6]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_6_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1392), .B(Key_s1[6]), .S(rst), .Z(
        new_AGEMA_signal_1396) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_6_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1393), .B(Key_s2[6]), .S(rst), .Z(
        new_AGEMA_signal_1397) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_7_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[7]), .B(Key_s0[7]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[7]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_7_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1398), .B(Key_s1[7]), .S(rst), .Z(
        new_AGEMA_signal_1402) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_7_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1399), .B(Key_s2[7]), .S(rst), .Z(
        new_AGEMA_signal_1403) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_8_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[8]), .B(Key_s0[8]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[8]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_8_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1404), .B(Key_s1[8]), .S(rst), .Z(
        new_AGEMA_signal_1408) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_8_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1405), .B(Key_s2[8]), .S(rst), .Z(
        new_AGEMA_signal_1409) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_9_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[9]), .B(Key_s0[9]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[9]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_9_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1410), .B(Key_s1[9]), .S(rst), .Z(
        new_AGEMA_signal_1414) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_9_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1411), .B(Key_s2[9]), .S(rst), .Z(
        new_AGEMA_signal_1415) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_10_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[10]), .B(Key_s0[10]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[10]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_10_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1416), .B(Key_s1[10]), .S(rst), .Z(
        new_AGEMA_signal_1420) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_10_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1417), .B(Key_s2[10]), .S(rst), .Z(
        new_AGEMA_signal_1421) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_11_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[11]), .B(Key_s0[11]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[11]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_11_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1422), .B(Key_s1[11]), .S(rst), .Z(
        new_AGEMA_signal_1426) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_11_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1423), .B(Key_s2[11]), .S(rst), .Z(
        new_AGEMA_signal_1427) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_12_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[12]), .B(Key_s0[12]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[12]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_12_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1428), .B(Key_s1[12]), .S(rst), .Z(
        new_AGEMA_signal_1432) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_12_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1429), .B(Key_s2[12]), .S(rst), .Z(
        new_AGEMA_signal_1433) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_13_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[13]), .B(Key_s0[13]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[13]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_13_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1434), .B(Key_s1[13]), .S(rst), .Z(
        new_AGEMA_signal_1438) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_13_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1435), .B(Key_s2[13]), .S(rst), .Z(
        new_AGEMA_signal_1439) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_14_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[14]), .B(Key_s0[14]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[14]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_14_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1440), .B(Key_s1[14]), .S(rst), .Z(
        new_AGEMA_signal_1444) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_14_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1441), .B(Key_s2[14]), .S(rst), .Z(
        new_AGEMA_signal_1445) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_15_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[15]), .B(Key_s0[15]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[15]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_15_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1446), .B(Key_s1[15]), .S(rst), .Z(
        new_AGEMA_signal_1450) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_15_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1447), .B(Key_s2[15]), .S(rst), .Z(
        new_AGEMA_signal_1451) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_16_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[16]), .B(Key_s0[16]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[16]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_16_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1452), .B(Key_s1[16]), .S(rst), .Z(
        new_AGEMA_signal_1456) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_16_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1453), .B(Key_s2[16]), .S(rst), .Z(
        new_AGEMA_signal_1457) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_17_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[17]), .B(Key_s0[17]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[17]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_17_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1458), .B(Key_s1[17]), .S(rst), .Z(
        new_AGEMA_signal_1462) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_17_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1459), .B(Key_s2[17]), .S(rst), .Z(
        new_AGEMA_signal_1463) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_18_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[18]), .B(Key_s0[18]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[18]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_18_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1464), .B(Key_s1[18]), .S(rst), .Z(
        new_AGEMA_signal_1468) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_18_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1465), .B(Key_s2[18]), .S(rst), .Z(
        new_AGEMA_signal_1469) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_19_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[19]), .B(Key_s0[19]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[19]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_19_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1470), .B(Key_s1[19]), .S(rst), .Z(
        new_AGEMA_signal_1474) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_19_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1471), .B(Key_s2[19]), .S(rst), .Z(
        new_AGEMA_signal_1475) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_20_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[20]), .B(Key_s0[20]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[20]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_20_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1476), .B(Key_s1[20]), .S(rst), .Z(
        new_AGEMA_signal_1480) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_20_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1477), .B(Key_s2[20]), .S(rst), .Z(
        new_AGEMA_signal_1481) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_21_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[21]), .B(Key_s0[21]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[21]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_21_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1482), .B(Key_s1[21]), .S(rst), .Z(
        new_AGEMA_signal_1486) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_21_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1483), .B(Key_s2[21]), .S(rst), .Z(
        new_AGEMA_signal_1487) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_22_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[22]), .B(Key_s0[22]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[22]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_22_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1488), .B(Key_s1[22]), .S(rst), .Z(
        new_AGEMA_signal_1492) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_22_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1489), .B(Key_s2[22]), .S(rst), .Z(
        new_AGEMA_signal_1493) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_23_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[23]), .B(Key_s0[23]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[23]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_23_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1494), .B(Key_s1[23]), .S(rst), .Z(
        new_AGEMA_signal_1498) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_23_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1495), .B(Key_s2[23]), .S(rst), .Z(
        new_AGEMA_signal_1499) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_24_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[24]), .B(Key_s0[24]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[24]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_24_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1500), .B(Key_s1[24]), .S(rst), .Z(
        new_AGEMA_signal_1504) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_24_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1501), .B(Key_s2[24]), .S(rst), .Z(
        new_AGEMA_signal_1505) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_25_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[25]), .B(Key_s0[25]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[25]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_25_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1506), .B(Key_s1[25]), .S(rst), .Z(
        new_AGEMA_signal_1510) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_25_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1507), .B(Key_s2[25]), .S(rst), .Z(
        new_AGEMA_signal_1511) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_26_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[26]), .B(Key_s0[26]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[26]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_26_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1512), .B(Key_s1[26]), .S(rst), .Z(
        new_AGEMA_signal_1516) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_26_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1513), .B(Key_s2[26]), .S(rst), .Z(
        new_AGEMA_signal_1517) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_27_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[27]), .B(Key_s0[27]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[27]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_27_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1518), .B(Key_s1[27]), .S(rst), .Z(
        new_AGEMA_signal_1522) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_27_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1519), .B(Key_s2[27]), .S(rst), .Z(
        new_AGEMA_signal_1523) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_28_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[28]), .B(Key_s0[28]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[28]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_28_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1524), .B(Key_s1[28]), .S(rst), .Z(
        new_AGEMA_signal_1528) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_28_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1525), .B(Key_s2[28]), .S(rst), .Z(
        new_AGEMA_signal_1529) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_29_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[29]), .B(Key_s0[29]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[29]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_29_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1530), .B(Key_s1[29]), .S(rst), .Z(
        new_AGEMA_signal_1534) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_29_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1531), .B(Key_s2[29]), .S(rst), .Z(
        new_AGEMA_signal_1535) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_30_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[30]), .B(Key_s0[30]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[30]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_30_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1536), .B(Key_s1[30]), .S(rst), .Z(
        new_AGEMA_signal_1540) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_30_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1537), .B(Key_s2[30]), .S(rst), .Z(
        new_AGEMA_signal_1541) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_31_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[31]), .B(Key_s0[31]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[31]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_31_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1542), .B(Key_s1[31]), .S(rst), .Z(
        new_AGEMA_signal_1546) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_31_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1543), .B(Key_s2[31]), .S(rst), .Z(
        new_AGEMA_signal_1547) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_32_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[32]), .B(Key_s0[32]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[32]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_32_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1548), .B(Key_s1[32]), .S(rst), .Z(
        new_AGEMA_signal_1552) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_32_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1549), .B(Key_s2[32]), .S(rst), .Z(
        new_AGEMA_signal_1553) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_33_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[33]), .B(Key_s0[33]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[33]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_33_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1554), .B(Key_s1[33]), .S(rst), .Z(
        new_AGEMA_signal_1558) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_33_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1555), .B(Key_s2[33]), .S(rst), .Z(
        new_AGEMA_signal_1559) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_34_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[34]), .B(Key_s0[34]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[34]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_34_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1560), .B(Key_s1[34]), .S(rst), .Z(
        new_AGEMA_signal_1564) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_34_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1561), .B(Key_s2[34]), .S(rst), .Z(
        new_AGEMA_signal_1565) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_35_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[35]), .B(Key_s0[35]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[35]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_35_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1566), .B(Key_s1[35]), .S(rst), .Z(
        new_AGEMA_signal_1570) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_35_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1567), .B(Key_s2[35]), .S(rst), .Z(
        new_AGEMA_signal_1571) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_36_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[36]), .B(Key_s0[36]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[36]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_36_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1572), .B(Key_s1[36]), .S(rst), .Z(
        new_AGEMA_signal_1576) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_36_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1573), .B(Key_s2[36]), .S(rst), .Z(
        new_AGEMA_signal_1577) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_37_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[37]), .B(Key_s0[37]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[37]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_37_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1578), .B(Key_s1[37]), .S(rst), .Z(
        new_AGEMA_signal_1582) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_37_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1579), .B(Key_s2[37]), .S(rst), .Z(
        new_AGEMA_signal_1583) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_38_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[38]), .B(Key_s0[38]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[38]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_38_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1584), .B(Key_s1[38]), .S(rst), .Z(
        new_AGEMA_signal_1588) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_38_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1585), .B(Key_s2[38]), .S(rst), .Z(
        new_AGEMA_signal_1589) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_39_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[39]), .B(Key_s0[39]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[39]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_39_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1590), .B(Key_s1[39]), .S(rst), .Z(
        new_AGEMA_signal_1594) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_39_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1591), .B(Key_s2[39]), .S(rst), .Z(
        new_AGEMA_signal_1595) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_40_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[40]), .B(Key_s0[40]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[40]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_40_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1596), .B(Key_s1[40]), .S(rst), .Z(
        new_AGEMA_signal_1600) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_40_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1597), .B(Key_s2[40]), .S(rst), .Z(
        new_AGEMA_signal_1601) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_41_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[41]), .B(Key_s0[41]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[41]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_41_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1602), .B(Key_s1[41]), .S(rst), .Z(
        new_AGEMA_signal_1606) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_41_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1603), .B(Key_s2[41]), .S(rst), .Z(
        new_AGEMA_signal_1607) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_42_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[42]), .B(Key_s0[42]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[42]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_42_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1608), .B(Key_s1[42]), .S(rst), .Z(
        new_AGEMA_signal_1612) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_42_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1609), .B(Key_s2[42]), .S(rst), .Z(
        new_AGEMA_signal_1613) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_43_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[43]), .B(Key_s0[43]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[43]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_43_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1614), .B(Key_s1[43]), .S(rst), .Z(
        new_AGEMA_signal_1618) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_43_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1615), .B(Key_s2[43]), .S(rst), .Z(
        new_AGEMA_signal_1619) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_44_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[44]), .B(Key_s0[44]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[44]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_44_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1620), .B(Key_s1[44]), .S(rst), .Z(
        new_AGEMA_signal_1624) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_44_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1621), .B(Key_s2[44]), .S(rst), .Z(
        new_AGEMA_signal_1625) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_45_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[45]), .B(Key_s0[45]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[45]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_45_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1626), .B(Key_s1[45]), .S(rst), .Z(
        new_AGEMA_signal_1630) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_45_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1627), .B(Key_s2[45]), .S(rst), .Z(
        new_AGEMA_signal_1631) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_46_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[46]), .B(Key_s0[46]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[46]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_46_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1632), .B(Key_s1[46]), .S(rst), .Z(
        new_AGEMA_signal_1636) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_46_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1633), .B(Key_s2[46]), .S(rst), .Z(
        new_AGEMA_signal_1637) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_47_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[47]), .B(Key_s0[47]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[47]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_47_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1638), .B(Key_s1[47]), .S(rst), .Z(
        new_AGEMA_signal_1642) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_47_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1639), .B(Key_s2[47]), .S(rst), .Z(
        new_AGEMA_signal_1643) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_48_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[48]), .B(Key_s0[48]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[48]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_48_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1644), .B(Key_s1[48]), .S(rst), .Z(
        new_AGEMA_signal_1648) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_48_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1645), .B(Key_s2[48]), .S(rst), .Z(
        new_AGEMA_signal_1649) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_49_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[49]), .B(Key_s0[49]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[49]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_49_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1650), .B(Key_s1[49]), .S(rst), .Z(
        new_AGEMA_signal_1654) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_49_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1651), .B(Key_s2[49]), .S(rst), .Z(
        new_AGEMA_signal_1655) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_50_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[50]), .B(Key_s0[50]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[50]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_50_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1656), .B(Key_s1[50]), .S(rst), .Z(
        new_AGEMA_signal_1660) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_50_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1657), .B(Key_s2[50]), .S(rst), .Z(
        new_AGEMA_signal_1661) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_51_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[51]), .B(Key_s0[51]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[51]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_51_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1662), .B(Key_s1[51]), .S(rst), .Z(
        new_AGEMA_signal_1666) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_51_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1663), .B(Key_s2[51]), .S(rst), .Z(
        new_AGEMA_signal_1667) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_52_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[52]), .B(Key_s0[52]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[52]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_52_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1668), .B(Key_s1[52]), .S(rst), .Z(
        new_AGEMA_signal_1672) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_52_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1669), .B(Key_s2[52]), .S(rst), .Z(
        new_AGEMA_signal_1673) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_53_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[53]), .B(Key_s0[53]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[53]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_53_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1674), .B(Key_s1[53]), .S(rst), .Z(
        new_AGEMA_signal_1678) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_53_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1675), .B(Key_s2[53]), .S(rst), .Z(
        new_AGEMA_signal_1679) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_54_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[54]), .B(Key_s0[54]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[54]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_54_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1680), .B(Key_s1[54]), .S(rst), .Z(
        new_AGEMA_signal_1684) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_54_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1681), .B(Key_s2[54]), .S(rst), .Z(
        new_AGEMA_signal_1685) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_55_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[55]), .B(Key_s0[55]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[55]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_55_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1686), .B(Key_s1[55]), .S(rst), .Z(
        new_AGEMA_signal_1690) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_55_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1687), .B(Key_s2[55]), .S(rst), .Z(
        new_AGEMA_signal_1691) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_56_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[56]), .B(Key_s0[56]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[56]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_56_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1692), .B(Key_s1[56]), .S(rst), .Z(
        new_AGEMA_signal_1696) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_56_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1693), .B(Key_s2[56]), .S(rst), .Z(
        new_AGEMA_signal_1697) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_57_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[57]), .B(Key_s0[57]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[57]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_57_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1698), .B(Key_s1[57]), .S(rst), .Z(
        new_AGEMA_signal_1702) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_57_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1699), .B(Key_s2[57]), .S(rst), .Z(
        new_AGEMA_signal_1703) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_58_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[58]), .B(Key_s0[58]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[58]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_58_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1704), .B(Key_s1[58]), .S(rst), .Z(
        new_AGEMA_signal_1708) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_58_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1705), .B(Key_s2[58]), .S(rst), .Z(
        new_AGEMA_signal_1709) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_59_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[59]), .B(Key_s0[59]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[59]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_59_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1710), .B(Key_s1[59]), .S(rst), .Z(
        new_AGEMA_signal_1714) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_59_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1711), .B(Key_s2[59]), .S(rst), .Z(
        new_AGEMA_signal_1715) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_60_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[60]), .B(Key_s0[60]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[60]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_60_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1716), .B(Key_s1[60]), .S(rst), .Z(
        new_AGEMA_signal_1720) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_60_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1717), .B(Key_s2[60]), .S(rst), .Z(
        new_AGEMA_signal_1721) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_61_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[61]), .B(Key_s0[61]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[61]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_61_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1722), .B(Key_s1[61]), .S(rst), .Z(
        new_AGEMA_signal_1726) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_61_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1723), .B(Key_s2[61]), .S(rst), .Z(
        new_AGEMA_signal_1727) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_62_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[62]), .B(Key_s0[62]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[62]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_62_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1728), .B(Key_s1[62]), .S(rst), .Z(
        new_AGEMA_signal_1732) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_62_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1729), .B(Key_s2[62]), .S(rst), .Z(
        new_AGEMA_signal_1733) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_63_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[63]), .B(Key_s0[63]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[63]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_63_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1734), .B(Key_s1[63]), .S(rst), .Z(
        new_AGEMA_signal_1738) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_63_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_1735), .B(Key_s2[63]), .S(rst), .Z(
        new_AGEMA_signal_1739) );
  DFF_X1 new_AGEMA_reg_buffer_1000_s_current_state_reg ( .D(rst), .CK(clk), 
        .Q(new_AGEMA_signal_3278), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1002_s_current_state_reg ( .D(Plaintext_s0[2]), 
        .CK(clk), .Q(new_AGEMA_signal_3280), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1004_s_current_state_reg ( .D(Plaintext_s1[2]), 
        .CK(clk), .Q(new_AGEMA_signal_3282), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1006_s_current_state_reg ( .D(Plaintext_s2[2]), 
        .CK(clk), .Q(new_AGEMA_signal_3284), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1008_s_current_state_reg ( .D(Plaintext_s0[3]), 
        .CK(clk), .Q(new_AGEMA_signal_3286), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1010_s_current_state_reg ( .D(Plaintext_s1[3]), 
        .CK(clk), .Q(new_AGEMA_signal_3288), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1012_s_current_state_reg ( .D(Plaintext_s2[3]), 
        .CK(clk), .Q(new_AGEMA_signal_3290), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1014_s_current_state_reg ( .D(Plaintext_s0[6]), 
        .CK(clk), .Q(new_AGEMA_signal_3292), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1016_s_current_state_reg ( .D(Plaintext_s1[6]), 
        .CK(clk), .Q(new_AGEMA_signal_3294), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1018_s_current_state_reg ( .D(Plaintext_s2[6]), 
        .CK(clk), .Q(new_AGEMA_signal_3296), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1020_s_current_state_reg ( .D(Plaintext_s0[7]), 
        .CK(clk), .Q(new_AGEMA_signal_3298), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1022_s_current_state_reg ( .D(Plaintext_s1[7]), 
        .CK(clk), .Q(new_AGEMA_signal_3300), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1024_s_current_state_reg ( .D(Plaintext_s2[7]), 
        .CK(clk), .Q(new_AGEMA_signal_3302), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1026_s_current_state_reg ( .D(Plaintext_s0[10]), 
        .CK(clk), .Q(new_AGEMA_signal_3304), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1028_s_current_state_reg ( .D(Plaintext_s1[10]), 
        .CK(clk), .Q(new_AGEMA_signal_3306), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1030_s_current_state_reg ( .D(Plaintext_s2[10]), 
        .CK(clk), .Q(new_AGEMA_signal_3308), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1032_s_current_state_reg ( .D(Plaintext_s0[11]), 
        .CK(clk), .Q(new_AGEMA_signal_3310), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1034_s_current_state_reg ( .D(Plaintext_s1[11]), 
        .CK(clk), .Q(new_AGEMA_signal_3312), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1036_s_current_state_reg ( .D(Plaintext_s2[11]), 
        .CK(clk), .Q(new_AGEMA_signal_3314), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1038_s_current_state_reg ( .D(Plaintext_s0[14]), 
        .CK(clk), .Q(new_AGEMA_signal_3316), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1040_s_current_state_reg ( .D(Plaintext_s1[14]), 
        .CK(clk), .Q(new_AGEMA_signal_3318), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1042_s_current_state_reg ( .D(Plaintext_s2[14]), 
        .CK(clk), .Q(new_AGEMA_signal_3320), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1044_s_current_state_reg ( .D(Plaintext_s0[15]), 
        .CK(clk), .Q(new_AGEMA_signal_3322), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1046_s_current_state_reg ( .D(Plaintext_s1[15]), 
        .CK(clk), .Q(new_AGEMA_signal_3324), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1048_s_current_state_reg ( .D(Plaintext_s2[15]), 
        .CK(clk), .Q(new_AGEMA_signal_3326), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1050_s_current_state_reg ( .D(Plaintext_s0[18]), 
        .CK(clk), .Q(new_AGEMA_signal_3328), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1052_s_current_state_reg ( .D(Plaintext_s1[18]), 
        .CK(clk), .Q(new_AGEMA_signal_3330), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1054_s_current_state_reg ( .D(Plaintext_s2[18]), 
        .CK(clk), .Q(new_AGEMA_signal_3332), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1056_s_current_state_reg ( .D(Plaintext_s0[19]), 
        .CK(clk), .Q(new_AGEMA_signal_3334), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1058_s_current_state_reg ( .D(Plaintext_s1[19]), 
        .CK(clk), .Q(new_AGEMA_signal_3336), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1060_s_current_state_reg ( .D(Plaintext_s2[19]), 
        .CK(clk), .Q(new_AGEMA_signal_3338), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1062_s_current_state_reg ( .D(Plaintext_s0[22]), 
        .CK(clk), .Q(new_AGEMA_signal_3340), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1064_s_current_state_reg ( .D(Plaintext_s1[22]), 
        .CK(clk), .Q(new_AGEMA_signal_3342), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1066_s_current_state_reg ( .D(Plaintext_s2[22]), 
        .CK(clk), .Q(new_AGEMA_signal_3344), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1068_s_current_state_reg ( .D(Plaintext_s0[23]), 
        .CK(clk), .Q(new_AGEMA_signal_3346), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1070_s_current_state_reg ( .D(Plaintext_s1[23]), 
        .CK(clk), .Q(new_AGEMA_signal_3348), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1072_s_current_state_reg ( .D(Plaintext_s2[23]), 
        .CK(clk), .Q(new_AGEMA_signal_3350), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1074_s_current_state_reg ( .D(Plaintext_s0[26]), 
        .CK(clk), .Q(new_AGEMA_signal_3352), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1076_s_current_state_reg ( .D(Plaintext_s1[26]), 
        .CK(clk), .Q(new_AGEMA_signal_3354), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1078_s_current_state_reg ( .D(Plaintext_s2[26]), 
        .CK(clk), .Q(new_AGEMA_signal_3356), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1080_s_current_state_reg ( .D(Plaintext_s0[27]), 
        .CK(clk), .Q(new_AGEMA_signal_3358), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1082_s_current_state_reg ( .D(Plaintext_s1[27]), 
        .CK(clk), .Q(new_AGEMA_signal_3360), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1084_s_current_state_reg ( .D(Plaintext_s2[27]), 
        .CK(clk), .Q(new_AGEMA_signal_3362), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1086_s_current_state_reg ( .D(Plaintext_s0[30]), 
        .CK(clk), .Q(new_AGEMA_signal_3364), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1088_s_current_state_reg ( .D(Plaintext_s1[30]), 
        .CK(clk), .Q(new_AGEMA_signal_3366), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1090_s_current_state_reg ( .D(Plaintext_s2[30]), 
        .CK(clk), .Q(new_AGEMA_signal_3368), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1092_s_current_state_reg ( .D(Plaintext_s0[31]), 
        .CK(clk), .Q(new_AGEMA_signal_3370), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1094_s_current_state_reg ( .D(Plaintext_s1[31]), 
        .CK(clk), .Q(new_AGEMA_signal_3372), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1096_s_current_state_reg ( .D(Plaintext_s2[31]), 
        .CK(clk), .Q(new_AGEMA_signal_3374), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1098_s_current_state_reg ( .D(Plaintext_s0[34]), 
        .CK(clk), .Q(new_AGEMA_signal_3376), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1100_s_current_state_reg ( .D(Plaintext_s1[34]), 
        .CK(clk), .Q(new_AGEMA_signal_3378), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1102_s_current_state_reg ( .D(Plaintext_s2[34]), 
        .CK(clk), .Q(new_AGEMA_signal_3380), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1104_s_current_state_reg ( .D(Plaintext_s0[35]), 
        .CK(clk), .Q(new_AGEMA_signal_3382), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1106_s_current_state_reg ( .D(Plaintext_s1[35]), 
        .CK(clk), .Q(new_AGEMA_signal_3384), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1108_s_current_state_reg ( .D(Plaintext_s2[35]), 
        .CK(clk), .Q(new_AGEMA_signal_3386), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1110_s_current_state_reg ( .D(Plaintext_s0[38]), 
        .CK(clk), .Q(new_AGEMA_signal_3388), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1112_s_current_state_reg ( .D(Plaintext_s1[38]), 
        .CK(clk), .Q(new_AGEMA_signal_3390), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1114_s_current_state_reg ( .D(Plaintext_s2[38]), 
        .CK(clk), .Q(new_AGEMA_signal_3392), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1116_s_current_state_reg ( .D(Plaintext_s0[39]), 
        .CK(clk), .Q(new_AGEMA_signal_3394), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1118_s_current_state_reg ( .D(Plaintext_s1[39]), 
        .CK(clk), .Q(new_AGEMA_signal_3396), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1120_s_current_state_reg ( .D(Plaintext_s2[39]), 
        .CK(clk), .Q(new_AGEMA_signal_3398), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1122_s_current_state_reg ( .D(Plaintext_s0[42]), 
        .CK(clk), .Q(new_AGEMA_signal_3400), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1124_s_current_state_reg ( .D(Plaintext_s1[42]), 
        .CK(clk), .Q(new_AGEMA_signal_3402), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1126_s_current_state_reg ( .D(Plaintext_s2[42]), 
        .CK(clk), .Q(new_AGEMA_signal_3404), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1128_s_current_state_reg ( .D(Plaintext_s0[43]), 
        .CK(clk), .Q(new_AGEMA_signal_3406), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1130_s_current_state_reg ( .D(Plaintext_s1[43]), 
        .CK(clk), .Q(new_AGEMA_signal_3408), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1132_s_current_state_reg ( .D(Plaintext_s2[43]), 
        .CK(clk), .Q(new_AGEMA_signal_3410), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1134_s_current_state_reg ( .D(Plaintext_s0[46]), 
        .CK(clk), .Q(new_AGEMA_signal_3412), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1136_s_current_state_reg ( .D(Plaintext_s1[46]), 
        .CK(clk), .Q(new_AGEMA_signal_3414), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1138_s_current_state_reg ( .D(Plaintext_s2[46]), 
        .CK(clk), .Q(new_AGEMA_signal_3416), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1140_s_current_state_reg ( .D(Plaintext_s0[47]), 
        .CK(clk), .Q(new_AGEMA_signal_3418), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1142_s_current_state_reg ( .D(Plaintext_s1[47]), 
        .CK(clk), .Q(new_AGEMA_signal_3420), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1144_s_current_state_reg ( .D(Plaintext_s2[47]), 
        .CK(clk), .Q(new_AGEMA_signal_3422), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1146_s_current_state_reg ( .D(Plaintext_s0[50]), 
        .CK(clk), .Q(new_AGEMA_signal_3424), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1148_s_current_state_reg ( .D(Plaintext_s1[50]), 
        .CK(clk), .Q(new_AGEMA_signal_3426), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1150_s_current_state_reg ( .D(Plaintext_s2[50]), 
        .CK(clk), .Q(new_AGEMA_signal_3428), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1152_s_current_state_reg ( .D(Plaintext_s0[51]), 
        .CK(clk), .Q(new_AGEMA_signal_3430), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1154_s_current_state_reg ( .D(Plaintext_s1[51]), 
        .CK(clk), .Q(new_AGEMA_signal_3432), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1156_s_current_state_reg ( .D(Plaintext_s2[51]), 
        .CK(clk), .Q(new_AGEMA_signal_3434), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1158_s_current_state_reg ( .D(Plaintext_s0[54]), 
        .CK(clk), .Q(new_AGEMA_signal_3436), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1160_s_current_state_reg ( .D(Plaintext_s1[54]), 
        .CK(clk), .Q(new_AGEMA_signal_3438), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1162_s_current_state_reg ( .D(Plaintext_s2[54]), 
        .CK(clk), .Q(new_AGEMA_signal_3440), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1164_s_current_state_reg ( .D(Plaintext_s0[55]), 
        .CK(clk), .Q(new_AGEMA_signal_3442), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1166_s_current_state_reg ( .D(Plaintext_s1[55]), 
        .CK(clk), .Q(new_AGEMA_signal_3444), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1168_s_current_state_reg ( .D(Plaintext_s2[55]), 
        .CK(clk), .Q(new_AGEMA_signal_3446), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1170_s_current_state_reg ( .D(Plaintext_s0[58]), 
        .CK(clk), .Q(new_AGEMA_signal_3448), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1172_s_current_state_reg ( .D(Plaintext_s1[58]), 
        .CK(clk), .Q(new_AGEMA_signal_3450), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1174_s_current_state_reg ( .D(Plaintext_s2[58]), 
        .CK(clk), .Q(new_AGEMA_signal_3452), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1176_s_current_state_reg ( .D(Plaintext_s0[59]), 
        .CK(clk), .Q(new_AGEMA_signal_3454), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1178_s_current_state_reg ( .D(Plaintext_s1[59]), 
        .CK(clk), .Q(new_AGEMA_signal_3456), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1180_s_current_state_reg ( .D(Plaintext_s2[59]), 
        .CK(clk), .Q(new_AGEMA_signal_3458), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1182_s_current_state_reg ( .D(Plaintext_s0[62]), 
        .CK(clk), .Q(new_AGEMA_signal_3460), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1184_s_current_state_reg ( .D(Plaintext_s1[62]), 
        .CK(clk), .Q(new_AGEMA_signal_3462), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1186_s_current_state_reg ( .D(Plaintext_s2[62]), 
        .CK(clk), .Q(new_AGEMA_signal_3464), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1188_s_current_state_reg ( .D(Plaintext_s0[63]), 
        .CK(clk), .Q(new_AGEMA_signal_3466), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1190_s_current_state_reg ( .D(Plaintext_s1[63]), 
        .CK(clk), .Q(new_AGEMA_signal_3468), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1192_s_current_state_reg ( .D(Plaintext_s2[63]), 
        .CK(clk), .Q(new_AGEMA_signal_3470), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1194_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_Q0), .CK(clk), .Q(new_AGEMA_signal_3472), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1196_s_current_state_reg ( .D(
        new_AGEMA_signal_1742), .CK(clk), .Q(new_AGEMA_signal_3474), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1198_s_current_state_reg ( .D(
        new_AGEMA_signal_1743), .CK(clk), .Q(new_AGEMA_signal_3476), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1200_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_L1), .CK(clk), .Q(new_AGEMA_signal_3478), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1202_s_current_state_reg ( .D(
        new_AGEMA_signal_1936), .CK(clk), .Q(new_AGEMA_signal_3480), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1204_s_current_state_reg ( .D(
        new_AGEMA_signal_1937), .CK(clk), .Q(new_AGEMA_signal_3482), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1206_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_XX_2_), .CK(clk), .Q(new_AGEMA_signal_3484), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1208_s_current_state_reg ( .D(
        new_AGEMA_signal_1174), .CK(clk), .Q(new_AGEMA_signal_3486), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1210_s_current_state_reg ( .D(
        new_AGEMA_signal_1175), .CK(clk), .Q(new_AGEMA_signal_3488), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1212_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_XX_1_), .CK(clk), .Q(new_AGEMA_signal_3490), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1214_s_current_state_reg ( .D(
        new_AGEMA_signal_1170), .CK(clk), .Q(new_AGEMA_signal_3492), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1216_s_current_state_reg ( .D(
        new_AGEMA_signal_1171), .CK(clk), .Q(new_AGEMA_signal_3494), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1218_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_Q0), .CK(clk), .Q(new_AGEMA_signal_3496), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1220_s_current_state_reg ( .D(
        new_AGEMA_signal_1754), .CK(clk), .Q(new_AGEMA_signal_3498), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1222_s_current_state_reg ( .D(
        new_AGEMA_signal_1755), .CK(clk), .Q(new_AGEMA_signal_3500), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1224_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_L1), .CK(clk), .Q(new_AGEMA_signal_3502), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1226_s_current_state_reg ( .D(
        new_AGEMA_signal_1942), .CK(clk), .Q(new_AGEMA_signal_3504), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1228_s_current_state_reg ( .D(
        new_AGEMA_signal_1943), .CK(clk), .Q(new_AGEMA_signal_3506), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1230_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_XX_2_), .CK(clk), .Q(new_AGEMA_signal_3508), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1232_s_current_state_reg ( .D(
        new_AGEMA_signal_1186), .CK(clk), .Q(new_AGEMA_signal_3510), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1234_s_current_state_reg ( .D(
        new_AGEMA_signal_1187), .CK(clk), .Q(new_AGEMA_signal_3512), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1236_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_XX_1_), .CK(clk), .Q(new_AGEMA_signal_3514), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1238_s_current_state_reg ( .D(
        new_AGEMA_signal_1182), .CK(clk), .Q(new_AGEMA_signal_3516), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1240_s_current_state_reg ( .D(
        new_AGEMA_signal_1183), .CK(clk), .Q(new_AGEMA_signal_3518), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1242_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_Q0), .CK(clk), .Q(new_AGEMA_signal_3520), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1244_s_current_state_reg ( .D(
        new_AGEMA_signal_1766), .CK(clk), .Q(new_AGEMA_signal_3522), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1246_s_current_state_reg ( .D(
        new_AGEMA_signal_1767), .CK(clk), .Q(new_AGEMA_signal_3524), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1248_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_L1), .CK(clk), .Q(new_AGEMA_signal_3526), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1250_s_current_state_reg ( .D(
        new_AGEMA_signal_1948), .CK(clk), .Q(new_AGEMA_signal_3528), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1252_s_current_state_reg ( .D(
        new_AGEMA_signal_1949), .CK(clk), .Q(new_AGEMA_signal_3530), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1254_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_XX_2_), .CK(clk), .Q(new_AGEMA_signal_3532), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1256_s_current_state_reg ( .D(
        new_AGEMA_signal_1198), .CK(clk), .Q(new_AGEMA_signal_3534), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1258_s_current_state_reg ( .D(
        new_AGEMA_signal_1199), .CK(clk), .Q(new_AGEMA_signal_3536), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1260_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_XX_1_), .CK(clk), .Q(new_AGEMA_signal_3538), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1262_s_current_state_reg ( .D(
        new_AGEMA_signal_1194), .CK(clk), .Q(new_AGEMA_signal_3540), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1264_s_current_state_reg ( .D(
        new_AGEMA_signal_1195), .CK(clk), .Q(new_AGEMA_signal_3542), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1266_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_Q0), .CK(clk), .Q(new_AGEMA_signal_3544), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1268_s_current_state_reg ( .D(
        new_AGEMA_signal_1778), .CK(clk), .Q(new_AGEMA_signal_3546), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1270_s_current_state_reg ( .D(
        new_AGEMA_signal_1779), .CK(clk), .Q(new_AGEMA_signal_3548), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1272_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_L1), .CK(clk), .Q(new_AGEMA_signal_3550), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1274_s_current_state_reg ( .D(
        new_AGEMA_signal_1954), .CK(clk), .Q(new_AGEMA_signal_3552), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1276_s_current_state_reg ( .D(
        new_AGEMA_signal_1955), .CK(clk), .Q(new_AGEMA_signal_3554), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1278_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_XX_2_), .CK(clk), .Q(new_AGEMA_signal_3556), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1280_s_current_state_reg ( .D(
        new_AGEMA_signal_1210), .CK(clk), .Q(new_AGEMA_signal_3558), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1282_s_current_state_reg ( .D(
        new_AGEMA_signal_1211), .CK(clk), .Q(new_AGEMA_signal_3560), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1284_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_XX_1_), .CK(clk), .Q(new_AGEMA_signal_3562), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1286_s_current_state_reg ( .D(
        new_AGEMA_signal_1206), .CK(clk), .Q(new_AGEMA_signal_3564), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1288_s_current_state_reg ( .D(
        new_AGEMA_signal_1207), .CK(clk), .Q(new_AGEMA_signal_3566), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1290_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_Q0), .CK(clk), .Q(new_AGEMA_signal_3568), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1292_s_current_state_reg ( .D(
        new_AGEMA_signal_1790), .CK(clk), .Q(new_AGEMA_signal_3570), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1294_s_current_state_reg ( .D(
        new_AGEMA_signal_1791), .CK(clk), .Q(new_AGEMA_signal_3572), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1296_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_L1), .CK(clk), .Q(new_AGEMA_signal_3574), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1298_s_current_state_reg ( .D(
        new_AGEMA_signal_1960), .CK(clk), .Q(new_AGEMA_signal_3576), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1300_s_current_state_reg ( .D(
        new_AGEMA_signal_1961), .CK(clk), .Q(new_AGEMA_signal_3578), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1302_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_XX_2_), .CK(clk), .Q(new_AGEMA_signal_3580), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1304_s_current_state_reg ( .D(
        new_AGEMA_signal_1222), .CK(clk), .Q(new_AGEMA_signal_3582), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1306_s_current_state_reg ( .D(
        new_AGEMA_signal_1223), .CK(clk), .Q(new_AGEMA_signal_3584), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1308_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_XX_1_), .CK(clk), .Q(new_AGEMA_signal_3586), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1310_s_current_state_reg ( .D(
        new_AGEMA_signal_1218), .CK(clk), .Q(new_AGEMA_signal_3588), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1312_s_current_state_reg ( .D(
        new_AGEMA_signal_1219), .CK(clk), .Q(new_AGEMA_signal_3590), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1314_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_Q0), .CK(clk), .Q(new_AGEMA_signal_3592), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1316_s_current_state_reg ( .D(
        new_AGEMA_signal_1802), .CK(clk), .Q(new_AGEMA_signal_3594), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1318_s_current_state_reg ( .D(
        new_AGEMA_signal_1803), .CK(clk), .Q(new_AGEMA_signal_3596), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1320_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_L1), .CK(clk), .Q(new_AGEMA_signal_3598), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1322_s_current_state_reg ( .D(
        new_AGEMA_signal_1966), .CK(clk), .Q(new_AGEMA_signal_3600), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1324_s_current_state_reg ( .D(
        new_AGEMA_signal_1967), .CK(clk), .Q(new_AGEMA_signal_3602), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1326_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_XX_2_), .CK(clk), .Q(new_AGEMA_signal_3604), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1328_s_current_state_reg ( .D(
        new_AGEMA_signal_1234), .CK(clk), .Q(new_AGEMA_signal_3606), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1330_s_current_state_reg ( .D(
        new_AGEMA_signal_1235), .CK(clk), .Q(new_AGEMA_signal_3608), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1332_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_XX_1_), .CK(clk), .Q(new_AGEMA_signal_3610), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1334_s_current_state_reg ( .D(
        new_AGEMA_signal_1230), .CK(clk), .Q(new_AGEMA_signal_3612), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1336_s_current_state_reg ( .D(
        new_AGEMA_signal_1231), .CK(clk), .Q(new_AGEMA_signal_3614), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1338_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_Q0), .CK(clk), .Q(new_AGEMA_signal_3616), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1340_s_current_state_reg ( .D(
        new_AGEMA_signal_1814), .CK(clk), .Q(new_AGEMA_signal_3618), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1342_s_current_state_reg ( .D(
        new_AGEMA_signal_1815), .CK(clk), .Q(new_AGEMA_signal_3620), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1344_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_L1), .CK(clk), .Q(new_AGEMA_signal_3622), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1346_s_current_state_reg ( .D(
        new_AGEMA_signal_1972), .CK(clk), .Q(new_AGEMA_signal_3624), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1348_s_current_state_reg ( .D(
        new_AGEMA_signal_1973), .CK(clk), .Q(new_AGEMA_signal_3626), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1350_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_XX_2_), .CK(clk), .Q(new_AGEMA_signal_3628), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1352_s_current_state_reg ( .D(
        new_AGEMA_signal_1246), .CK(clk), .Q(new_AGEMA_signal_3630), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1354_s_current_state_reg ( .D(
        new_AGEMA_signal_1247), .CK(clk), .Q(new_AGEMA_signal_3632), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1356_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_XX_1_), .CK(clk), .Q(new_AGEMA_signal_3634), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1358_s_current_state_reg ( .D(
        new_AGEMA_signal_1242), .CK(clk), .Q(new_AGEMA_signal_3636), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1360_s_current_state_reg ( .D(
        new_AGEMA_signal_1243), .CK(clk), .Q(new_AGEMA_signal_3638), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1362_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_Q0), .CK(clk), .Q(new_AGEMA_signal_3640), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1364_s_current_state_reg ( .D(
        new_AGEMA_signal_1826), .CK(clk), .Q(new_AGEMA_signal_3642), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1366_s_current_state_reg ( .D(
        new_AGEMA_signal_1827), .CK(clk), .Q(new_AGEMA_signal_3644), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1368_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_L1), .CK(clk), .Q(new_AGEMA_signal_3646), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1370_s_current_state_reg ( .D(
        new_AGEMA_signal_1978), .CK(clk), .Q(new_AGEMA_signal_3648), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1372_s_current_state_reg ( .D(
        new_AGEMA_signal_1979), .CK(clk), .Q(new_AGEMA_signal_3650), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1374_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_XX_2_), .CK(clk), .Q(new_AGEMA_signal_3652), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1376_s_current_state_reg ( .D(
        new_AGEMA_signal_1258), .CK(clk), .Q(new_AGEMA_signal_3654), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1378_s_current_state_reg ( .D(
        new_AGEMA_signal_1259), .CK(clk), .Q(new_AGEMA_signal_3656), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1380_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_XX_1_), .CK(clk), .Q(new_AGEMA_signal_3658), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1382_s_current_state_reg ( .D(
        new_AGEMA_signal_1254), .CK(clk), .Q(new_AGEMA_signal_3660), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1384_s_current_state_reg ( .D(
        new_AGEMA_signal_1255), .CK(clk), .Q(new_AGEMA_signal_3662), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1386_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_Q0), .CK(clk), .Q(new_AGEMA_signal_3664), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1388_s_current_state_reg ( .D(
        new_AGEMA_signal_1838), .CK(clk), .Q(new_AGEMA_signal_3666), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1390_s_current_state_reg ( .D(
        new_AGEMA_signal_1839), .CK(clk), .Q(new_AGEMA_signal_3668), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1392_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_L1), .CK(clk), .Q(new_AGEMA_signal_3670), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1394_s_current_state_reg ( .D(
        new_AGEMA_signal_1984), .CK(clk), .Q(new_AGEMA_signal_3672), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1396_s_current_state_reg ( .D(
        new_AGEMA_signal_1985), .CK(clk), .Q(new_AGEMA_signal_3674), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1398_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_XX_2_), .CK(clk), .Q(new_AGEMA_signal_3676), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1400_s_current_state_reg ( .D(
        new_AGEMA_signal_1270), .CK(clk), .Q(new_AGEMA_signal_3678), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1402_s_current_state_reg ( .D(
        new_AGEMA_signal_1271), .CK(clk), .Q(new_AGEMA_signal_3680), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1404_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_XX_1_), .CK(clk), .Q(new_AGEMA_signal_3682), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1406_s_current_state_reg ( .D(
        new_AGEMA_signal_1266), .CK(clk), .Q(new_AGEMA_signal_3684), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1408_s_current_state_reg ( .D(
        new_AGEMA_signal_1267), .CK(clk), .Q(new_AGEMA_signal_3686), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1410_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_Q0), .CK(clk), .Q(new_AGEMA_signal_3688), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1412_s_current_state_reg ( .D(
        new_AGEMA_signal_1850), .CK(clk), .Q(new_AGEMA_signal_3690), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1414_s_current_state_reg ( .D(
        new_AGEMA_signal_1851), .CK(clk), .Q(new_AGEMA_signal_3692), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1416_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_L1), .CK(clk), .Q(new_AGEMA_signal_3694), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_1418_s_current_state_reg ( .D(
        new_AGEMA_signal_1990), .CK(clk), .Q(new_AGEMA_signal_3696), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1420_s_current_state_reg ( .D(
        new_AGEMA_signal_1991), .CK(clk), .Q(new_AGEMA_signal_3698), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1422_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_XX_2_), .CK(clk), .Q(new_AGEMA_signal_3700), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1424_s_current_state_reg ( .D(
        new_AGEMA_signal_1282), .CK(clk), .Q(new_AGEMA_signal_3702), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1426_s_current_state_reg ( .D(
        new_AGEMA_signal_1283), .CK(clk), .Q(new_AGEMA_signal_3704), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1428_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_XX_1_), .CK(clk), .Q(new_AGEMA_signal_3706), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1430_s_current_state_reg ( .D(
        new_AGEMA_signal_1278), .CK(clk), .Q(new_AGEMA_signal_3708), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1432_s_current_state_reg ( .D(
        new_AGEMA_signal_1279), .CK(clk), .Q(new_AGEMA_signal_3710), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1434_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_Q0), .CK(clk), .Q(new_AGEMA_signal_3712), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1436_s_current_state_reg ( .D(
        new_AGEMA_signal_1862), .CK(clk), .Q(new_AGEMA_signal_3714), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1438_s_current_state_reg ( .D(
        new_AGEMA_signal_1863), .CK(clk), .Q(new_AGEMA_signal_3716), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1440_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_L1), .CK(clk), .Q(new_AGEMA_signal_3718), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1442_s_current_state_reg ( .D(
        new_AGEMA_signal_1996), .CK(clk), .Q(new_AGEMA_signal_3720), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1444_s_current_state_reg ( .D(
        new_AGEMA_signal_1997), .CK(clk), .Q(new_AGEMA_signal_3722), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1446_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_XX_2_), .CK(clk), .Q(new_AGEMA_signal_3724), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1448_s_current_state_reg ( .D(
        new_AGEMA_signal_1294), .CK(clk), .Q(new_AGEMA_signal_3726), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1450_s_current_state_reg ( .D(
        new_AGEMA_signal_1295), .CK(clk), .Q(new_AGEMA_signal_3728), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1452_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_XX_1_), .CK(clk), .Q(new_AGEMA_signal_3730), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1454_s_current_state_reg ( .D(
        new_AGEMA_signal_1290), .CK(clk), .Q(new_AGEMA_signal_3732), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1456_s_current_state_reg ( .D(
        new_AGEMA_signal_1291), .CK(clk), .Q(new_AGEMA_signal_3734), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1458_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_Q0), .CK(clk), .Q(new_AGEMA_signal_3736), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1460_s_current_state_reg ( .D(
        new_AGEMA_signal_1874), .CK(clk), .Q(new_AGEMA_signal_3738), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1462_s_current_state_reg ( .D(
        new_AGEMA_signal_1875), .CK(clk), .Q(new_AGEMA_signal_3740), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1464_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_L1), .CK(clk), .Q(new_AGEMA_signal_3742), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1466_s_current_state_reg ( .D(
        new_AGEMA_signal_2002), .CK(clk), .Q(new_AGEMA_signal_3744), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1468_s_current_state_reg ( .D(
        new_AGEMA_signal_2003), .CK(clk), .Q(new_AGEMA_signal_3746), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1470_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_XX_2_), .CK(clk), .Q(new_AGEMA_signal_3748), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1472_s_current_state_reg ( .D(
        new_AGEMA_signal_1306), .CK(clk), .Q(new_AGEMA_signal_3750), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1474_s_current_state_reg ( .D(
        new_AGEMA_signal_1307), .CK(clk), .Q(new_AGEMA_signal_3752), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1476_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_XX_1_), .CK(clk), .Q(new_AGEMA_signal_3754), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1478_s_current_state_reg ( .D(
        new_AGEMA_signal_1302), .CK(clk), .Q(new_AGEMA_signal_3756), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1480_s_current_state_reg ( .D(
        new_AGEMA_signal_1303), .CK(clk), .Q(new_AGEMA_signal_3758), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1482_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_Q0), .CK(clk), .Q(new_AGEMA_signal_3760), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1484_s_current_state_reg ( .D(
        new_AGEMA_signal_1886), .CK(clk), .Q(new_AGEMA_signal_3762), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1486_s_current_state_reg ( .D(
        new_AGEMA_signal_1887), .CK(clk), .Q(new_AGEMA_signal_3764), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1488_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_L1), .CK(clk), .Q(new_AGEMA_signal_3766), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1490_s_current_state_reg ( .D(
        new_AGEMA_signal_2008), .CK(clk), .Q(new_AGEMA_signal_3768), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1492_s_current_state_reg ( .D(
        new_AGEMA_signal_2009), .CK(clk), .Q(new_AGEMA_signal_3770), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1494_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_XX_2_), .CK(clk), .Q(new_AGEMA_signal_3772), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1496_s_current_state_reg ( .D(
        new_AGEMA_signal_1318), .CK(clk), .Q(new_AGEMA_signal_3774), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1498_s_current_state_reg ( .D(
        new_AGEMA_signal_1319), .CK(clk), .Q(new_AGEMA_signal_3776), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1500_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_XX_1_), .CK(clk), .Q(new_AGEMA_signal_3778), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1502_s_current_state_reg ( .D(
        new_AGEMA_signal_1314), .CK(clk), .Q(new_AGEMA_signal_3780), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1504_s_current_state_reg ( .D(
        new_AGEMA_signal_1315), .CK(clk), .Q(new_AGEMA_signal_3782), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1506_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_Q0), .CK(clk), .Q(new_AGEMA_signal_3784), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1508_s_current_state_reg ( .D(
        new_AGEMA_signal_1898), .CK(clk), .Q(new_AGEMA_signal_3786), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1510_s_current_state_reg ( .D(
        new_AGEMA_signal_1899), .CK(clk), .Q(new_AGEMA_signal_3788), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1512_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_L1), .CK(clk), .Q(new_AGEMA_signal_3790), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1514_s_current_state_reg ( .D(
        new_AGEMA_signal_2014), .CK(clk), .Q(new_AGEMA_signal_3792), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1516_s_current_state_reg ( .D(
        new_AGEMA_signal_2015), .CK(clk), .Q(new_AGEMA_signal_3794), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1518_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_XX_2_), .CK(clk), .Q(new_AGEMA_signal_3796), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1520_s_current_state_reg ( .D(
        new_AGEMA_signal_1330), .CK(clk), .Q(new_AGEMA_signal_3798), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1522_s_current_state_reg ( .D(
        new_AGEMA_signal_1331), .CK(clk), .Q(new_AGEMA_signal_3800), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1524_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_XX_1_), .CK(clk), .Q(new_AGEMA_signal_3802), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1526_s_current_state_reg ( .D(
        new_AGEMA_signal_1326), .CK(clk), .Q(new_AGEMA_signal_3804), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1528_s_current_state_reg ( .D(
        new_AGEMA_signal_1327), .CK(clk), .Q(new_AGEMA_signal_3806), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1530_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_Q0), .CK(clk), .Q(new_AGEMA_signal_3808), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1532_s_current_state_reg ( .D(
        new_AGEMA_signal_1910), .CK(clk), .Q(new_AGEMA_signal_3810), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1534_s_current_state_reg ( .D(
        new_AGEMA_signal_1911), .CK(clk), .Q(new_AGEMA_signal_3812), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1536_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_L1), .CK(clk), .Q(new_AGEMA_signal_3814), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1538_s_current_state_reg ( .D(
        new_AGEMA_signal_2020), .CK(clk), .Q(new_AGEMA_signal_3816), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1540_s_current_state_reg ( .D(
        new_AGEMA_signal_2021), .CK(clk), .Q(new_AGEMA_signal_3818), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1542_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_XX_2_), .CK(clk), .Q(new_AGEMA_signal_3820), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1544_s_current_state_reg ( .D(
        new_AGEMA_signal_1342), .CK(clk), .Q(new_AGEMA_signal_3822), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1546_s_current_state_reg ( .D(
        new_AGEMA_signal_1343), .CK(clk), .Q(new_AGEMA_signal_3824), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1548_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_XX_1_), .CK(clk), .Q(new_AGEMA_signal_3826), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1550_s_current_state_reg ( .D(
        new_AGEMA_signal_1338), .CK(clk), .Q(new_AGEMA_signal_3828), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1552_s_current_state_reg ( .D(
        new_AGEMA_signal_1339), .CK(clk), .Q(new_AGEMA_signal_3830), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1554_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_Q0), .CK(clk), .Q(new_AGEMA_signal_3832), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1556_s_current_state_reg ( .D(
        new_AGEMA_signal_1922), .CK(clk), .Q(new_AGEMA_signal_3834), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1558_s_current_state_reg ( .D(
        new_AGEMA_signal_1923), .CK(clk), .Q(new_AGEMA_signal_3836), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1560_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_L1), .CK(clk), .Q(new_AGEMA_signal_3838), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1562_s_current_state_reg ( .D(
        new_AGEMA_signal_2026), .CK(clk), .Q(new_AGEMA_signal_3840), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1564_s_current_state_reg ( .D(
        new_AGEMA_signal_2027), .CK(clk), .Q(new_AGEMA_signal_3842), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1566_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_XX_2_), .CK(clk), .Q(new_AGEMA_signal_3844), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1568_s_current_state_reg ( .D(
        new_AGEMA_signal_1354), .CK(clk), .Q(new_AGEMA_signal_3846), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1570_s_current_state_reg ( .D(
        new_AGEMA_signal_1355), .CK(clk), .Q(new_AGEMA_signal_3848), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1572_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_XX_1_), .CK(clk), .Q(new_AGEMA_signal_3850), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1574_s_current_state_reg ( .D(
        new_AGEMA_signal_1350), .CK(clk), .Q(new_AGEMA_signal_3852), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1576_s_current_state_reg ( .D(
        new_AGEMA_signal_1351), .CK(clk), .Q(new_AGEMA_signal_3854), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1578_s_current_state_reg ( .D(FSMUpdate[3]), 
        .CK(clk), .Q(new_AGEMA_signal_3856), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1580_s_current_state_reg ( .D(FSMUpdate[4]), 
        .CK(clk), .Q(new_AGEMA_signal_3858), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1582_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[2]), .CK(clk), .Q(new_AGEMA_signal_3860), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1584_s_current_state_reg ( .D(
        new_AGEMA_signal_1368), .CK(clk), .Q(new_AGEMA_signal_3862), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1586_s_current_state_reg ( .D(
        new_AGEMA_signal_1369), .CK(clk), .Q(new_AGEMA_signal_3864), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1588_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[3]), .CK(clk), .Q(new_AGEMA_signal_3866), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1590_s_current_state_reg ( .D(
        new_AGEMA_signal_1374), .CK(clk), .Q(new_AGEMA_signal_3868), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1592_s_current_state_reg ( .D(
        new_AGEMA_signal_1375), .CK(clk), .Q(new_AGEMA_signal_3870), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1594_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[6]), .CK(clk), .Q(new_AGEMA_signal_3872), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1596_s_current_state_reg ( .D(
        new_AGEMA_signal_1392), .CK(clk), .Q(new_AGEMA_signal_3874), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1598_s_current_state_reg ( .D(
        new_AGEMA_signal_1393), .CK(clk), .Q(new_AGEMA_signal_3876), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1600_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[7]), .CK(clk), .Q(new_AGEMA_signal_3878), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1602_s_current_state_reg ( .D(
        new_AGEMA_signal_1398), .CK(clk), .Q(new_AGEMA_signal_3880), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1604_s_current_state_reg ( .D(
        new_AGEMA_signal_1399), .CK(clk), .Q(new_AGEMA_signal_3882), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1606_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[10]), .CK(clk), .Q(
        new_AGEMA_signal_3884), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1608_s_current_state_reg ( .D(
        new_AGEMA_signal_1416), .CK(clk), .Q(new_AGEMA_signal_3886), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1610_s_current_state_reg ( .D(
        new_AGEMA_signal_1417), .CK(clk), .Q(new_AGEMA_signal_3888), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1612_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[11]), .CK(clk), .Q(
        new_AGEMA_signal_3890), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1614_s_current_state_reg ( .D(
        new_AGEMA_signal_1422), .CK(clk), .Q(new_AGEMA_signal_3892), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1616_s_current_state_reg ( .D(
        new_AGEMA_signal_1423), .CK(clk), .Q(new_AGEMA_signal_3894), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1618_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[14]), .CK(clk), .Q(
        new_AGEMA_signal_3896), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1620_s_current_state_reg ( .D(
        new_AGEMA_signal_1440), .CK(clk), .Q(new_AGEMA_signal_3898), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1622_s_current_state_reg ( .D(
        new_AGEMA_signal_1441), .CK(clk), .Q(new_AGEMA_signal_3900), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1624_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[15]), .CK(clk), .Q(
        new_AGEMA_signal_3902), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1626_s_current_state_reg ( .D(
        new_AGEMA_signal_1446), .CK(clk), .Q(new_AGEMA_signal_3904), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1628_s_current_state_reg ( .D(
        new_AGEMA_signal_1447), .CK(clk), .Q(new_AGEMA_signal_3906), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1630_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[18]), .CK(clk), .Q(
        new_AGEMA_signal_3908), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1632_s_current_state_reg ( .D(
        new_AGEMA_signal_1464), .CK(clk), .Q(new_AGEMA_signal_3910), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1634_s_current_state_reg ( .D(
        new_AGEMA_signal_1465), .CK(clk), .Q(new_AGEMA_signal_3912), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1636_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[19]), .CK(clk), .Q(
        new_AGEMA_signal_3914), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1638_s_current_state_reg ( .D(
        new_AGEMA_signal_1470), .CK(clk), .Q(new_AGEMA_signal_3916), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1640_s_current_state_reg ( .D(
        new_AGEMA_signal_1471), .CK(clk), .Q(new_AGEMA_signal_3918), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1642_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[22]), .CK(clk), .Q(
        new_AGEMA_signal_3920), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1644_s_current_state_reg ( .D(
        new_AGEMA_signal_1488), .CK(clk), .Q(new_AGEMA_signal_3922), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1646_s_current_state_reg ( .D(
        new_AGEMA_signal_1489), .CK(clk), .Q(new_AGEMA_signal_3924), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1648_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[23]), .CK(clk), .Q(
        new_AGEMA_signal_3926), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1650_s_current_state_reg ( .D(
        new_AGEMA_signal_1494), .CK(clk), .Q(new_AGEMA_signal_3928), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1652_s_current_state_reg ( .D(
        new_AGEMA_signal_1495), .CK(clk), .Q(new_AGEMA_signal_3930), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1654_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[26]), .CK(clk), .Q(
        new_AGEMA_signal_3932), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1656_s_current_state_reg ( .D(
        new_AGEMA_signal_1512), .CK(clk), .Q(new_AGEMA_signal_3934), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1658_s_current_state_reg ( .D(
        new_AGEMA_signal_1513), .CK(clk), .Q(new_AGEMA_signal_3936), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1660_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[27]), .CK(clk), .Q(
        new_AGEMA_signal_3938), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1662_s_current_state_reg ( .D(
        new_AGEMA_signal_1518), .CK(clk), .Q(new_AGEMA_signal_3940), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1664_s_current_state_reg ( .D(
        new_AGEMA_signal_1519), .CK(clk), .Q(new_AGEMA_signal_3942), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1666_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[30]), .CK(clk), .Q(
        new_AGEMA_signal_3944), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1668_s_current_state_reg ( .D(
        new_AGEMA_signal_1536), .CK(clk), .Q(new_AGEMA_signal_3946), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1670_s_current_state_reg ( .D(
        new_AGEMA_signal_1537), .CK(clk), .Q(new_AGEMA_signal_3948), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1672_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[31]), .CK(clk), .Q(
        new_AGEMA_signal_3950), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1674_s_current_state_reg ( .D(
        new_AGEMA_signal_1542), .CK(clk), .Q(new_AGEMA_signal_3952), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1676_s_current_state_reg ( .D(
        new_AGEMA_signal_1543), .CK(clk), .Q(new_AGEMA_signal_3954), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1680_s_current_state_reg ( .D(Plaintext_s0[0]), 
        .CK(clk), .Q(new_AGEMA_signal_3958), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1684_s_current_state_reg ( .D(Plaintext_s1[0]), 
        .CK(clk), .Q(new_AGEMA_signal_3962), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1688_s_current_state_reg ( .D(Plaintext_s2[0]), 
        .CK(clk), .Q(new_AGEMA_signal_3966), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1692_s_current_state_reg ( .D(Plaintext_s0[1]), 
        .CK(clk), .Q(new_AGEMA_signal_3970), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1696_s_current_state_reg ( .D(Plaintext_s1[1]), 
        .CK(clk), .Q(new_AGEMA_signal_3974), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1700_s_current_state_reg ( .D(Plaintext_s2[1]), 
        .CK(clk), .Q(new_AGEMA_signal_3978), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1704_s_current_state_reg ( .D(Plaintext_s0[4]), 
        .CK(clk), .Q(new_AGEMA_signal_3982), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1708_s_current_state_reg ( .D(Plaintext_s1[4]), 
        .CK(clk), .Q(new_AGEMA_signal_3986), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1712_s_current_state_reg ( .D(Plaintext_s2[4]), 
        .CK(clk), .Q(new_AGEMA_signal_3990), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1716_s_current_state_reg ( .D(Plaintext_s0[5]), 
        .CK(clk), .Q(new_AGEMA_signal_3994), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1720_s_current_state_reg ( .D(Plaintext_s1[5]), 
        .CK(clk), .Q(new_AGEMA_signal_3998), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1724_s_current_state_reg ( .D(Plaintext_s2[5]), 
        .CK(clk), .Q(new_AGEMA_signal_4002), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1728_s_current_state_reg ( .D(Plaintext_s0[8]), 
        .CK(clk), .Q(new_AGEMA_signal_4006), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1732_s_current_state_reg ( .D(Plaintext_s1[8]), 
        .CK(clk), .Q(new_AGEMA_signal_4010), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1736_s_current_state_reg ( .D(Plaintext_s2[8]), 
        .CK(clk), .Q(new_AGEMA_signal_4014), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1740_s_current_state_reg ( .D(Plaintext_s0[9]), 
        .CK(clk), .Q(new_AGEMA_signal_4018), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1744_s_current_state_reg ( .D(Plaintext_s1[9]), 
        .CK(clk), .Q(new_AGEMA_signal_4022), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1748_s_current_state_reg ( .D(Plaintext_s2[9]), 
        .CK(clk), .Q(new_AGEMA_signal_4026), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1752_s_current_state_reg ( .D(Plaintext_s0[12]), 
        .CK(clk), .Q(new_AGEMA_signal_4030), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1756_s_current_state_reg ( .D(Plaintext_s1[12]), 
        .CK(clk), .Q(new_AGEMA_signal_4034), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1760_s_current_state_reg ( .D(Plaintext_s2[12]), 
        .CK(clk), .Q(new_AGEMA_signal_4038), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1764_s_current_state_reg ( .D(Plaintext_s0[13]), 
        .CK(clk), .Q(new_AGEMA_signal_4042), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1768_s_current_state_reg ( .D(Plaintext_s1[13]), 
        .CK(clk), .Q(new_AGEMA_signal_4046), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1772_s_current_state_reg ( .D(Plaintext_s2[13]), 
        .CK(clk), .Q(new_AGEMA_signal_4050), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1776_s_current_state_reg ( .D(Plaintext_s0[16]), 
        .CK(clk), .Q(new_AGEMA_signal_4054), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1780_s_current_state_reg ( .D(Plaintext_s1[16]), 
        .CK(clk), .Q(new_AGEMA_signal_4058), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1784_s_current_state_reg ( .D(Plaintext_s2[16]), 
        .CK(clk), .Q(new_AGEMA_signal_4062), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1788_s_current_state_reg ( .D(Plaintext_s0[17]), 
        .CK(clk), .Q(new_AGEMA_signal_4066), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1792_s_current_state_reg ( .D(Plaintext_s1[17]), 
        .CK(clk), .Q(new_AGEMA_signal_4070), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1796_s_current_state_reg ( .D(Plaintext_s2[17]), 
        .CK(clk), .Q(new_AGEMA_signal_4074), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1800_s_current_state_reg ( .D(Plaintext_s0[20]), 
        .CK(clk), .Q(new_AGEMA_signal_4078), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1804_s_current_state_reg ( .D(Plaintext_s1[20]), 
        .CK(clk), .Q(new_AGEMA_signal_4082), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1808_s_current_state_reg ( .D(Plaintext_s2[20]), 
        .CK(clk), .Q(new_AGEMA_signal_4086), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1812_s_current_state_reg ( .D(Plaintext_s0[21]), 
        .CK(clk), .Q(new_AGEMA_signal_4090), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1816_s_current_state_reg ( .D(Plaintext_s1[21]), 
        .CK(clk), .Q(new_AGEMA_signal_4094), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1820_s_current_state_reg ( .D(Plaintext_s2[21]), 
        .CK(clk), .Q(new_AGEMA_signal_4098), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1824_s_current_state_reg ( .D(Plaintext_s0[24]), 
        .CK(clk), .Q(new_AGEMA_signal_4102), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1828_s_current_state_reg ( .D(Plaintext_s1[24]), 
        .CK(clk), .Q(new_AGEMA_signal_4106), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1832_s_current_state_reg ( .D(Plaintext_s2[24]), 
        .CK(clk), .Q(new_AGEMA_signal_4110), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1836_s_current_state_reg ( .D(Plaintext_s0[25]), 
        .CK(clk), .Q(new_AGEMA_signal_4114), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1840_s_current_state_reg ( .D(Plaintext_s1[25]), 
        .CK(clk), .Q(new_AGEMA_signal_4118), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1844_s_current_state_reg ( .D(Plaintext_s2[25]), 
        .CK(clk), .Q(new_AGEMA_signal_4122), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1848_s_current_state_reg ( .D(Plaintext_s0[28]), 
        .CK(clk), .Q(new_AGEMA_signal_4126), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1852_s_current_state_reg ( .D(Plaintext_s1[28]), 
        .CK(clk), .Q(new_AGEMA_signal_4130), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1856_s_current_state_reg ( .D(Plaintext_s2[28]), 
        .CK(clk), .Q(new_AGEMA_signal_4134), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1860_s_current_state_reg ( .D(Plaintext_s0[29]), 
        .CK(clk), .Q(new_AGEMA_signal_4138), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1864_s_current_state_reg ( .D(Plaintext_s1[29]), 
        .CK(clk), .Q(new_AGEMA_signal_4142), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1868_s_current_state_reg ( .D(Plaintext_s2[29]), 
        .CK(clk), .Q(new_AGEMA_signal_4146), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1872_s_current_state_reg ( .D(Plaintext_s0[32]), 
        .CK(clk), .Q(new_AGEMA_signal_4150), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1876_s_current_state_reg ( .D(Plaintext_s1[32]), 
        .CK(clk), .Q(new_AGEMA_signal_4154), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1880_s_current_state_reg ( .D(Plaintext_s2[32]), 
        .CK(clk), .Q(new_AGEMA_signal_4158), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1884_s_current_state_reg ( .D(Plaintext_s0[33]), 
        .CK(clk), .Q(new_AGEMA_signal_4162), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1888_s_current_state_reg ( .D(Plaintext_s1[33]), 
        .CK(clk), .Q(new_AGEMA_signal_4166), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1892_s_current_state_reg ( .D(Plaintext_s2[33]), 
        .CK(clk), .Q(new_AGEMA_signal_4170), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1896_s_current_state_reg ( .D(Plaintext_s0[36]), 
        .CK(clk), .Q(new_AGEMA_signal_4174), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1900_s_current_state_reg ( .D(Plaintext_s1[36]), 
        .CK(clk), .Q(new_AGEMA_signal_4178), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1904_s_current_state_reg ( .D(Plaintext_s2[36]), 
        .CK(clk), .Q(new_AGEMA_signal_4182), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1908_s_current_state_reg ( .D(Plaintext_s0[37]), 
        .CK(clk), .Q(new_AGEMA_signal_4186), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1912_s_current_state_reg ( .D(Plaintext_s1[37]), 
        .CK(clk), .Q(new_AGEMA_signal_4190), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1916_s_current_state_reg ( .D(Plaintext_s2[37]), 
        .CK(clk), .Q(new_AGEMA_signal_4194), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1920_s_current_state_reg ( .D(Plaintext_s0[40]), 
        .CK(clk), .Q(new_AGEMA_signal_4198), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1924_s_current_state_reg ( .D(Plaintext_s1[40]), 
        .CK(clk), .Q(new_AGEMA_signal_4202), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1928_s_current_state_reg ( .D(Plaintext_s2[40]), 
        .CK(clk), .Q(new_AGEMA_signal_4206), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1932_s_current_state_reg ( .D(Plaintext_s0[41]), 
        .CK(clk), .Q(new_AGEMA_signal_4210), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1936_s_current_state_reg ( .D(Plaintext_s1[41]), 
        .CK(clk), .Q(new_AGEMA_signal_4214), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1940_s_current_state_reg ( .D(Plaintext_s2[41]), 
        .CK(clk), .Q(new_AGEMA_signal_4218), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1944_s_current_state_reg ( .D(Plaintext_s0[44]), 
        .CK(clk), .Q(new_AGEMA_signal_4222), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1948_s_current_state_reg ( .D(Plaintext_s1[44]), 
        .CK(clk), .Q(new_AGEMA_signal_4226), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1952_s_current_state_reg ( .D(Plaintext_s2[44]), 
        .CK(clk), .Q(new_AGEMA_signal_4230), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1956_s_current_state_reg ( .D(Plaintext_s0[45]), 
        .CK(clk), .Q(new_AGEMA_signal_4234), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1960_s_current_state_reg ( .D(Plaintext_s1[45]), 
        .CK(clk), .Q(new_AGEMA_signal_4238), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1964_s_current_state_reg ( .D(Plaintext_s2[45]), 
        .CK(clk), .Q(new_AGEMA_signal_4242), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1968_s_current_state_reg ( .D(Plaintext_s0[48]), 
        .CK(clk), .Q(new_AGEMA_signal_4246), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1972_s_current_state_reg ( .D(Plaintext_s1[48]), 
        .CK(clk), .Q(new_AGEMA_signal_4250), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1976_s_current_state_reg ( .D(Plaintext_s2[48]), 
        .CK(clk), .Q(new_AGEMA_signal_4254), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1980_s_current_state_reg ( .D(Plaintext_s0[49]), 
        .CK(clk), .Q(new_AGEMA_signal_4258), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1984_s_current_state_reg ( .D(Plaintext_s1[49]), 
        .CK(clk), .Q(new_AGEMA_signal_4262), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1988_s_current_state_reg ( .D(Plaintext_s2[49]), 
        .CK(clk), .Q(new_AGEMA_signal_4266), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1992_s_current_state_reg ( .D(Plaintext_s0[52]), 
        .CK(clk), .Q(new_AGEMA_signal_4270), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1996_s_current_state_reg ( .D(Plaintext_s1[52]), 
        .CK(clk), .Q(new_AGEMA_signal_4274), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2000_s_current_state_reg ( .D(Plaintext_s2[52]), 
        .CK(clk), .Q(new_AGEMA_signal_4278), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2004_s_current_state_reg ( .D(Plaintext_s0[53]), 
        .CK(clk), .Q(new_AGEMA_signal_4282), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2008_s_current_state_reg ( .D(Plaintext_s1[53]), 
        .CK(clk), .Q(new_AGEMA_signal_4286), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2012_s_current_state_reg ( .D(Plaintext_s2[53]), 
        .CK(clk), .Q(new_AGEMA_signal_4290), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2016_s_current_state_reg ( .D(Plaintext_s0[56]), 
        .CK(clk), .Q(new_AGEMA_signal_4294), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2020_s_current_state_reg ( .D(Plaintext_s1[56]), 
        .CK(clk), .Q(new_AGEMA_signal_4298), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2024_s_current_state_reg ( .D(Plaintext_s2[56]), 
        .CK(clk), .Q(new_AGEMA_signal_4302), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2028_s_current_state_reg ( .D(Plaintext_s0[57]), 
        .CK(clk), .Q(new_AGEMA_signal_4306), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2032_s_current_state_reg ( .D(Plaintext_s1[57]), 
        .CK(clk), .Q(new_AGEMA_signal_4310), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2036_s_current_state_reg ( .D(Plaintext_s2[57]), 
        .CK(clk), .Q(new_AGEMA_signal_4314), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2040_s_current_state_reg ( .D(Plaintext_s0[60]), 
        .CK(clk), .Q(new_AGEMA_signal_4318), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2044_s_current_state_reg ( .D(Plaintext_s1[60]), 
        .CK(clk), .Q(new_AGEMA_signal_4322), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2048_s_current_state_reg ( .D(Plaintext_s2[60]), 
        .CK(clk), .Q(new_AGEMA_signal_4326), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2052_s_current_state_reg ( .D(Plaintext_s0[61]), 
        .CK(clk), .Q(new_AGEMA_signal_4330), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2056_s_current_state_reg ( .D(Plaintext_s1[61]), 
        .CK(clk), .Q(new_AGEMA_signal_4334), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2060_s_current_state_reg ( .D(Plaintext_s2[61]), 
        .CK(clk), .Q(new_AGEMA_signal_4338), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2064_s_current_state_reg ( .D(Ciphertext_s0[1]), 
        .CK(clk), .Q(new_AGEMA_signal_4342), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2066_s_current_state_reg ( .D(Ciphertext_s1[1]), 
        .CK(clk), .Q(new_AGEMA_signal_4344), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2068_s_current_state_reg ( .D(Ciphertext_s2[1]), 
        .CK(clk), .Q(new_AGEMA_signal_4346), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2076_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_Q6), .CK(clk), .Q(new_AGEMA_signal_4354), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2078_s_current_state_reg ( .D(
        new_AGEMA_signal_1748), .CK(clk), .Q(new_AGEMA_signal_4356), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2080_s_current_state_reg ( .D(
        new_AGEMA_signal_1749), .CK(clk), .Q(new_AGEMA_signal_4358), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2082_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_L2), .CK(clk), .Q(new_AGEMA_signal_4360), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2086_s_current_state_reg ( .D(
        new_AGEMA_signal_1750), .CK(clk), .Q(new_AGEMA_signal_4364), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2090_s_current_state_reg ( .D(
        new_AGEMA_signal_1751), .CK(clk), .Q(new_AGEMA_signal_4368), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2100_s_current_state_reg ( .D(Ciphertext_s0[5]), 
        .CK(clk), .Q(new_AGEMA_signal_4378), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2102_s_current_state_reg ( .D(Ciphertext_s1[5]), 
        .CK(clk), .Q(new_AGEMA_signal_4380), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2104_s_current_state_reg ( .D(Ciphertext_s2[5]), 
        .CK(clk), .Q(new_AGEMA_signal_4382), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2112_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_Q6), .CK(clk), .Q(new_AGEMA_signal_4390), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2114_s_current_state_reg ( .D(
        new_AGEMA_signal_1760), .CK(clk), .Q(new_AGEMA_signal_4392), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2116_s_current_state_reg ( .D(
        new_AGEMA_signal_1761), .CK(clk), .Q(new_AGEMA_signal_4394), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2118_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_L2), .CK(clk), .Q(new_AGEMA_signal_4396), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2122_s_current_state_reg ( .D(
        new_AGEMA_signal_1762), .CK(clk), .Q(new_AGEMA_signal_4400), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2126_s_current_state_reg ( .D(
        new_AGEMA_signal_1763), .CK(clk), .Q(new_AGEMA_signal_4404), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2136_s_current_state_reg ( .D(Ciphertext_s0[9]), 
        .CK(clk), .Q(new_AGEMA_signal_4414), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2138_s_current_state_reg ( .D(Ciphertext_s1[9]), 
        .CK(clk), .Q(new_AGEMA_signal_4416), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2140_s_current_state_reg ( .D(Ciphertext_s2[9]), 
        .CK(clk), .Q(new_AGEMA_signal_4418), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2148_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_Q6), .CK(clk), .Q(new_AGEMA_signal_4426), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2150_s_current_state_reg ( .D(
        new_AGEMA_signal_1772), .CK(clk), .Q(new_AGEMA_signal_4428), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2152_s_current_state_reg ( .D(
        new_AGEMA_signal_1773), .CK(clk), .Q(new_AGEMA_signal_4430), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2154_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_L2), .CK(clk), .Q(new_AGEMA_signal_4432), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2158_s_current_state_reg ( .D(
        new_AGEMA_signal_1774), .CK(clk), .Q(new_AGEMA_signal_4436), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2162_s_current_state_reg ( .D(
        new_AGEMA_signal_1775), .CK(clk), .Q(new_AGEMA_signal_4440), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2172_s_current_state_reg ( .D(Ciphertext_s0[13]), 
        .CK(clk), .Q(new_AGEMA_signal_4450), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2174_s_current_state_reg ( .D(Ciphertext_s1[13]), 
        .CK(clk), .Q(new_AGEMA_signal_4452), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2176_s_current_state_reg ( .D(Ciphertext_s2[13]), 
        .CK(clk), .Q(new_AGEMA_signal_4454), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2184_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_Q6), .CK(clk), .Q(new_AGEMA_signal_4462), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2186_s_current_state_reg ( .D(
        new_AGEMA_signal_1784), .CK(clk), .Q(new_AGEMA_signal_4464), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2188_s_current_state_reg ( .D(
        new_AGEMA_signal_1785), .CK(clk), .Q(new_AGEMA_signal_4466), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2190_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_L2), .CK(clk), .Q(new_AGEMA_signal_4468), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2194_s_current_state_reg ( .D(
        new_AGEMA_signal_1786), .CK(clk), .Q(new_AGEMA_signal_4472), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2198_s_current_state_reg ( .D(
        new_AGEMA_signal_1787), .CK(clk), .Q(new_AGEMA_signal_4476), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2208_s_current_state_reg ( .D(Ciphertext_s0[17]), 
        .CK(clk), .Q(new_AGEMA_signal_4486), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2210_s_current_state_reg ( .D(Ciphertext_s1[17]), 
        .CK(clk), .Q(new_AGEMA_signal_4488), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2212_s_current_state_reg ( .D(Ciphertext_s2[17]), 
        .CK(clk), .Q(new_AGEMA_signal_4490), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2220_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_Q6), .CK(clk), .Q(new_AGEMA_signal_4498), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2222_s_current_state_reg ( .D(
        new_AGEMA_signal_1796), .CK(clk), .Q(new_AGEMA_signal_4500), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2224_s_current_state_reg ( .D(
        new_AGEMA_signal_1797), .CK(clk), .Q(new_AGEMA_signal_4502), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2226_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_L2), .CK(clk), .Q(new_AGEMA_signal_4504), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2230_s_current_state_reg ( .D(
        new_AGEMA_signal_1798), .CK(clk), .Q(new_AGEMA_signal_4508), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2234_s_current_state_reg ( .D(
        new_AGEMA_signal_1799), .CK(clk), .Q(new_AGEMA_signal_4512), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2244_s_current_state_reg ( .D(Ciphertext_s0[21]), 
        .CK(clk), .Q(new_AGEMA_signal_4522), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2246_s_current_state_reg ( .D(Ciphertext_s1[21]), 
        .CK(clk), .Q(new_AGEMA_signal_4524), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2248_s_current_state_reg ( .D(Ciphertext_s2[21]), 
        .CK(clk), .Q(new_AGEMA_signal_4526), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2256_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_Q6), .CK(clk), .Q(new_AGEMA_signal_4534), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2258_s_current_state_reg ( .D(
        new_AGEMA_signal_1808), .CK(clk), .Q(new_AGEMA_signal_4536), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2260_s_current_state_reg ( .D(
        new_AGEMA_signal_1809), .CK(clk), .Q(new_AGEMA_signal_4538), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2262_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_L2), .CK(clk), .Q(new_AGEMA_signal_4540), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2266_s_current_state_reg ( .D(
        new_AGEMA_signal_1810), .CK(clk), .Q(new_AGEMA_signal_4544), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2270_s_current_state_reg ( .D(
        new_AGEMA_signal_1811), .CK(clk), .Q(new_AGEMA_signal_4548), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2280_s_current_state_reg ( .D(Ciphertext_s0[25]), 
        .CK(clk), .Q(new_AGEMA_signal_4558), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2282_s_current_state_reg ( .D(Ciphertext_s1[25]), 
        .CK(clk), .Q(new_AGEMA_signal_4560), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2284_s_current_state_reg ( .D(Ciphertext_s2[25]), 
        .CK(clk), .Q(new_AGEMA_signal_4562), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2292_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_Q6), .CK(clk), .Q(new_AGEMA_signal_4570), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2294_s_current_state_reg ( .D(
        new_AGEMA_signal_1820), .CK(clk), .Q(new_AGEMA_signal_4572), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2296_s_current_state_reg ( .D(
        new_AGEMA_signal_1821), .CK(clk), .Q(new_AGEMA_signal_4574), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2298_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_L2), .CK(clk), .Q(new_AGEMA_signal_4576), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2302_s_current_state_reg ( .D(
        new_AGEMA_signal_1822), .CK(clk), .Q(new_AGEMA_signal_4580), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2306_s_current_state_reg ( .D(
        new_AGEMA_signal_1823), .CK(clk), .Q(new_AGEMA_signal_4584), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2316_s_current_state_reg ( .D(Ciphertext_s0[29]), 
        .CK(clk), .Q(new_AGEMA_signal_4594), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2318_s_current_state_reg ( .D(Ciphertext_s1[29]), 
        .CK(clk), .Q(new_AGEMA_signal_4596), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2320_s_current_state_reg ( .D(Ciphertext_s2[29]), 
        .CK(clk), .Q(new_AGEMA_signal_4598), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2328_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_Q6), .CK(clk), .Q(new_AGEMA_signal_4606), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2330_s_current_state_reg ( .D(
        new_AGEMA_signal_1832), .CK(clk), .Q(new_AGEMA_signal_4608), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2332_s_current_state_reg ( .D(
        new_AGEMA_signal_1833), .CK(clk), .Q(new_AGEMA_signal_4610), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2334_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_L2), .CK(clk), .Q(new_AGEMA_signal_4612), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2338_s_current_state_reg ( .D(
        new_AGEMA_signal_1834), .CK(clk), .Q(new_AGEMA_signal_4616), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2342_s_current_state_reg ( .D(
        new_AGEMA_signal_1835), .CK(clk), .Q(new_AGEMA_signal_4620), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2352_s_current_state_reg ( .D(Ciphertext_s0[33]), 
        .CK(clk), .Q(new_AGEMA_signal_4630), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2354_s_current_state_reg ( .D(Ciphertext_s1[33]), 
        .CK(clk), .Q(new_AGEMA_signal_4632), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2356_s_current_state_reg ( .D(Ciphertext_s2[33]), 
        .CK(clk), .Q(new_AGEMA_signal_4634), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2364_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_Q6), .CK(clk), .Q(new_AGEMA_signal_4642), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2366_s_current_state_reg ( .D(
        new_AGEMA_signal_1844), .CK(clk), .Q(new_AGEMA_signal_4644), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2368_s_current_state_reg ( .D(
        new_AGEMA_signal_1845), .CK(clk), .Q(new_AGEMA_signal_4646), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2370_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_L2), .CK(clk), .Q(new_AGEMA_signal_4648), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2374_s_current_state_reg ( .D(
        new_AGEMA_signal_1846), .CK(clk), .Q(new_AGEMA_signal_4652), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2378_s_current_state_reg ( .D(
        new_AGEMA_signal_1847), .CK(clk), .Q(new_AGEMA_signal_4656), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2388_s_current_state_reg ( .D(Ciphertext_s0[37]), 
        .CK(clk), .Q(new_AGEMA_signal_4666), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2390_s_current_state_reg ( .D(Ciphertext_s1[37]), 
        .CK(clk), .Q(new_AGEMA_signal_4668), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2392_s_current_state_reg ( .D(Ciphertext_s2[37]), 
        .CK(clk), .Q(new_AGEMA_signal_4670), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2400_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_Q6), .CK(clk), .Q(new_AGEMA_signal_4678), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2402_s_current_state_reg ( .D(
        new_AGEMA_signal_1856), .CK(clk), .Q(new_AGEMA_signal_4680), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2404_s_current_state_reg ( .D(
        new_AGEMA_signal_1857), .CK(clk), .Q(new_AGEMA_signal_4682), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2406_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_L2), .CK(clk), .Q(new_AGEMA_signal_4684), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2410_s_current_state_reg ( .D(
        new_AGEMA_signal_1858), .CK(clk), .Q(new_AGEMA_signal_4688), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2414_s_current_state_reg ( .D(
        new_AGEMA_signal_1859), .CK(clk), .Q(new_AGEMA_signal_4692), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2424_s_current_state_reg ( .D(Ciphertext_s0[41]), 
        .CK(clk), .Q(new_AGEMA_signal_4702), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2426_s_current_state_reg ( .D(Ciphertext_s1[41]), 
        .CK(clk), .Q(new_AGEMA_signal_4704), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2428_s_current_state_reg ( .D(Ciphertext_s2[41]), 
        .CK(clk), .Q(new_AGEMA_signal_4706), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2436_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_Q6), .CK(clk), .Q(new_AGEMA_signal_4714), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2438_s_current_state_reg ( .D(
        new_AGEMA_signal_1868), .CK(clk), .Q(new_AGEMA_signal_4716), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2440_s_current_state_reg ( .D(
        new_AGEMA_signal_1869), .CK(clk), .Q(new_AGEMA_signal_4718), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2442_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_L2), .CK(clk), .Q(new_AGEMA_signal_4720), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2446_s_current_state_reg ( .D(
        new_AGEMA_signal_1870), .CK(clk), .Q(new_AGEMA_signal_4724), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2450_s_current_state_reg ( .D(
        new_AGEMA_signal_1871), .CK(clk), .Q(new_AGEMA_signal_4728), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2460_s_current_state_reg ( .D(Ciphertext_s0[45]), 
        .CK(clk), .Q(new_AGEMA_signal_4738), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2462_s_current_state_reg ( .D(Ciphertext_s1[45]), 
        .CK(clk), .Q(new_AGEMA_signal_4740), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2464_s_current_state_reg ( .D(Ciphertext_s2[45]), 
        .CK(clk), .Q(new_AGEMA_signal_4742), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2472_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_Q6), .CK(clk), .Q(new_AGEMA_signal_4750), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2474_s_current_state_reg ( .D(
        new_AGEMA_signal_1880), .CK(clk), .Q(new_AGEMA_signal_4752), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2476_s_current_state_reg ( .D(
        new_AGEMA_signal_1881), .CK(clk), .Q(new_AGEMA_signal_4754), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2478_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_L2), .CK(clk), .Q(new_AGEMA_signal_4756), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2482_s_current_state_reg ( .D(
        new_AGEMA_signal_1882), .CK(clk), .Q(new_AGEMA_signal_4760), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2486_s_current_state_reg ( .D(
        new_AGEMA_signal_1883), .CK(clk), .Q(new_AGEMA_signal_4764), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2496_s_current_state_reg ( .D(Ciphertext_s0[49]), 
        .CK(clk), .Q(new_AGEMA_signal_4774), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2498_s_current_state_reg ( .D(Ciphertext_s1[49]), 
        .CK(clk), .Q(new_AGEMA_signal_4776), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2500_s_current_state_reg ( .D(Ciphertext_s2[49]), 
        .CK(clk), .Q(new_AGEMA_signal_4778), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2508_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_Q6), .CK(clk), .Q(new_AGEMA_signal_4786), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2510_s_current_state_reg ( .D(
        new_AGEMA_signal_1892), .CK(clk), .Q(new_AGEMA_signal_4788), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2512_s_current_state_reg ( .D(
        new_AGEMA_signal_1893), .CK(clk), .Q(new_AGEMA_signal_4790), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2514_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_L2), .CK(clk), .Q(new_AGEMA_signal_4792), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2518_s_current_state_reg ( .D(
        new_AGEMA_signal_1894), .CK(clk), .Q(new_AGEMA_signal_4796), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2522_s_current_state_reg ( .D(
        new_AGEMA_signal_1895), .CK(clk), .Q(new_AGEMA_signal_4800), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2532_s_current_state_reg ( .D(Ciphertext_s0[53]), 
        .CK(clk), .Q(new_AGEMA_signal_4810), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2534_s_current_state_reg ( .D(Ciphertext_s1[53]), 
        .CK(clk), .Q(new_AGEMA_signal_4812), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2536_s_current_state_reg ( .D(Ciphertext_s2[53]), 
        .CK(clk), .Q(new_AGEMA_signal_4814), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2544_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_Q6), .CK(clk), .Q(new_AGEMA_signal_4822), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2546_s_current_state_reg ( .D(
        new_AGEMA_signal_1904), .CK(clk), .Q(new_AGEMA_signal_4824), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2548_s_current_state_reg ( .D(
        new_AGEMA_signal_1905), .CK(clk), .Q(new_AGEMA_signal_4826), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2550_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_L2), .CK(clk), .Q(new_AGEMA_signal_4828), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2554_s_current_state_reg ( .D(
        new_AGEMA_signal_1906), .CK(clk), .Q(new_AGEMA_signal_4832), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2558_s_current_state_reg ( .D(
        new_AGEMA_signal_1907), .CK(clk), .Q(new_AGEMA_signal_4836), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2568_s_current_state_reg ( .D(Ciphertext_s0[57]), 
        .CK(clk), .Q(new_AGEMA_signal_4846), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2570_s_current_state_reg ( .D(Ciphertext_s1[57]), 
        .CK(clk), .Q(new_AGEMA_signal_4848), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2572_s_current_state_reg ( .D(Ciphertext_s2[57]), 
        .CK(clk), .Q(new_AGEMA_signal_4850), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2580_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_Q6), .CK(clk), .Q(new_AGEMA_signal_4858), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2582_s_current_state_reg ( .D(
        new_AGEMA_signal_1916), .CK(clk), .Q(new_AGEMA_signal_4860), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2584_s_current_state_reg ( .D(
        new_AGEMA_signal_1917), .CK(clk), .Q(new_AGEMA_signal_4862), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2586_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_L2), .CK(clk), .Q(new_AGEMA_signal_4864), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2590_s_current_state_reg ( .D(
        new_AGEMA_signal_1918), .CK(clk), .Q(new_AGEMA_signal_4868), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2594_s_current_state_reg ( .D(
        new_AGEMA_signal_1919), .CK(clk), .Q(new_AGEMA_signal_4872), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2604_s_current_state_reg ( .D(Ciphertext_s0[61]), 
        .CK(clk), .Q(new_AGEMA_signal_4882), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2606_s_current_state_reg ( .D(Ciphertext_s1[61]), 
        .CK(clk), .Q(new_AGEMA_signal_4884), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2608_s_current_state_reg ( .D(Ciphertext_s2[61]), 
        .CK(clk), .Q(new_AGEMA_signal_4886), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2616_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_Q6), .CK(clk), .Q(new_AGEMA_signal_4894), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2618_s_current_state_reg ( .D(
        new_AGEMA_signal_1928), .CK(clk), .Q(new_AGEMA_signal_4896), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2620_s_current_state_reg ( .D(
        new_AGEMA_signal_1929), .CK(clk), .Q(new_AGEMA_signal_4898), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2622_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_L2), .CK(clk), .Q(new_AGEMA_signal_4900), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2626_s_current_state_reg ( .D(
        new_AGEMA_signal_1930), .CK(clk), .Q(new_AGEMA_signal_4904), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2630_s_current_state_reg ( .D(
        new_AGEMA_signal_1931), .CK(clk), .Q(new_AGEMA_signal_4908), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2640_s_current_state_reg ( .D(FSMUpdate[1]), 
        .CK(clk), .Q(new_AGEMA_signal_4918), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2644_s_current_state_reg ( .D(FSM_1), .CK(clk), 
        .Q(new_AGEMA_signal_4922), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2648_s_current_state_reg ( .D(FSM[4]), .CK(clk), 
        .Q(new_AGEMA_signal_4926), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2652_s_current_state_reg ( .D(FSM[5]), .CK(clk), 
        .Q(new_AGEMA_signal_4930), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2656_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[0]), .CK(clk), .Q(new_AGEMA_signal_4934), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2660_s_current_state_reg ( .D(
        new_AGEMA_signal_1356), .CK(clk), .Q(new_AGEMA_signal_4938), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2664_s_current_state_reg ( .D(
        new_AGEMA_signal_1357), .CK(clk), .Q(new_AGEMA_signal_4942), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2668_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[1]), .CK(clk), .Q(new_AGEMA_signal_4946), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2672_s_current_state_reg ( .D(
        new_AGEMA_signal_1362), .CK(clk), .Q(new_AGEMA_signal_4950), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2676_s_current_state_reg ( .D(
        new_AGEMA_signal_1363), .CK(clk), .Q(new_AGEMA_signal_4954), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2680_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[4]), .CK(clk), .Q(new_AGEMA_signal_4958), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2684_s_current_state_reg ( .D(
        new_AGEMA_signal_1380), .CK(clk), .Q(new_AGEMA_signal_4962), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2688_s_current_state_reg ( .D(
        new_AGEMA_signal_1381), .CK(clk), .Q(new_AGEMA_signal_4966), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2692_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[5]), .CK(clk), .Q(new_AGEMA_signal_4970), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2696_s_current_state_reg ( .D(
        new_AGEMA_signal_1386), .CK(clk), .Q(new_AGEMA_signal_4974), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2700_s_current_state_reg ( .D(
        new_AGEMA_signal_1387), .CK(clk), .Q(new_AGEMA_signal_4978), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2704_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[8]), .CK(clk), .Q(new_AGEMA_signal_4982), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2708_s_current_state_reg ( .D(
        new_AGEMA_signal_1404), .CK(clk), .Q(new_AGEMA_signal_4986), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2712_s_current_state_reg ( .D(
        new_AGEMA_signal_1405), .CK(clk), .Q(new_AGEMA_signal_4990), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2716_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[9]), .CK(clk), .Q(new_AGEMA_signal_4994), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2720_s_current_state_reg ( .D(
        new_AGEMA_signal_1410), .CK(clk), .Q(new_AGEMA_signal_4998), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2724_s_current_state_reg ( .D(
        new_AGEMA_signal_1411), .CK(clk), .Q(new_AGEMA_signal_5002), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2728_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[12]), .CK(clk), .Q(
        new_AGEMA_signal_5006), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2732_s_current_state_reg ( .D(
        new_AGEMA_signal_1428), .CK(clk), .Q(new_AGEMA_signal_5010), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2736_s_current_state_reg ( .D(
        new_AGEMA_signal_1429), .CK(clk), .Q(new_AGEMA_signal_5014), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2740_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[13]), .CK(clk), .Q(
        new_AGEMA_signal_5018), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2744_s_current_state_reg ( .D(
        new_AGEMA_signal_1434), .CK(clk), .Q(new_AGEMA_signal_5022), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2748_s_current_state_reg ( .D(
        new_AGEMA_signal_1435), .CK(clk), .Q(new_AGEMA_signal_5026), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2752_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[16]), .CK(clk), .Q(
        new_AGEMA_signal_5030), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2756_s_current_state_reg ( .D(
        new_AGEMA_signal_1452), .CK(clk), .Q(new_AGEMA_signal_5034), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2760_s_current_state_reg ( .D(
        new_AGEMA_signal_1453), .CK(clk), .Q(new_AGEMA_signal_5038), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2764_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[17]), .CK(clk), .Q(
        new_AGEMA_signal_5042), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2768_s_current_state_reg ( .D(
        new_AGEMA_signal_1458), .CK(clk), .Q(new_AGEMA_signal_5046), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2772_s_current_state_reg ( .D(
        new_AGEMA_signal_1459), .CK(clk), .Q(new_AGEMA_signal_5050), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2776_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[20]), .CK(clk), .Q(
        new_AGEMA_signal_5054), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2780_s_current_state_reg ( .D(
        new_AGEMA_signal_1476), .CK(clk), .Q(new_AGEMA_signal_5058), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2784_s_current_state_reg ( .D(
        new_AGEMA_signal_1477), .CK(clk), .Q(new_AGEMA_signal_5062), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2788_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[21]), .CK(clk), .Q(
        new_AGEMA_signal_5066), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2792_s_current_state_reg ( .D(
        new_AGEMA_signal_1482), .CK(clk), .Q(new_AGEMA_signal_5070), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2796_s_current_state_reg ( .D(
        new_AGEMA_signal_1483), .CK(clk), .Q(new_AGEMA_signal_5074), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2800_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[24]), .CK(clk), .Q(
        new_AGEMA_signal_5078), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2804_s_current_state_reg ( .D(
        new_AGEMA_signal_1500), .CK(clk), .Q(new_AGEMA_signal_5082), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2808_s_current_state_reg ( .D(
        new_AGEMA_signal_1501), .CK(clk), .Q(new_AGEMA_signal_5086), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2812_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[25]), .CK(clk), .Q(
        new_AGEMA_signal_5090), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2816_s_current_state_reg ( .D(
        new_AGEMA_signal_1506), .CK(clk), .Q(new_AGEMA_signal_5094), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2820_s_current_state_reg ( .D(
        new_AGEMA_signal_1507), .CK(clk), .Q(new_AGEMA_signal_5098), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2824_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[28]), .CK(clk), .Q(
        new_AGEMA_signal_5102), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2828_s_current_state_reg ( .D(
        new_AGEMA_signal_1524), .CK(clk), .Q(new_AGEMA_signal_5106), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2832_s_current_state_reg ( .D(
        new_AGEMA_signal_1525), .CK(clk), .Q(new_AGEMA_signal_5110), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2836_s_current_state_reg ( .D(
        TweakeyGeneration_key_Feedback[29]), .CK(clk), .Q(
        new_AGEMA_signal_5114), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2840_s_current_state_reg ( .D(
        new_AGEMA_signal_1530), .CK(clk), .Q(new_AGEMA_signal_5118), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2844_s_current_state_reg ( .D(
        new_AGEMA_signal_1531), .CK(clk), .Q(new_AGEMA_signal_5122), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3040_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[63]), .CK(clk), .Q(
        new_AGEMA_signal_5318), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3044_s_current_state_reg ( .D(
        new_AGEMA_signal_1738), .CK(clk), .Q(new_AGEMA_signal_5322), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3048_s_current_state_reg ( .D(
        new_AGEMA_signal_1739), .CK(clk), .Q(new_AGEMA_signal_5326), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3052_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[62]), .CK(clk), .Q(
        new_AGEMA_signal_5330), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3056_s_current_state_reg ( .D(
        new_AGEMA_signal_1732), .CK(clk), .Q(new_AGEMA_signal_5334), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3060_s_current_state_reg ( .D(
        new_AGEMA_signal_1733), .CK(clk), .Q(new_AGEMA_signal_5338), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3064_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[61]), .CK(clk), .Q(
        new_AGEMA_signal_5342), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3068_s_current_state_reg ( .D(
        new_AGEMA_signal_1726), .CK(clk), .Q(new_AGEMA_signal_5346), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3072_s_current_state_reg ( .D(
        new_AGEMA_signal_1727), .CK(clk), .Q(new_AGEMA_signal_5350), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3076_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[60]), .CK(clk), .Q(
        new_AGEMA_signal_5354), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3080_s_current_state_reg ( .D(
        new_AGEMA_signal_1720), .CK(clk), .Q(new_AGEMA_signal_5358), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3084_s_current_state_reg ( .D(
        new_AGEMA_signal_1721), .CK(clk), .Q(new_AGEMA_signal_5362), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3088_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[59]), .CK(clk), .Q(
        new_AGEMA_signal_5366), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3092_s_current_state_reg ( .D(
        new_AGEMA_signal_1714), .CK(clk), .Q(new_AGEMA_signal_5370), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3096_s_current_state_reg ( .D(
        new_AGEMA_signal_1715), .CK(clk), .Q(new_AGEMA_signal_5374), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3100_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[58]), .CK(clk), .Q(
        new_AGEMA_signal_5378), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3104_s_current_state_reg ( .D(
        new_AGEMA_signal_1708), .CK(clk), .Q(new_AGEMA_signal_5382), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3108_s_current_state_reg ( .D(
        new_AGEMA_signal_1709), .CK(clk), .Q(new_AGEMA_signal_5386), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3112_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[57]), .CK(clk), .Q(
        new_AGEMA_signal_5390), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3116_s_current_state_reg ( .D(
        new_AGEMA_signal_1702), .CK(clk), .Q(new_AGEMA_signal_5394), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3120_s_current_state_reg ( .D(
        new_AGEMA_signal_1703), .CK(clk), .Q(new_AGEMA_signal_5398), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3124_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[56]), .CK(clk), .Q(
        new_AGEMA_signal_5402), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3128_s_current_state_reg ( .D(
        new_AGEMA_signal_1696), .CK(clk), .Q(new_AGEMA_signal_5406), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3132_s_current_state_reg ( .D(
        new_AGEMA_signal_1697), .CK(clk), .Q(new_AGEMA_signal_5410), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3136_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[55]), .CK(clk), .Q(
        new_AGEMA_signal_5414), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3140_s_current_state_reg ( .D(
        new_AGEMA_signal_1690), .CK(clk), .Q(new_AGEMA_signal_5418), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3144_s_current_state_reg ( .D(
        new_AGEMA_signal_1691), .CK(clk), .Q(new_AGEMA_signal_5422), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3148_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[54]), .CK(clk), .Q(
        new_AGEMA_signal_5426), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3152_s_current_state_reg ( .D(
        new_AGEMA_signal_1684), .CK(clk), .Q(new_AGEMA_signal_5430), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3156_s_current_state_reg ( .D(
        new_AGEMA_signal_1685), .CK(clk), .Q(new_AGEMA_signal_5434), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3160_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[53]), .CK(clk), .Q(
        new_AGEMA_signal_5438), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3164_s_current_state_reg ( .D(
        new_AGEMA_signal_1678), .CK(clk), .Q(new_AGEMA_signal_5442), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3168_s_current_state_reg ( .D(
        new_AGEMA_signal_1679), .CK(clk), .Q(new_AGEMA_signal_5446), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3172_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[52]), .CK(clk), .Q(
        new_AGEMA_signal_5450), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3176_s_current_state_reg ( .D(
        new_AGEMA_signal_1672), .CK(clk), .Q(new_AGEMA_signal_5454), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3180_s_current_state_reg ( .D(
        new_AGEMA_signal_1673), .CK(clk), .Q(new_AGEMA_signal_5458), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3184_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[51]), .CK(clk), .Q(
        new_AGEMA_signal_5462), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3188_s_current_state_reg ( .D(
        new_AGEMA_signal_1666), .CK(clk), .Q(new_AGEMA_signal_5466), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3192_s_current_state_reg ( .D(
        new_AGEMA_signal_1667), .CK(clk), .Q(new_AGEMA_signal_5470), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3196_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[50]), .CK(clk), .Q(
        new_AGEMA_signal_5474), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3200_s_current_state_reg ( .D(
        new_AGEMA_signal_1660), .CK(clk), .Q(new_AGEMA_signal_5478), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3204_s_current_state_reg ( .D(
        new_AGEMA_signal_1661), .CK(clk), .Q(new_AGEMA_signal_5482), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3208_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[49]), .CK(clk), .Q(
        new_AGEMA_signal_5486), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3212_s_current_state_reg ( .D(
        new_AGEMA_signal_1654), .CK(clk), .Q(new_AGEMA_signal_5490), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3216_s_current_state_reg ( .D(
        new_AGEMA_signal_1655), .CK(clk), .Q(new_AGEMA_signal_5494), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3220_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[48]), .CK(clk), .Q(
        new_AGEMA_signal_5498), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3224_s_current_state_reg ( .D(
        new_AGEMA_signal_1648), .CK(clk), .Q(new_AGEMA_signal_5502), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3228_s_current_state_reg ( .D(
        new_AGEMA_signal_1649), .CK(clk), .Q(new_AGEMA_signal_5506), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3232_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[47]), .CK(clk), .Q(
        new_AGEMA_signal_5510), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3236_s_current_state_reg ( .D(
        new_AGEMA_signal_1642), .CK(clk), .Q(new_AGEMA_signal_5514), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3240_s_current_state_reg ( .D(
        new_AGEMA_signal_1643), .CK(clk), .Q(new_AGEMA_signal_5518), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3244_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[46]), .CK(clk), .Q(
        new_AGEMA_signal_5522), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3248_s_current_state_reg ( .D(
        new_AGEMA_signal_1636), .CK(clk), .Q(new_AGEMA_signal_5526), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3252_s_current_state_reg ( .D(
        new_AGEMA_signal_1637), .CK(clk), .Q(new_AGEMA_signal_5530), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3256_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[45]), .CK(clk), .Q(
        new_AGEMA_signal_5534), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3260_s_current_state_reg ( .D(
        new_AGEMA_signal_1630), .CK(clk), .Q(new_AGEMA_signal_5538), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3264_s_current_state_reg ( .D(
        new_AGEMA_signal_1631), .CK(clk), .Q(new_AGEMA_signal_5542), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3268_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[44]), .CK(clk), .Q(
        new_AGEMA_signal_5546), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3272_s_current_state_reg ( .D(
        new_AGEMA_signal_1624), .CK(clk), .Q(new_AGEMA_signal_5550), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3276_s_current_state_reg ( .D(
        new_AGEMA_signal_1625), .CK(clk), .Q(new_AGEMA_signal_5554), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3280_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[43]), .CK(clk), .Q(
        new_AGEMA_signal_5558), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3284_s_current_state_reg ( .D(
        new_AGEMA_signal_1618), .CK(clk), .Q(new_AGEMA_signal_5562), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3288_s_current_state_reg ( .D(
        new_AGEMA_signal_1619), .CK(clk), .Q(new_AGEMA_signal_5566), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3292_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[42]), .CK(clk), .Q(
        new_AGEMA_signal_5570), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3296_s_current_state_reg ( .D(
        new_AGEMA_signal_1612), .CK(clk), .Q(new_AGEMA_signal_5574), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3300_s_current_state_reg ( .D(
        new_AGEMA_signal_1613), .CK(clk), .Q(new_AGEMA_signal_5578), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3304_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[41]), .CK(clk), .Q(
        new_AGEMA_signal_5582), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3308_s_current_state_reg ( .D(
        new_AGEMA_signal_1606), .CK(clk), .Q(new_AGEMA_signal_5586), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3312_s_current_state_reg ( .D(
        new_AGEMA_signal_1607), .CK(clk), .Q(new_AGEMA_signal_5590), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3316_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[40]), .CK(clk), .Q(
        new_AGEMA_signal_5594), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3320_s_current_state_reg ( .D(
        new_AGEMA_signal_1600), .CK(clk), .Q(new_AGEMA_signal_5598), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3324_s_current_state_reg ( .D(
        new_AGEMA_signal_1601), .CK(clk), .Q(new_AGEMA_signal_5602), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3328_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[39]), .CK(clk), .Q(
        new_AGEMA_signal_5606), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3332_s_current_state_reg ( .D(
        new_AGEMA_signal_1594), .CK(clk), .Q(new_AGEMA_signal_5610), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3336_s_current_state_reg ( .D(
        new_AGEMA_signal_1595), .CK(clk), .Q(new_AGEMA_signal_5614), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3340_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[38]), .CK(clk), .Q(
        new_AGEMA_signal_5618), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3344_s_current_state_reg ( .D(
        new_AGEMA_signal_1588), .CK(clk), .Q(new_AGEMA_signal_5622), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3348_s_current_state_reg ( .D(
        new_AGEMA_signal_1589), .CK(clk), .Q(new_AGEMA_signal_5626), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3352_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[37]), .CK(clk), .Q(
        new_AGEMA_signal_5630), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3356_s_current_state_reg ( .D(
        new_AGEMA_signal_1582), .CK(clk), .Q(new_AGEMA_signal_5634), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3360_s_current_state_reg ( .D(
        new_AGEMA_signal_1583), .CK(clk), .Q(new_AGEMA_signal_5638), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3364_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[36]), .CK(clk), .Q(
        new_AGEMA_signal_5642), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3368_s_current_state_reg ( .D(
        new_AGEMA_signal_1576), .CK(clk), .Q(new_AGEMA_signal_5646), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3372_s_current_state_reg ( .D(
        new_AGEMA_signal_1577), .CK(clk), .Q(new_AGEMA_signal_5650), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3376_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[35]), .CK(clk), .Q(
        new_AGEMA_signal_5654), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3380_s_current_state_reg ( .D(
        new_AGEMA_signal_1570), .CK(clk), .Q(new_AGEMA_signal_5658), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3384_s_current_state_reg ( .D(
        new_AGEMA_signal_1571), .CK(clk), .Q(new_AGEMA_signal_5662), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3388_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[34]), .CK(clk), .Q(
        new_AGEMA_signal_5666), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3392_s_current_state_reg ( .D(
        new_AGEMA_signal_1564), .CK(clk), .Q(new_AGEMA_signal_5670), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3396_s_current_state_reg ( .D(
        new_AGEMA_signal_1565), .CK(clk), .Q(new_AGEMA_signal_5674), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3400_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[33]), .CK(clk), .Q(
        new_AGEMA_signal_5678), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3404_s_current_state_reg ( .D(
        new_AGEMA_signal_1558), .CK(clk), .Q(new_AGEMA_signal_5682), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3408_s_current_state_reg ( .D(
        new_AGEMA_signal_1559), .CK(clk), .Q(new_AGEMA_signal_5686), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3412_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[32]), .CK(clk), .Q(
        new_AGEMA_signal_5690), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3416_s_current_state_reg ( .D(
        new_AGEMA_signal_1552), .CK(clk), .Q(new_AGEMA_signal_5694), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3420_s_current_state_reg ( .D(
        new_AGEMA_signal_1553), .CK(clk), .Q(new_AGEMA_signal_5698), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3424_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[31]), .CK(clk), .Q(
        new_AGEMA_signal_5702), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3428_s_current_state_reg ( .D(
        new_AGEMA_signal_1546), .CK(clk), .Q(new_AGEMA_signal_5706), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3432_s_current_state_reg ( .D(
        new_AGEMA_signal_1547), .CK(clk), .Q(new_AGEMA_signal_5710), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3436_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[30]), .CK(clk), .Q(
        new_AGEMA_signal_5714), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3440_s_current_state_reg ( .D(
        new_AGEMA_signal_1540), .CK(clk), .Q(new_AGEMA_signal_5718), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3444_s_current_state_reg ( .D(
        new_AGEMA_signal_1541), .CK(clk), .Q(new_AGEMA_signal_5722), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3448_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[29]), .CK(clk), .Q(
        new_AGEMA_signal_5726), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3452_s_current_state_reg ( .D(
        new_AGEMA_signal_1534), .CK(clk), .Q(new_AGEMA_signal_5730), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3456_s_current_state_reg ( .D(
        new_AGEMA_signal_1535), .CK(clk), .Q(new_AGEMA_signal_5734), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3460_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[28]), .CK(clk), .Q(
        new_AGEMA_signal_5738), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3464_s_current_state_reg ( .D(
        new_AGEMA_signal_1528), .CK(clk), .Q(new_AGEMA_signal_5742), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3468_s_current_state_reg ( .D(
        new_AGEMA_signal_1529), .CK(clk), .Q(new_AGEMA_signal_5746), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3472_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[27]), .CK(clk), .Q(
        new_AGEMA_signal_5750), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3476_s_current_state_reg ( .D(
        new_AGEMA_signal_1522), .CK(clk), .Q(new_AGEMA_signal_5754), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3480_s_current_state_reg ( .D(
        new_AGEMA_signal_1523), .CK(clk), .Q(new_AGEMA_signal_5758), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3484_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[26]), .CK(clk), .Q(
        new_AGEMA_signal_5762), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3488_s_current_state_reg ( .D(
        new_AGEMA_signal_1516), .CK(clk), .Q(new_AGEMA_signal_5766), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3492_s_current_state_reg ( .D(
        new_AGEMA_signal_1517), .CK(clk), .Q(new_AGEMA_signal_5770), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3496_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[25]), .CK(clk), .Q(
        new_AGEMA_signal_5774), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3500_s_current_state_reg ( .D(
        new_AGEMA_signal_1510), .CK(clk), .Q(new_AGEMA_signal_5778), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3504_s_current_state_reg ( .D(
        new_AGEMA_signal_1511), .CK(clk), .Q(new_AGEMA_signal_5782), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3508_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[24]), .CK(clk), .Q(
        new_AGEMA_signal_5786), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3512_s_current_state_reg ( .D(
        new_AGEMA_signal_1504), .CK(clk), .Q(new_AGEMA_signal_5790), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3516_s_current_state_reg ( .D(
        new_AGEMA_signal_1505), .CK(clk), .Q(new_AGEMA_signal_5794), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3520_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[23]), .CK(clk), .Q(
        new_AGEMA_signal_5798), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3524_s_current_state_reg ( .D(
        new_AGEMA_signal_1498), .CK(clk), .Q(new_AGEMA_signal_5802), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3528_s_current_state_reg ( .D(
        new_AGEMA_signal_1499), .CK(clk), .Q(new_AGEMA_signal_5806), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3532_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[22]), .CK(clk), .Q(
        new_AGEMA_signal_5810), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3536_s_current_state_reg ( .D(
        new_AGEMA_signal_1492), .CK(clk), .Q(new_AGEMA_signal_5814), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3540_s_current_state_reg ( .D(
        new_AGEMA_signal_1493), .CK(clk), .Q(new_AGEMA_signal_5818), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3544_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[21]), .CK(clk), .Q(
        new_AGEMA_signal_5822), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3548_s_current_state_reg ( .D(
        new_AGEMA_signal_1486), .CK(clk), .Q(new_AGEMA_signal_5826), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3552_s_current_state_reg ( .D(
        new_AGEMA_signal_1487), .CK(clk), .Q(new_AGEMA_signal_5830), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3556_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[20]), .CK(clk), .Q(
        new_AGEMA_signal_5834), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3560_s_current_state_reg ( .D(
        new_AGEMA_signal_1480), .CK(clk), .Q(new_AGEMA_signal_5838), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3564_s_current_state_reg ( .D(
        new_AGEMA_signal_1481), .CK(clk), .Q(new_AGEMA_signal_5842), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3568_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[19]), .CK(clk), .Q(
        new_AGEMA_signal_5846), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3572_s_current_state_reg ( .D(
        new_AGEMA_signal_1474), .CK(clk), .Q(new_AGEMA_signal_5850), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3576_s_current_state_reg ( .D(
        new_AGEMA_signal_1475), .CK(clk), .Q(new_AGEMA_signal_5854), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3580_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[18]), .CK(clk), .Q(
        new_AGEMA_signal_5858), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3584_s_current_state_reg ( .D(
        new_AGEMA_signal_1468), .CK(clk), .Q(new_AGEMA_signal_5862), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3588_s_current_state_reg ( .D(
        new_AGEMA_signal_1469), .CK(clk), .Q(new_AGEMA_signal_5866), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3592_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[17]), .CK(clk), .Q(
        new_AGEMA_signal_5870), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3596_s_current_state_reg ( .D(
        new_AGEMA_signal_1462), .CK(clk), .Q(new_AGEMA_signal_5874), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3600_s_current_state_reg ( .D(
        new_AGEMA_signal_1463), .CK(clk), .Q(new_AGEMA_signal_5878), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3604_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[16]), .CK(clk), .Q(
        new_AGEMA_signal_5882), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3608_s_current_state_reg ( .D(
        new_AGEMA_signal_1456), .CK(clk), .Q(new_AGEMA_signal_5886), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3612_s_current_state_reg ( .D(
        new_AGEMA_signal_1457), .CK(clk), .Q(new_AGEMA_signal_5890), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3616_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[15]), .CK(clk), .Q(
        new_AGEMA_signal_5894), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3620_s_current_state_reg ( .D(
        new_AGEMA_signal_1450), .CK(clk), .Q(new_AGEMA_signal_5898), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3624_s_current_state_reg ( .D(
        new_AGEMA_signal_1451), .CK(clk), .Q(new_AGEMA_signal_5902), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3628_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[14]), .CK(clk), .Q(
        new_AGEMA_signal_5906), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3632_s_current_state_reg ( .D(
        new_AGEMA_signal_1444), .CK(clk), .Q(new_AGEMA_signal_5910), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3636_s_current_state_reg ( .D(
        new_AGEMA_signal_1445), .CK(clk), .Q(new_AGEMA_signal_5914), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3640_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[13]), .CK(clk), .Q(
        new_AGEMA_signal_5918), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3644_s_current_state_reg ( .D(
        new_AGEMA_signal_1438), .CK(clk), .Q(new_AGEMA_signal_5922), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3648_s_current_state_reg ( .D(
        new_AGEMA_signal_1439), .CK(clk), .Q(new_AGEMA_signal_5926), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3652_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[12]), .CK(clk), .Q(
        new_AGEMA_signal_5930), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3656_s_current_state_reg ( .D(
        new_AGEMA_signal_1432), .CK(clk), .Q(new_AGEMA_signal_5934), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3660_s_current_state_reg ( .D(
        new_AGEMA_signal_1433), .CK(clk), .Q(new_AGEMA_signal_5938), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3664_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[11]), .CK(clk), .Q(
        new_AGEMA_signal_5942), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3668_s_current_state_reg ( .D(
        new_AGEMA_signal_1426), .CK(clk), .Q(new_AGEMA_signal_5946), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3672_s_current_state_reg ( .D(
        new_AGEMA_signal_1427), .CK(clk), .Q(new_AGEMA_signal_5950), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3676_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[10]), .CK(clk), .Q(
        new_AGEMA_signal_5954), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3680_s_current_state_reg ( .D(
        new_AGEMA_signal_1420), .CK(clk), .Q(new_AGEMA_signal_5958), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3684_s_current_state_reg ( .D(
        new_AGEMA_signal_1421), .CK(clk), .Q(new_AGEMA_signal_5962), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3688_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[9]), .CK(clk), .Q(
        new_AGEMA_signal_5966), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3692_s_current_state_reg ( .D(
        new_AGEMA_signal_1414), .CK(clk), .Q(new_AGEMA_signal_5970), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3696_s_current_state_reg ( .D(
        new_AGEMA_signal_1415), .CK(clk), .Q(new_AGEMA_signal_5974), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3700_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[8]), .CK(clk), .Q(
        new_AGEMA_signal_5978), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3704_s_current_state_reg ( .D(
        new_AGEMA_signal_1408), .CK(clk), .Q(new_AGEMA_signal_5982), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3708_s_current_state_reg ( .D(
        new_AGEMA_signal_1409), .CK(clk), .Q(new_AGEMA_signal_5986), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3712_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[7]), .CK(clk), .Q(
        new_AGEMA_signal_5990), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3716_s_current_state_reg ( .D(
        new_AGEMA_signal_1402), .CK(clk), .Q(new_AGEMA_signal_5994), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3720_s_current_state_reg ( .D(
        new_AGEMA_signal_1403), .CK(clk), .Q(new_AGEMA_signal_5998), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3724_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[6]), .CK(clk), .Q(
        new_AGEMA_signal_6002), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3728_s_current_state_reg ( .D(
        new_AGEMA_signal_1396), .CK(clk), .Q(new_AGEMA_signal_6006), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3732_s_current_state_reg ( .D(
        new_AGEMA_signal_1397), .CK(clk), .Q(new_AGEMA_signal_6010), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3736_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[5]), .CK(clk), .Q(
        new_AGEMA_signal_6014), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3740_s_current_state_reg ( .D(
        new_AGEMA_signal_1390), .CK(clk), .Q(new_AGEMA_signal_6018), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3744_s_current_state_reg ( .D(
        new_AGEMA_signal_1391), .CK(clk), .Q(new_AGEMA_signal_6022), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3748_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[4]), .CK(clk), .Q(
        new_AGEMA_signal_6026), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3752_s_current_state_reg ( .D(
        new_AGEMA_signal_1384), .CK(clk), .Q(new_AGEMA_signal_6030), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3756_s_current_state_reg ( .D(
        new_AGEMA_signal_1385), .CK(clk), .Q(new_AGEMA_signal_6034), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3760_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[3]), .CK(clk), .Q(
        new_AGEMA_signal_6038), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3764_s_current_state_reg ( .D(
        new_AGEMA_signal_1378), .CK(clk), .Q(new_AGEMA_signal_6042), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3768_s_current_state_reg ( .D(
        new_AGEMA_signal_1379), .CK(clk), .Q(new_AGEMA_signal_6046), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3772_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[2]), .CK(clk), .Q(
        new_AGEMA_signal_6050), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3776_s_current_state_reg ( .D(
        new_AGEMA_signal_1372), .CK(clk), .Q(new_AGEMA_signal_6054), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3780_s_current_state_reg ( .D(
        new_AGEMA_signal_1373), .CK(clk), .Q(new_AGEMA_signal_6058), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3784_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[1]), .CK(clk), .Q(
        new_AGEMA_signal_6062), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3788_s_current_state_reg ( .D(
        new_AGEMA_signal_1366), .CK(clk), .Q(new_AGEMA_signal_6066), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3792_s_current_state_reg ( .D(
        new_AGEMA_signal_1367), .CK(clk), .Q(new_AGEMA_signal_6070), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3796_s_current_state_reg ( .D(
        TweakeyGeneration_StateRegInput[0]), .CK(clk), .Q(
        new_AGEMA_signal_6074), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3800_s_current_state_reg ( .D(
        new_AGEMA_signal_1360), .CK(clk), .Q(new_AGEMA_signal_6078), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3804_s_current_state_reg ( .D(
        new_AGEMA_signal_1361), .CK(clk), .Q(new_AGEMA_signal_6082), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3808_s_current_state_reg ( .D(FSMSelected[5]), 
        .CK(clk), .Q(new_AGEMA_signal_6086), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3812_s_current_state_reg ( .D(FSMSelected[4]), 
        .CK(clk), .Q(new_AGEMA_signal_6090), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3816_s_current_state_reg ( .D(FSMSelected[3]), 
        .CK(clk), .Q(new_AGEMA_signal_6094), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3820_s_current_state_reg ( .D(FSMSelected[2]), 
        .CK(clk), .Q(new_AGEMA_signal_6098), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3824_s_current_state_reg ( .D(FSMSelected[1]), 
        .CK(clk), .Q(new_AGEMA_signal_6102), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3828_s_current_state_reg ( .D(FSMSelected[0]), 
        .CK(clk), .Q(new_AGEMA_signal_6106), .QN() );
  MUX2_X1 PlaintextMUX_MUXInst_2_U1_Ins_0_U1 ( .A(MCOutput[2]), .B(
        new_AGEMA_signal_3281), .S(new_AGEMA_signal_3279), .Z(StateRegInput[2]) );
  MUX2_X1 PlaintextMUX_MUXInst_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2666), .B(
        new_AGEMA_signal_3283), .S(new_AGEMA_signal_3279), .Z(
        new_AGEMA_signal_2680) );
  MUX2_X1 PlaintextMUX_MUXInst_2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2667), .B(
        new_AGEMA_signal_3285), .S(new_AGEMA_signal_3279), .Z(
        new_AGEMA_signal_2681) );
  MUX2_X1 PlaintextMUX_MUXInst_3_U1_Ins_0_U1 ( .A(MCOutput[3]), .B(
        new_AGEMA_signal_3287), .S(new_AGEMA_signal_3279), .Z(StateRegInput[3]) );
  MUX2_X1 PlaintextMUX_MUXInst_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2786), .B(
        new_AGEMA_signal_3289), .S(new_AGEMA_signal_3279), .Z(
        new_AGEMA_signal_2800) );
  MUX2_X1 PlaintextMUX_MUXInst_3_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2787), .B(
        new_AGEMA_signal_3291), .S(new_AGEMA_signal_3279), .Z(
        new_AGEMA_signal_2801) );
  MUX2_X1 PlaintextMUX_MUXInst_6_U1_Ins_0_U1 ( .A(MCOutput[6]), .B(
        new_AGEMA_signal_3293), .S(new_AGEMA_signal_3279), .Z(StateRegInput[6]) );
  MUX2_X1 PlaintextMUX_MUXInst_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2670), .B(
        new_AGEMA_signal_3295), .S(new_AGEMA_signal_3279), .Z(
        new_AGEMA_signal_2684) );
  MUX2_X1 PlaintextMUX_MUXInst_6_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2671), .B(
        new_AGEMA_signal_3297), .S(new_AGEMA_signal_3279), .Z(
        new_AGEMA_signal_2685) );
  MUX2_X1 PlaintextMUX_MUXInst_7_U1_Ins_0_U1 ( .A(MCOutput[7]), .B(
        new_AGEMA_signal_3299), .S(n46), .Z(StateRegInput[7]) );
  MUX2_X1 PlaintextMUX_MUXInst_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2790), .B(
        new_AGEMA_signal_3301), .S(n46), .Z(new_AGEMA_signal_2804) );
  MUX2_X1 PlaintextMUX_MUXInst_7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2791), .B(
        new_AGEMA_signal_3303), .S(n46), .Z(new_AGEMA_signal_2805) );
  MUX2_X1 PlaintextMUX_MUXInst_10_U1_Ins_0_U1 ( .A(MCOutput[10]), .B(
        new_AGEMA_signal_3305), .S(n47), .Z(StateRegInput[10]) );
  MUX2_X1 PlaintextMUX_MUXInst_10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2674), .B(
        new_AGEMA_signal_3307), .S(n47), .Z(new_AGEMA_signal_2688) );
  MUX2_X1 PlaintextMUX_MUXInst_10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2675), .B(
        new_AGEMA_signal_3309), .S(n47), .Z(new_AGEMA_signal_2689) );
  MUX2_X1 PlaintextMUX_MUXInst_11_U1_Ins_0_U1 ( .A(MCOutput[11]), .B(
        new_AGEMA_signal_3311), .S(n47), .Z(StateRegInput[11]) );
  MUX2_X1 PlaintextMUX_MUXInst_11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2794), .B(
        new_AGEMA_signal_3313), .S(n47), .Z(new_AGEMA_signal_2808) );
  MUX2_X1 PlaintextMUX_MUXInst_11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2795), .B(
        new_AGEMA_signal_3315), .S(n47), .Z(new_AGEMA_signal_2809) );
  MUX2_X1 PlaintextMUX_MUXInst_14_U1_Ins_0_U1 ( .A(MCOutput[14]), .B(
        new_AGEMA_signal_3317), .S(n47), .Z(StateRegInput[14]) );
  MUX2_X1 PlaintextMUX_MUXInst_14_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2902), .B(
        new_AGEMA_signal_3319), .S(n47), .Z(new_AGEMA_signal_2920) );
  MUX2_X1 PlaintextMUX_MUXInst_14_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2903), .B(
        new_AGEMA_signal_3321), .S(n47), .Z(new_AGEMA_signal_2921) );
  MUX2_X1 PlaintextMUX_MUXInst_15_U1_Ins_0_U1 ( .A(MCOutput[15]), .B(
        new_AGEMA_signal_3323), .S(n47), .Z(StateRegInput[15]) );
  MUX2_X1 PlaintextMUX_MUXInst_15_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2990), .B(
        new_AGEMA_signal_3325), .S(n47), .Z(new_AGEMA_signal_3006) );
  MUX2_X1 PlaintextMUX_MUXInst_15_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2991), .B(
        new_AGEMA_signal_3327), .S(n47), .Z(new_AGEMA_signal_3007) );
  MUX2_X1 PlaintextMUX_MUXInst_18_U1_Ins_0_U1 ( .A(MCOutput[18]), .B(
        new_AGEMA_signal_3329), .S(n47), .Z(StateRegInput[18]) );
  MUX2_X1 PlaintextMUX_MUXInst_18_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2654), .B(
        new_AGEMA_signal_3331), .S(n47), .Z(new_AGEMA_signal_2692) );
  MUX2_X1 PlaintextMUX_MUXInst_18_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2655), .B(
        new_AGEMA_signal_3333), .S(n47), .Z(new_AGEMA_signal_2693) );
  MUX2_X1 PlaintextMUX_MUXInst_19_U1_Ins_0_U1 ( .A(MCOutput[19]), .B(
        new_AGEMA_signal_3335), .S(n47), .Z(StateRegInput[19]) );
  MUX2_X1 PlaintextMUX_MUXInst_19_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2772), .B(
        new_AGEMA_signal_3337), .S(n47), .Z(new_AGEMA_signal_2812) );
  MUX2_X1 PlaintextMUX_MUXInst_19_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2773), .B(
        new_AGEMA_signal_3339), .S(n47), .Z(new_AGEMA_signal_2813) );
  MUX2_X1 PlaintextMUX_MUXInst_22_U1_Ins_0_U1 ( .A(MCOutput[22]), .B(
        new_AGEMA_signal_3341), .S(n47), .Z(StateRegInput[22]) );
  MUX2_X1 PlaintextMUX_MUXInst_22_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2658), .B(
        new_AGEMA_signal_3343), .S(n47), .Z(new_AGEMA_signal_2696) );
  MUX2_X1 PlaintextMUX_MUXInst_22_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2659), .B(
        new_AGEMA_signal_3345), .S(n47), .Z(new_AGEMA_signal_2697) );
  MUX2_X1 PlaintextMUX_MUXInst_23_U1_Ins_0_U1 ( .A(MCOutput[23]), .B(
        new_AGEMA_signal_3347), .S(n47), .Z(StateRegInput[23]) );
  MUX2_X1 PlaintextMUX_MUXInst_23_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2776), .B(
        new_AGEMA_signal_3349), .S(n47), .Z(new_AGEMA_signal_2816) );
  MUX2_X1 PlaintextMUX_MUXInst_23_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2777), .B(
        new_AGEMA_signal_3351), .S(n47), .Z(new_AGEMA_signal_2817) );
  MUX2_X1 PlaintextMUX_MUXInst_26_U1_Ins_0_U1 ( .A(MCOutput[26]), .B(
        new_AGEMA_signal_3353), .S(n47), .Z(StateRegInput[26]) );
  MUX2_X1 PlaintextMUX_MUXInst_26_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2882), .B(
        new_AGEMA_signal_3355), .S(n47), .Z(new_AGEMA_signal_2932) );
  MUX2_X1 PlaintextMUX_MUXInst_26_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2883), .B(
        new_AGEMA_signal_3357), .S(n47), .Z(new_AGEMA_signal_2933) );
  MUX2_X1 PlaintextMUX_MUXInst_27_U1_Ins_0_U1 ( .A(MCOutput[27]), .B(
        new_AGEMA_signal_3359), .S(n47), .Z(StateRegInput[27]) );
  MUX2_X1 PlaintextMUX_MUXInst_27_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2978), .B(
        new_AGEMA_signal_3361), .S(n47), .Z(new_AGEMA_signal_3018) );
  MUX2_X1 PlaintextMUX_MUXInst_27_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2979), .B(
        new_AGEMA_signal_3363), .S(n47), .Z(new_AGEMA_signal_3019) );
  MUX2_X1 PlaintextMUX_MUXInst_30_U1_Ins_0_U1 ( .A(MCOutput[30]), .B(
        new_AGEMA_signal_3365), .S(n46), .Z(StateRegInput[30]) );
  MUX2_X1 PlaintextMUX_MUXInst_30_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2662), .B(
        new_AGEMA_signal_3367), .S(n46), .Z(new_AGEMA_signal_2700) );
  MUX2_X1 PlaintextMUX_MUXInst_30_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2663), .B(
        new_AGEMA_signal_3369), .S(n46), .Z(new_AGEMA_signal_2701) );
  MUX2_X1 PlaintextMUX_MUXInst_31_U1_Ins_0_U1 ( .A(MCOutput[31]), .B(
        new_AGEMA_signal_3371), .S(n46), .Z(StateRegInput[31]) );
  MUX2_X1 PlaintextMUX_MUXInst_31_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2782), .B(
        new_AGEMA_signal_3373), .S(n46), .Z(new_AGEMA_signal_2820) );
  MUX2_X1 PlaintextMUX_MUXInst_31_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2783), .B(
        new_AGEMA_signal_3375), .S(n46), .Z(new_AGEMA_signal_2821) );
  MUX2_X1 PlaintextMUX_MUXInst_34_U1_Ins_0_U1 ( .A(MCOutput[34]), .B(
        new_AGEMA_signal_3377), .S(n46), .Z(StateRegInput[34]) );
  MUX2_X1 PlaintextMUX_MUXInst_34_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2456), .B(
        new_AGEMA_signal_3379), .S(n46), .Z(new_AGEMA_signal_2478) );
  MUX2_X1 PlaintextMUX_MUXInst_34_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2457), .B(
        new_AGEMA_signal_3381), .S(n46), .Z(new_AGEMA_signal_2479) );
  MUX2_X1 PlaintextMUX_MUXInst_35_U1_Ins_0_U1 ( .A(MCOutput[35]), .B(
        new_AGEMA_signal_3383), .S(n46), .Z(StateRegInput[35]) );
  MUX2_X1 PlaintextMUX_MUXInst_35_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2544), .B(
        new_AGEMA_signal_3385), .S(n46), .Z(new_AGEMA_signal_2584) );
  MUX2_X1 PlaintextMUX_MUXInst_35_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2545), .B(
        new_AGEMA_signal_3387), .S(n46), .Z(new_AGEMA_signal_2585) );
  MUX2_X1 PlaintextMUX_MUXInst_38_U1_Ins_0_U1 ( .A(MCOutput[38]), .B(
        new_AGEMA_signal_3389), .S(n46), .Z(StateRegInput[38]) );
  MUX2_X1 PlaintextMUX_MUXInst_38_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2460), .B(
        new_AGEMA_signal_3391), .S(n46), .Z(new_AGEMA_signal_2482) );
  MUX2_X1 PlaintextMUX_MUXInst_38_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2461), .B(
        new_AGEMA_signal_3393), .S(n46), .Z(new_AGEMA_signal_2483) );
  MUX2_X1 PlaintextMUX_MUXInst_39_U1_Ins_0_U1 ( .A(MCOutput[39]), .B(
        new_AGEMA_signal_3395), .S(n46), .Z(StateRegInput[39]) );
  MUX2_X1 PlaintextMUX_MUXInst_39_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2548), .B(
        new_AGEMA_signal_3397), .S(n46), .Z(new_AGEMA_signal_2588) );
  MUX2_X1 PlaintextMUX_MUXInst_39_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2549), .B(
        new_AGEMA_signal_3399), .S(n46), .Z(new_AGEMA_signal_2589) );
  MUX2_X1 PlaintextMUX_MUXInst_42_U1_Ins_0_U1 ( .A(MCOutput[42]), .B(
        new_AGEMA_signal_3401), .S(n46), .Z(StateRegInput[42]) );
  MUX2_X1 PlaintextMUX_MUXInst_42_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2464), .B(
        new_AGEMA_signal_3403), .S(n46), .Z(new_AGEMA_signal_2486) );
  MUX2_X1 PlaintextMUX_MUXInst_42_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2465), .B(
        new_AGEMA_signal_3405), .S(n46), .Z(new_AGEMA_signal_2487) );
  MUX2_X1 PlaintextMUX_MUXInst_43_U1_Ins_0_U1 ( .A(MCOutput[43]), .B(
        new_AGEMA_signal_3407), .S(n46), .Z(StateRegInput[43]) );
  MUX2_X1 PlaintextMUX_MUXInst_43_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2552), .B(
        new_AGEMA_signal_3409), .S(n46), .Z(new_AGEMA_signal_2592) );
  MUX2_X1 PlaintextMUX_MUXInst_43_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2553), .B(
        new_AGEMA_signal_3411), .S(n46), .Z(new_AGEMA_signal_2593) );
  MUX2_X1 PlaintextMUX_MUXInst_46_U1_Ins_0_U1 ( .A(MCOutput[46]), .B(
        new_AGEMA_signal_3413), .S(n46), .Z(StateRegInput[46]) );
  MUX2_X1 PlaintextMUX_MUXInst_46_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2632), .B(
        new_AGEMA_signal_3415), .S(n46), .Z(new_AGEMA_signal_2716) );
  MUX2_X1 PlaintextMUX_MUXInst_46_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2633), .B(
        new_AGEMA_signal_3417), .S(n46), .Z(new_AGEMA_signal_2717) );
  MUX2_X1 PlaintextMUX_MUXInst_47_U1_Ins_0_U1 ( .A(MCOutput[47]), .B(
        new_AGEMA_signal_3419), .S(n45), .Z(StateRegInput[47]) );
  MUX2_X1 PlaintextMUX_MUXInst_47_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2752), .B(
        new_AGEMA_signal_3421), .S(n45), .Z(new_AGEMA_signal_2836) );
  MUX2_X1 PlaintextMUX_MUXInst_47_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2753), .B(
        new_AGEMA_signal_3423), .S(n45), .Z(new_AGEMA_signal_2837) );
  MUX2_X1 PlaintextMUX_MUXInst_50_U1_Ins_0_U1 ( .A(MCOutput[50]), .B(
        new_AGEMA_signal_3425), .S(n45), .Z(StateRegInput[50]) );
  MUX2_X1 PlaintextMUX_MUXInst_50_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2638), .B(
        new_AGEMA_signal_3427), .S(n45), .Z(new_AGEMA_signal_2720) );
  MUX2_X1 PlaintextMUX_MUXInst_50_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2639), .B(
        new_AGEMA_signal_3429), .S(n45), .Z(new_AGEMA_signal_2721) );
  MUX2_X1 PlaintextMUX_MUXInst_51_U1_Ins_0_U1 ( .A(MCOutput[51]), .B(
        new_AGEMA_signal_3431), .S(n45), .Z(StateRegInput[51]) );
  MUX2_X1 PlaintextMUX_MUXInst_51_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2756), .B(
        new_AGEMA_signal_3433), .S(n45), .Z(new_AGEMA_signal_2840) );
  MUX2_X1 PlaintextMUX_MUXInst_51_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2757), .B(
        new_AGEMA_signal_3435), .S(n45), .Z(new_AGEMA_signal_2841) );
  MUX2_X1 PlaintextMUX_MUXInst_54_U1_Ins_0_U1 ( .A(MCOutput[54]), .B(
        new_AGEMA_signal_3437), .S(n45), .Z(StateRegInput[54]) );
  MUX2_X1 PlaintextMUX_MUXInst_54_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2642), .B(
        new_AGEMA_signal_3439), .S(n45), .Z(new_AGEMA_signal_2724) );
  MUX2_X1 PlaintextMUX_MUXInst_54_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2643), .B(
        new_AGEMA_signal_3441), .S(n45), .Z(new_AGEMA_signal_2725) );
  MUX2_X1 PlaintextMUX_MUXInst_55_U1_Ins_0_U1 ( .A(MCOutput[55]), .B(
        new_AGEMA_signal_3443), .S(n45), .Z(StateRegInput[55]) );
  MUX2_X1 PlaintextMUX_MUXInst_55_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2762), .B(
        new_AGEMA_signal_3445), .S(n45), .Z(new_AGEMA_signal_2844) );
  MUX2_X1 PlaintextMUX_MUXInst_55_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2763), .B(
        new_AGEMA_signal_3447), .S(n45), .Z(new_AGEMA_signal_2845) );
  MUX2_X1 PlaintextMUX_MUXInst_58_U1_Ins_0_U1 ( .A(MCOutput[58]), .B(
        new_AGEMA_signal_3449), .S(n45), .Z(StateRegInput[58]) );
  MUX2_X1 PlaintextMUX_MUXInst_58_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2648), .B(
        new_AGEMA_signal_3451), .S(n45), .Z(new_AGEMA_signal_2728) );
  MUX2_X1 PlaintextMUX_MUXInst_58_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2649), .B(
        new_AGEMA_signal_3453), .S(n45), .Z(new_AGEMA_signal_2729) );
  MUX2_X1 PlaintextMUX_MUXInst_59_U1_Ins_0_U1 ( .A(MCOutput[59]), .B(
        new_AGEMA_signal_3455), .S(n45), .Z(StateRegInput[59]) );
  MUX2_X1 PlaintextMUX_MUXInst_59_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2766), .B(
        new_AGEMA_signal_3457), .S(n45), .Z(new_AGEMA_signal_2848) );
  MUX2_X1 PlaintextMUX_MUXInst_59_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2767), .B(
        new_AGEMA_signal_3459), .S(n45), .Z(new_AGEMA_signal_2849) );
  MUX2_X1 PlaintextMUX_MUXInst_62_U1_Ins_0_U1 ( .A(MCOutput[62]), .B(
        new_AGEMA_signal_3461), .S(n45), .Z(StateRegInput[62]) );
  MUX2_X1 PlaintextMUX_MUXInst_62_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2870), .B(
        new_AGEMA_signal_3463), .S(n45), .Z(new_AGEMA_signal_2956) );
  MUX2_X1 PlaintextMUX_MUXInst_62_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2871), .B(
        new_AGEMA_signal_3465), .S(n45), .Z(new_AGEMA_signal_2957) );
  MUX2_X1 PlaintextMUX_MUXInst_63_U1_Ins_0_U1 ( .A(MCOutput[63]), .B(
        new_AGEMA_signal_3467), .S(n45), .Z(StateRegInput[63]) );
  MUX2_X1 PlaintextMUX_MUXInst_63_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2970), .B(
        new_AGEMA_signal_3469), .S(n45), .Z(new_AGEMA_signal_3042) );
  MUX2_X1 PlaintextMUX_MUXInst_63_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2971), .B(
        new_AGEMA_signal_3471), .S(n45), .Z(new_AGEMA_signal_3043) );
  INV_X1 SubCellInst_SboxInst_0_U3_U1 ( .A(SubCellInst_SboxInst_0_YY_1_), .ZN(
        ShiftRowsOutput[7]) );
  INV_X1 SubCellInst_SboxInst_0_U2_U1 ( .A(SubCellInst_SboxInst_0_YY_0_), .ZN(
        ShiftRowsOutput[6]) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U37 ( .A(new_AGEMA_signal_1744), .B(
        Fresh[2]), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U36 ( .A(Fresh[1]), .B(
        SubCellInst_SboxInst_0_Q1), .Z(
        SubCellInst_SboxInst_0_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U35 ( .A(new_AGEMA_signal_1745), .B(
        Fresh[2]), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U34 ( .A(Fresh[0]), .B(
        SubCellInst_SboxInst_0_Q1), .Z(
        SubCellInst_SboxInst_0_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U33 ( .A(Fresh[1]), .B(
        new_AGEMA_signal_1745), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U32 ( .A(new_AGEMA_signal_1744), .B(
        Fresh[0]), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U25 ( .A1(Ciphertext_s2[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U24 ( .A1(Ciphertext_s2[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U23 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND1_U1_U22 ( .A(Fresh[2]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U21 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND1_U1_U19 ( .A(Fresh[1]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND1_U1_U17 ( .A(Fresh[0]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U16 ( .A1(new_AGEMA_signal_1745), 
        .A2(Ciphertext_s2[2]), .ZN(SubCellInst_SboxInst_0_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U15 ( .A1(new_AGEMA_signal_1744), 
        .A2(Ciphertext_s1[2]), .ZN(SubCellInst_SboxInst_0_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_0_Q1), 
        .A2(SubCellInst_SboxInst_0_n3), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND1_U1_n33), .Z(new_AGEMA_signal_1933) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n32), .B(
        SubCellInst_SboxInst_0_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_0_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND1_U1_n30), .Z(new_AGEMA_signal_1932) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n29), .B(
        SubCellInst_SboxInst_0_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_0_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND1_U1_n27), .Z(SubCellInst_SboxInst_0_T0) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n26), .B(
        SubCellInst_SboxInst_0_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_0_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3473), 
        .B(SubCellInst_SboxInst_0_T0), .Z(SubCellInst_SboxInst_0_Q2) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3475), 
        .B(new_AGEMA_signal_1932), .Z(new_AGEMA_signal_2028) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3477), 
        .B(new_AGEMA_signal_1933), .Z(new_AGEMA_signal_2029) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U37 ( .A(new_AGEMA_signal_1746), .B(
        Fresh[5]), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U36 ( .A(Fresh[4]), .B(
        SubCellInst_SboxInst_0_Q4), .Z(
        SubCellInst_SboxInst_0_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U35 ( .A(new_AGEMA_signal_1747), .B(
        Fresh[5]), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U34 ( .A(Fresh[3]), .B(
        SubCellInst_SboxInst_0_Q4), .Z(
        SubCellInst_SboxInst_0_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U33 ( .A(Fresh[4]), .B(
        new_AGEMA_signal_1747), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U32 ( .A(new_AGEMA_signal_1746), .B(
        Fresh[3]), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U25 ( .A1(Ciphertext_s2[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U24 ( .A1(Ciphertext_s2[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U23 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND3_U1_U22 ( .A(Fresh[5]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U21 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND3_U1_U19 ( .A(Fresh[4]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND3_U1_U17 ( .A(Fresh[3]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U16 ( .A1(new_AGEMA_signal_1747), 
        .A2(Ciphertext_s2[2]), .ZN(SubCellInst_SboxInst_0_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U15 ( .A1(new_AGEMA_signal_1746), 
        .A2(Ciphertext_s1[2]), .ZN(SubCellInst_SboxInst_0_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_0_Q4), 
        .A2(SubCellInst_SboxInst_0_n3), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND3_U1_n33), .Z(new_AGEMA_signal_1935) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n32), .B(
        SubCellInst_SboxInst_0_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_0_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND3_U1_n30), .Z(new_AGEMA_signal_1934) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n29), .B(
        SubCellInst_SboxInst_0_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_0_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND3_U1_n27), .Z(SubCellInst_SboxInst_0_T2) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n26), .B(
        SubCellInst_SboxInst_0_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_0_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3479), 
        .B(SubCellInst_SboxInst_0_T2), .Z(SubCellInst_SboxInst_0_Q7) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3481), 
        .B(new_AGEMA_signal_1934), .Z(new_AGEMA_signal_2030) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3483), 
        .B(new_AGEMA_signal_1935), .Z(new_AGEMA_signal_2031) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3485), 
        .B(SubCellInst_SboxInst_0_T0), .Z(SubCellInst_SboxInst_0_L3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3487), 
        .B(new_AGEMA_signal_1932), .Z(new_AGEMA_signal_2032) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3489), 
        .B(new_AGEMA_signal_1933), .Z(new_AGEMA_signal_2033) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L3), .B(SubCellInst_SboxInst_0_T2), .Z(
        SubCellInst_SboxInst_0_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2032), 
        .B(new_AGEMA_signal_1934), .Z(new_AGEMA_signal_2284) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2033), 
        .B(new_AGEMA_signal_1935), .Z(new_AGEMA_signal_2285) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3491), 
        .B(SubCellInst_SboxInst_0_T2), .Z(SubCellInst_SboxInst_0_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3493), 
        .B(new_AGEMA_signal_1934), .Z(new_AGEMA_signal_2156) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3495), 
        .B(new_AGEMA_signal_1935), .Z(new_AGEMA_signal_2157) );
  INV_X1 SubCellInst_SboxInst_1_U3_U1 ( .A(SubCellInst_SboxInst_1_YY_1_), .ZN(
        ShiftRowsOutput[11]) );
  INV_X1 SubCellInst_SboxInst_1_U2_U1 ( .A(SubCellInst_SboxInst_1_YY_0_), .ZN(
        ShiftRowsOutput[10]) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U37 ( .A(new_AGEMA_signal_1756), .B(
        Fresh[8]), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U36 ( .A(Fresh[7]), .B(
        SubCellInst_SboxInst_1_Q1), .Z(
        SubCellInst_SboxInst_1_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U35 ( .A(new_AGEMA_signal_1757), .B(
        Fresh[8]), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U34 ( .A(Fresh[6]), .B(
        SubCellInst_SboxInst_1_Q1), .Z(
        SubCellInst_SboxInst_1_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U33 ( .A(Fresh[7]), .B(
        new_AGEMA_signal_1757), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U32 ( .A(new_AGEMA_signal_1756), .B(
        Fresh[6]), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U25 ( .A1(Ciphertext_s2[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U24 ( .A1(Ciphertext_s2[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U23 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND1_U1_U22 ( .A(Fresh[8]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U21 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND1_U1_U19 ( .A(Fresh[7]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND1_U1_U17 ( .A(Fresh[6]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U16 ( .A1(new_AGEMA_signal_1757), 
        .A2(Ciphertext_s2[6]), .ZN(SubCellInst_SboxInst_1_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U15 ( .A1(new_AGEMA_signal_1756), 
        .A2(Ciphertext_s1[6]), .ZN(SubCellInst_SboxInst_1_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_1_Q1), 
        .A2(SubCellInst_SboxInst_1_n3), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND1_U1_n33), .Z(new_AGEMA_signal_1939) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n32), .B(
        SubCellInst_SboxInst_1_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_1_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND1_U1_n30), .Z(new_AGEMA_signal_1938) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n29), .B(
        SubCellInst_SboxInst_1_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_1_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND1_U1_n27), .Z(SubCellInst_SboxInst_1_T0) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n26), .B(
        SubCellInst_SboxInst_1_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_1_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3497), 
        .B(SubCellInst_SboxInst_1_T0), .Z(SubCellInst_SboxInst_1_Q2) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3499), 
        .B(new_AGEMA_signal_1938), .Z(new_AGEMA_signal_2036) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3501), 
        .B(new_AGEMA_signal_1939), .Z(new_AGEMA_signal_2037) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U37 ( .A(new_AGEMA_signal_1758), .B(
        Fresh[11]), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U36 ( .A(Fresh[10]), .B(
        SubCellInst_SboxInst_1_Q4), .Z(
        SubCellInst_SboxInst_1_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U35 ( .A(new_AGEMA_signal_1759), .B(
        Fresh[11]), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U34 ( .A(Fresh[9]), .B(
        SubCellInst_SboxInst_1_Q4), .Z(
        SubCellInst_SboxInst_1_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U33 ( .A(Fresh[10]), .B(
        new_AGEMA_signal_1759), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U32 ( .A(new_AGEMA_signal_1758), .B(
        Fresh[9]), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U25 ( .A1(Ciphertext_s2[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U24 ( .A1(Ciphertext_s2[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U23 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND3_U1_U22 ( .A(Fresh[11]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U21 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND3_U1_U19 ( .A(Fresh[10]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND3_U1_U17 ( .A(Fresh[9]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U16 ( .A1(new_AGEMA_signal_1759), 
        .A2(Ciphertext_s2[6]), .ZN(SubCellInst_SboxInst_1_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U15 ( .A1(new_AGEMA_signal_1758), 
        .A2(Ciphertext_s1[6]), .ZN(SubCellInst_SboxInst_1_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_1_Q4), 
        .A2(SubCellInst_SboxInst_1_n3), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND3_U1_n33), .Z(new_AGEMA_signal_1941) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n32), .B(
        SubCellInst_SboxInst_1_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_1_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND3_U1_n30), .Z(new_AGEMA_signal_1940) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n29), .B(
        SubCellInst_SboxInst_1_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_1_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND3_U1_n27), .Z(SubCellInst_SboxInst_1_T2) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n26), .B(
        SubCellInst_SboxInst_1_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_1_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3503), 
        .B(SubCellInst_SboxInst_1_T2), .Z(SubCellInst_SboxInst_1_Q7) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3505), 
        .B(new_AGEMA_signal_1940), .Z(new_AGEMA_signal_2038) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3507), 
        .B(new_AGEMA_signal_1941), .Z(new_AGEMA_signal_2039) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3509), 
        .B(SubCellInst_SboxInst_1_T0), .Z(SubCellInst_SboxInst_1_L3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3511), 
        .B(new_AGEMA_signal_1938), .Z(new_AGEMA_signal_2040) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3513), 
        .B(new_AGEMA_signal_1939), .Z(new_AGEMA_signal_2041) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L3), .B(SubCellInst_SboxInst_1_T2), .Z(
        SubCellInst_SboxInst_1_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2040), 
        .B(new_AGEMA_signal_1940), .Z(new_AGEMA_signal_2288) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2041), 
        .B(new_AGEMA_signal_1941), .Z(new_AGEMA_signal_2289) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3515), 
        .B(SubCellInst_SboxInst_1_T2), .Z(SubCellInst_SboxInst_1_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3517), 
        .B(new_AGEMA_signal_1940), .Z(new_AGEMA_signal_2164) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3519), 
        .B(new_AGEMA_signal_1941), .Z(new_AGEMA_signal_2165) );
  INV_X1 SubCellInst_SboxInst_2_U3_U1 ( .A(SubCellInst_SboxInst_2_YY_1_), .ZN(
        ShiftRowsOutput[15]) );
  INV_X1 SubCellInst_SboxInst_2_U2_U1 ( .A(SubCellInst_SboxInst_2_YY_0_), .ZN(
        ShiftRowsOutput[14]) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U37 ( .A(new_AGEMA_signal_1768), .B(
        Fresh[14]), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U36 ( .A(Fresh[13]), .B(
        SubCellInst_SboxInst_2_Q1), .Z(
        SubCellInst_SboxInst_2_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U35 ( .A(new_AGEMA_signal_1769), .B(
        Fresh[14]), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U34 ( .A(Fresh[12]), .B(
        SubCellInst_SboxInst_2_Q1), .Z(
        SubCellInst_SboxInst_2_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U33 ( .A(Fresh[13]), .B(
        new_AGEMA_signal_1769), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U32 ( .A(new_AGEMA_signal_1768), .B(
        Fresh[12]), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U25 ( .A1(Ciphertext_s2[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U24 ( .A1(Ciphertext_s2[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U23 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND1_U1_U22 ( .A(Fresh[14]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U21 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND1_U1_U19 ( .A(Fresh[13]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND1_U1_U17 ( .A(Fresh[12]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U16 ( .A1(new_AGEMA_signal_1769), 
        .A2(Ciphertext_s2[10]), .ZN(SubCellInst_SboxInst_2_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U15 ( .A1(new_AGEMA_signal_1768), 
        .A2(Ciphertext_s1[10]), .ZN(SubCellInst_SboxInst_2_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_2_Q1), 
        .A2(SubCellInst_SboxInst_2_n3), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND1_U1_n33), .Z(new_AGEMA_signal_1945) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n32), .B(
        SubCellInst_SboxInst_2_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_2_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND1_U1_n30), .Z(new_AGEMA_signal_1944) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n29), .B(
        SubCellInst_SboxInst_2_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_2_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND1_U1_n27), .Z(SubCellInst_SboxInst_2_T0) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n26), .B(
        SubCellInst_SboxInst_2_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_2_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3521), 
        .B(SubCellInst_SboxInst_2_T0), .Z(SubCellInst_SboxInst_2_Q2) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3523), 
        .B(new_AGEMA_signal_1944), .Z(new_AGEMA_signal_2044) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3525), 
        .B(new_AGEMA_signal_1945), .Z(new_AGEMA_signal_2045) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U37 ( .A(new_AGEMA_signal_1770), .B(
        Fresh[17]), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U36 ( .A(Fresh[16]), .B(
        SubCellInst_SboxInst_2_Q4), .Z(
        SubCellInst_SboxInst_2_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U35 ( .A(new_AGEMA_signal_1771), .B(
        Fresh[17]), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U34 ( .A(Fresh[15]), .B(
        SubCellInst_SboxInst_2_Q4), .Z(
        SubCellInst_SboxInst_2_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U33 ( .A(Fresh[16]), .B(
        new_AGEMA_signal_1771), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U32 ( .A(new_AGEMA_signal_1770), .B(
        Fresh[15]), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U25 ( .A1(Ciphertext_s2[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U24 ( .A1(Ciphertext_s2[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U23 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND3_U1_U22 ( .A(Fresh[17]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U21 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND3_U1_U19 ( .A(Fresh[16]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND3_U1_U17 ( .A(Fresh[15]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U16 ( .A1(new_AGEMA_signal_1771), 
        .A2(Ciphertext_s2[10]), .ZN(SubCellInst_SboxInst_2_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U15 ( .A1(new_AGEMA_signal_1770), 
        .A2(Ciphertext_s1[10]), .ZN(SubCellInst_SboxInst_2_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_2_Q4), 
        .A2(SubCellInst_SboxInst_2_n3), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND3_U1_n33), .Z(new_AGEMA_signal_1947) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n32), .B(
        SubCellInst_SboxInst_2_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_2_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND3_U1_n30), .Z(new_AGEMA_signal_1946) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n29), .B(
        SubCellInst_SboxInst_2_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_2_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND3_U1_n27), .Z(SubCellInst_SboxInst_2_T2) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n26), .B(
        SubCellInst_SboxInst_2_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_2_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3527), 
        .B(SubCellInst_SboxInst_2_T2), .Z(SubCellInst_SboxInst_2_Q7) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3529), 
        .B(new_AGEMA_signal_1946), .Z(new_AGEMA_signal_2046) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3531), 
        .B(new_AGEMA_signal_1947), .Z(new_AGEMA_signal_2047) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3533), 
        .B(SubCellInst_SboxInst_2_T0), .Z(SubCellInst_SboxInst_2_L3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3535), 
        .B(new_AGEMA_signal_1944), .Z(new_AGEMA_signal_2048) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3537), 
        .B(new_AGEMA_signal_1945), .Z(new_AGEMA_signal_2049) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L3), .B(SubCellInst_SboxInst_2_T2), .Z(
        SubCellInst_SboxInst_2_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2048), 
        .B(new_AGEMA_signal_1946), .Z(new_AGEMA_signal_2292) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2049), 
        .B(new_AGEMA_signal_1947), .Z(new_AGEMA_signal_2293) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3539), 
        .B(SubCellInst_SboxInst_2_T2), .Z(SubCellInst_SboxInst_2_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3541), 
        .B(new_AGEMA_signal_1946), .Z(new_AGEMA_signal_2172) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3543), 
        .B(new_AGEMA_signal_1947), .Z(new_AGEMA_signal_2173) );
  INV_X1 SubCellInst_SboxInst_3_U3_U1 ( .A(SubCellInst_SboxInst_3_YY_1_), .ZN(
        ShiftRowsOutput[3]) );
  INV_X1 SubCellInst_SboxInst_3_U2_U1 ( .A(SubCellInst_SboxInst_3_YY_0_), .ZN(
        ShiftRowsOutput[2]) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U37 ( .A(new_AGEMA_signal_1780), .B(
        Fresh[20]), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U36 ( .A(Fresh[19]), .B(
        SubCellInst_SboxInst_3_Q1), .Z(
        SubCellInst_SboxInst_3_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U35 ( .A(new_AGEMA_signal_1781), .B(
        Fresh[20]), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U34 ( .A(Fresh[18]), .B(
        SubCellInst_SboxInst_3_Q1), .Z(
        SubCellInst_SboxInst_3_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U33 ( .A(Fresh[19]), .B(
        new_AGEMA_signal_1781), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U32 ( .A(new_AGEMA_signal_1780), .B(
        Fresh[18]), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U25 ( .A1(Ciphertext_s2[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U24 ( .A1(Ciphertext_s2[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U23 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND1_U1_U22 ( .A(Fresh[20]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U21 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND1_U1_U19 ( .A(Fresh[19]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND1_U1_U17 ( .A(Fresh[18]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U16 ( .A1(new_AGEMA_signal_1781), 
        .A2(Ciphertext_s2[14]), .ZN(SubCellInst_SboxInst_3_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U15 ( .A1(new_AGEMA_signal_1780), 
        .A2(Ciphertext_s1[14]), .ZN(SubCellInst_SboxInst_3_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_3_Q1), 
        .A2(SubCellInst_SboxInst_3_n3), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND1_U1_n33), .Z(new_AGEMA_signal_1951) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n32), .B(
        SubCellInst_SboxInst_3_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_3_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND1_U1_n30), .Z(new_AGEMA_signal_1950) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n29), .B(
        SubCellInst_SboxInst_3_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_3_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND1_U1_n27), .Z(SubCellInst_SboxInst_3_T0) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n26), .B(
        SubCellInst_SboxInst_3_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_3_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3545), 
        .B(SubCellInst_SboxInst_3_T0), .Z(SubCellInst_SboxInst_3_Q2) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3547), 
        .B(new_AGEMA_signal_1950), .Z(new_AGEMA_signal_2052) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3549), 
        .B(new_AGEMA_signal_1951), .Z(new_AGEMA_signal_2053) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U37 ( .A(new_AGEMA_signal_1782), .B(
        Fresh[23]), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U36 ( .A(Fresh[22]), .B(
        SubCellInst_SboxInst_3_Q4), .Z(
        SubCellInst_SboxInst_3_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U35 ( .A(new_AGEMA_signal_1783), .B(
        Fresh[23]), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U34 ( .A(Fresh[21]), .B(
        SubCellInst_SboxInst_3_Q4), .Z(
        SubCellInst_SboxInst_3_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U33 ( .A(Fresh[22]), .B(
        new_AGEMA_signal_1783), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U32 ( .A(new_AGEMA_signal_1782), .B(
        Fresh[21]), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U25 ( .A1(Ciphertext_s2[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U24 ( .A1(Ciphertext_s2[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U23 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND3_U1_U22 ( .A(Fresh[23]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U21 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND3_U1_U19 ( .A(Fresh[22]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND3_U1_U17 ( .A(Fresh[21]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U16 ( .A1(new_AGEMA_signal_1783), 
        .A2(Ciphertext_s2[14]), .ZN(SubCellInst_SboxInst_3_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U15 ( .A1(new_AGEMA_signal_1782), 
        .A2(Ciphertext_s1[14]), .ZN(SubCellInst_SboxInst_3_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_3_Q4), 
        .A2(SubCellInst_SboxInst_3_n3), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND3_U1_n33), .Z(new_AGEMA_signal_1953) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n32), .B(
        SubCellInst_SboxInst_3_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_3_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND3_U1_n30), .Z(new_AGEMA_signal_1952) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n29), .B(
        SubCellInst_SboxInst_3_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_3_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND3_U1_n27), .Z(SubCellInst_SboxInst_3_T2) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n26), .B(
        SubCellInst_SboxInst_3_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_3_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3551), 
        .B(SubCellInst_SboxInst_3_T2), .Z(SubCellInst_SboxInst_3_Q7) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3553), 
        .B(new_AGEMA_signal_1952), .Z(new_AGEMA_signal_2054) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3555), 
        .B(new_AGEMA_signal_1953), .Z(new_AGEMA_signal_2055) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3557), 
        .B(SubCellInst_SboxInst_3_T0), .Z(SubCellInst_SboxInst_3_L3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3559), 
        .B(new_AGEMA_signal_1950), .Z(new_AGEMA_signal_2056) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3561), 
        .B(new_AGEMA_signal_1951), .Z(new_AGEMA_signal_2057) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L3), .B(SubCellInst_SboxInst_3_T2), .Z(
        SubCellInst_SboxInst_3_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2056), 
        .B(new_AGEMA_signal_1952), .Z(new_AGEMA_signal_2296) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2057), 
        .B(new_AGEMA_signal_1953), .Z(new_AGEMA_signal_2297) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3563), 
        .B(SubCellInst_SboxInst_3_T2), .Z(SubCellInst_SboxInst_3_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3565), 
        .B(new_AGEMA_signal_1952), .Z(new_AGEMA_signal_2180) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3567), 
        .B(new_AGEMA_signal_1953), .Z(new_AGEMA_signal_2181) );
  INV_X1 SubCellInst_SboxInst_4_U3_U1 ( .A(SubCellInst_SboxInst_4_YY_1_), .ZN(
        ShiftRowsOutput[27]) );
  INV_X1 SubCellInst_SboxInst_4_U2_U1 ( .A(SubCellInst_SboxInst_4_YY_0_), .ZN(
        ShiftRowsOutput[26]) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U37 ( .A(new_AGEMA_signal_1792), .B(
        Fresh[26]), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U36 ( .A(Fresh[25]), .B(
        SubCellInst_SboxInst_4_Q1), .Z(
        SubCellInst_SboxInst_4_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U35 ( .A(new_AGEMA_signal_1793), .B(
        Fresh[26]), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U34 ( .A(Fresh[24]), .B(
        SubCellInst_SboxInst_4_Q1), .Z(
        SubCellInst_SboxInst_4_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U33 ( .A(Fresh[25]), .B(
        new_AGEMA_signal_1793), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U32 ( .A(new_AGEMA_signal_1792), .B(
        Fresh[24]), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U25 ( .A1(Ciphertext_s2[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U24 ( .A1(Ciphertext_s2[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U23 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND1_U1_U22 ( .A(Fresh[26]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U21 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND1_U1_U19 ( .A(Fresh[25]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND1_U1_U17 ( .A(Fresh[24]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U16 ( .A1(new_AGEMA_signal_1793), 
        .A2(Ciphertext_s2[18]), .ZN(SubCellInst_SboxInst_4_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U15 ( .A1(new_AGEMA_signal_1792), 
        .A2(Ciphertext_s1[18]), .ZN(SubCellInst_SboxInst_4_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_4_Q1), 
        .A2(SubCellInst_SboxInst_4_n3), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND1_U1_n33), .Z(new_AGEMA_signal_1957) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n32), .B(
        SubCellInst_SboxInst_4_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_4_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND1_U1_n30), .Z(new_AGEMA_signal_1956) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n29), .B(
        SubCellInst_SboxInst_4_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_4_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND1_U1_n27), .Z(SubCellInst_SboxInst_4_T0) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n26), .B(
        SubCellInst_SboxInst_4_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_4_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3569), 
        .B(SubCellInst_SboxInst_4_T0), .Z(SubCellInst_SboxInst_4_Q2) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3571), 
        .B(new_AGEMA_signal_1956), .Z(new_AGEMA_signal_2060) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3573), 
        .B(new_AGEMA_signal_1957), .Z(new_AGEMA_signal_2061) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U37 ( .A(new_AGEMA_signal_1794), .B(
        Fresh[29]), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U36 ( .A(Fresh[28]), .B(
        SubCellInst_SboxInst_4_Q4), .Z(
        SubCellInst_SboxInst_4_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U35 ( .A(new_AGEMA_signal_1795), .B(
        Fresh[29]), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U34 ( .A(Fresh[27]), .B(
        SubCellInst_SboxInst_4_Q4), .Z(
        SubCellInst_SboxInst_4_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U33 ( .A(Fresh[28]), .B(
        new_AGEMA_signal_1795), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U32 ( .A(new_AGEMA_signal_1794), .B(
        Fresh[27]), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U25 ( .A1(Ciphertext_s2[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U24 ( .A1(Ciphertext_s2[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U23 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND3_U1_U22 ( .A(Fresh[29]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U21 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND3_U1_U19 ( .A(Fresh[28]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND3_U1_U17 ( .A(Fresh[27]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U16 ( .A1(new_AGEMA_signal_1795), 
        .A2(Ciphertext_s2[18]), .ZN(SubCellInst_SboxInst_4_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U15 ( .A1(new_AGEMA_signal_1794), 
        .A2(Ciphertext_s1[18]), .ZN(SubCellInst_SboxInst_4_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_4_Q4), 
        .A2(SubCellInst_SboxInst_4_n3), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND3_U1_n33), .Z(new_AGEMA_signal_1959) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n32), .B(
        SubCellInst_SboxInst_4_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_4_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND3_U1_n30), .Z(new_AGEMA_signal_1958) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n29), .B(
        SubCellInst_SboxInst_4_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_4_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND3_U1_n27), .Z(SubCellInst_SboxInst_4_T2) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n26), .B(
        SubCellInst_SboxInst_4_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_4_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3575), 
        .B(SubCellInst_SboxInst_4_T2), .Z(SubCellInst_SboxInst_4_Q7) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3577), 
        .B(new_AGEMA_signal_1958), .Z(new_AGEMA_signal_2062) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3579), 
        .B(new_AGEMA_signal_1959), .Z(new_AGEMA_signal_2063) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3581), 
        .B(SubCellInst_SboxInst_4_T0), .Z(SubCellInst_SboxInst_4_L3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3583), 
        .B(new_AGEMA_signal_1956), .Z(new_AGEMA_signal_2064) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3585), 
        .B(new_AGEMA_signal_1957), .Z(new_AGEMA_signal_2065) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L3), .B(SubCellInst_SboxInst_4_T2), .Z(
        SubCellInst_SboxInst_4_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2064), 
        .B(new_AGEMA_signal_1958), .Z(new_AGEMA_signal_2300) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2065), 
        .B(new_AGEMA_signal_1959), .Z(new_AGEMA_signal_2301) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3587), 
        .B(SubCellInst_SboxInst_4_T2), .Z(SubCellInst_SboxInst_4_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3589), 
        .B(new_AGEMA_signal_1958), .Z(new_AGEMA_signal_2188) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3591), 
        .B(new_AGEMA_signal_1959), .Z(new_AGEMA_signal_2189) );
  INV_X1 SubCellInst_SboxInst_5_U3_U1 ( .A(SubCellInst_SboxInst_5_YY_1_), .ZN(
        ShiftRowsOutput[31]) );
  INV_X1 SubCellInst_SboxInst_5_U2_U1 ( .A(SubCellInst_SboxInst_5_YY_0_), .ZN(
        ShiftRowsOutput[30]) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U37 ( .A(new_AGEMA_signal_1804), .B(
        Fresh[32]), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U36 ( .A(Fresh[31]), .B(
        SubCellInst_SboxInst_5_Q1), .Z(
        SubCellInst_SboxInst_5_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U35 ( .A(new_AGEMA_signal_1805), .B(
        Fresh[32]), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U34 ( .A(Fresh[30]), .B(
        SubCellInst_SboxInst_5_Q1), .Z(
        SubCellInst_SboxInst_5_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U33 ( .A(Fresh[31]), .B(
        new_AGEMA_signal_1805), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U32 ( .A(new_AGEMA_signal_1804), .B(
        Fresh[30]), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U25 ( .A1(Ciphertext_s2[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U24 ( .A1(Ciphertext_s2[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U23 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND1_U1_U22 ( .A(Fresh[32]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U21 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND1_U1_U19 ( .A(Fresh[31]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND1_U1_U17 ( .A(Fresh[30]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U16 ( .A1(new_AGEMA_signal_1805), 
        .A2(Ciphertext_s2[22]), .ZN(SubCellInst_SboxInst_5_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U15 ( .A1(new_AGEMA_signal_1804), 
        .A2(Ciphertext_s1[22]), .ZN(SubCellInst_SboxInst_5_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_5_Q1), 
        .A2(SubCellInst_SboxInst_5_n3), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND1_U1_n33), .Z(new_AGEMA_signal_1963) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n32), .B(
        SubCellInst_SboxInst_5_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_5_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND1_U1_n30), .Z(new_AGEMA_signal_1962) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n29), .B(
        SubCellInst_SboxInst_5_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_5_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND1_U1_n27), .Z(SubCellInst_SboxInst_5_T0) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n26), .B(
        SubCellInst_SboxInst_5_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_5_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3593), 
        .B(SubCellInst_SboxInst_5_T0), .Z(SubCellInst_SboxInst_5_Q2) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3595), 
        .B(new_AGEMA_signal_1962), .Z(new_AGEMA_signal_2068) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3597), 
        .B(new_AGEMA_signal_1963), .Z(new_AGEMA_signal_2069) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U37 ( .A(new_AGEMA_signal_1806), .B(
        Fresh[35]), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U36 ( .A(Fresh[34]), .B(
        SubCellInst_SboxInst_5_Q4), .Z(
        SubCellInst_SboxInst_5_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U35 ( .A(new_AGEMA_signal_1807), .B(
        Fresh[35]), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U34 ( .A(Fresh[33]), .B(
        SubCellInst_SboxInst_5_Q4), .Z(
        SubCellInst_SboxInst_5_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U33 ( .A(Fresh[34]), .B(
        new_AGEMA_signal_1807), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U32 ( .A(new_AGEMA_signal_1806), .B(
        Fresh[33]), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U25 ( .A1(Ciphertext_s2[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U24 ( .A1(Ciphertext_s2[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U23 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND3_U1_U22 ( .A(Fresh[35]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U21 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND3_U1_U19 ( .A(Fresh[34]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND3_U1_U17 ( .A(Fresh[33]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U16 ( .A1(new_AGEMA_signal_1807), 
        .A2(Ciphertext_s2[22]), .ZN(SubCellInst_SboxInst_5_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U15 ( .A1(new_AGEMA_signal_1806), 
        .A2(Ciphertext_s1[22]), .ZN(SubCellInst_SboxInst_5_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_5_Q4), 
        .A2(SubCellInst_SboxInst_5_n3), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND3_U1_n33), .Z(new_AGEMA_signal_1965) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n32), .B(
        SubCellInst_SboxInst_5_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_5_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND3_U1_n30), .Z(new_AGEMA_signal_1964) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n29), .B(
        SubCellInst_SboxInst_5_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_5_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND3_U1_n27), .Z(SubCellInst_SboxInst_5_T2) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n26), .B(
        SubCellInst_SboxInst_5_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_5_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3599), 
        .B(SubCellInst_SboxInst_5_T2), .Z(SubCellInst_SboxInst_5_Q7) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3601), 
        .B(new_AGEMA_signal_1964), .Z(new_AGEMA_signal_2070) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3603), 
        .B(new_AGEMA_signal_1965), .Z(new_AGEMA_signal_2071) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3605), 
        .B(SubCellInst_SboxInst_5_T0), .Z(SubCellInst_SboxInst_5_L3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3607), 
        .B(new_AGEMA_signal_1962), .Z(new_AGEMA_signal_2072) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3609), 
        .B(new_AGEMA_signal_1963), .Z(new_AGEMA_signal_2073) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L3), .B(SubCellInst_SboxInst_5_T2), .Z(
        SubCellInst_SboxInst_5_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2072), 
        .B(new_AGEMA_signal_1964), .Z(new_AGEMA_signal_2304) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2073), 
        .B(new_AGEMA_signal_1965), .Z(new_AGEMA_signal_2305) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3611), 
        .B(SubCellInst_SboxInst_5_T2), .Z(SubCellInst_SboxInst_5_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3613), 
        .B(new_AGEMA_signal_1964), .Z(new_AGEMA_signal_2196) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3615), 
        .B(new_AGEMA_signal_1965), .Z(new_AGEMA_signal_2197) );
  INV_X1 SubCellInst_SboxInst_6_U3_U1 ( .A(SubCellInst_SboxInst_6_YY_1_), .ZN(
        ShiftRowsOutput[19]) );
  INV_X1 SubCellInst_SboxInst_6_U2_U1 ( .A(SubCellInst_SboxInst_6_YY_0_), .ZN(
        ShiftRowsOutput[18]) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U37 ( .A(new_AGEMA_signal_1816), .B(
        Fresh[38]), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U36 ( .A(Fresh[37]), .B(
        SubCellInst_SboxInst_6_Q1), .Z(
        SubCellInst_SboxInst_6_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U35 ( .A(new_AGEMA_signal_1817), .B(
        Fresh[38]), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U34 ( .A(Fresh[36]), .B(
        SubCellInst_SboxInst_6_Q1), .Z(
        SubCellInst_SboxInst_6_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U33 ( .A(Fresh[37]), .B(
        new_AGEMA_signal_1817), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U32 ( .A(new_AGEMA_signal_1816), .B(
        Fresh[36]), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U25 ( .A1(Ciphertext_s2[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U24 ( .A1(Ciphertext_s2[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U23 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND1_U1_U22 ( .A(Fresh[38]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U21 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND1_U1_U19 ( .A(Fresh[37]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND1_U1_U17 ( .A(Fresh[36]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U16 ( .A1(new_AGEMA_signal_1817), 
        .A2(Ciphertext_s2[26]), .ZN(SubCellInst_SboxInst_6_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U15 ( .A1(new_AGEMA_signal_1816), 
        .A2(Ciphertext_s1[26]), .ZN(SubCellInst_SboxInst_6_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_6_Q1), 
        .A2(SubCellInst_SboxInst_6_n3), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND1_U1_n33), .Z(new_AGEMA_signal_1969) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n32), .B(
        SubCellInst_SboxInst_6_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_6_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND1_U1_n30), .Z(new_AGEMA_signal_1968) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n29), .B(
        SubCellInst_SboxInst_6_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_6_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND1_U1_n27), .Z(SubCellInst_SboxInst_6_T0) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n26), .B(
        SubCellInst_SboxInst_6_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_6_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3617), 
        .B(SubCellInst_SboxInst_6_T0), .Z(SubCellInst_SboxInst_6_Q2) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3619), 
        .B(new_AGEMA_signal_1968), .Z(new_AGEMA_signal_2076) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3621), 
        .B(new_AGEMA_signal_1969), .Z(new_AGEMA_signal_2077) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U37 ( .A(new_AGEMA_signal_1818), .B(
        Fresh[41]), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U36 ( .A(Fresh[40]), .B(
        SubCellInst_SboxInst_6_Q4), .Z(
        SubCellInst_SboxInst_6_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U35 ( .A(new_AGEMA_signal_1819), .B(
        Fresh[41]), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U34 ( .A(Fresh[39]), .B(
        SubCellInst_SboxInst_6_Q4), .Z(
        SubCellInst_SboxInst_6_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U33 ( .A(Fresh[40]), .B(
        new_AGEMA_signal_1819), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U32 ( .A(new_AGEMA_signal_1818), .B(
        Fresh[39]), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U25 ( .A1(Ciphertext_s2[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U24 ( .A1(Ciphertext_s2[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U23 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND3_U1_U22 ( .A(Fresh[41]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U21 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND3_U1_U19 ( .A(Fresh[40]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND3_U1_U17 ( .A(Fresh[39]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U16 ( .A1(new_AGEMA_signal_1819), 
        .A2(Ciphertext_s2[26]), .ZN(SubCellInst_SboxInst_6_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U15 ( .A1(new_AGEMA_signal_1818), 
        .A2(Ciphertext_s1[26]), .ZN(SubCellInst_SboxInst_6_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_6_Q4), 
        .A2(SubCellInst_SboxInst_6_n3), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND3_U1_n33), .Z(new_AGEMA_signal_1971) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n32), .B(
        SubCellInst_SboxInst_6_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_6_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND3_U1_n30), .Z(new_AGEMA_signal_1970) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n29), .B(
        SubCellInst_SboxInst_6_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_6_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND3_U1_n27), .Z(SubCellInst_SboxInst_6_T2) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n26), .B(
        SubCellInst_SboxInst_6_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_6_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3623), 
        .B(SubCellInst_SboxInst_6_T2), .Z(SubCellInst_SboxInst_6_Q7) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3625), 
        .B(new_AGEMA_signal_1970), .Z(new_AGEMA_signal_2078) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3627), 
        .B(new_AGEMA_signal_1971), .Z(new_AGEMA_signal_2079) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3629), 
        .B(SubCellInst_SboxInst_6_T0), .Z(SubCellInst_SboxInst_6_L3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3631), 
        .B(new_AGEMA_signal_1968), .Z(new_AGEMA_signal_2080) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3633), 
        .B(new_AGEMA_signal_1969), .Z(new_AGEMA_signal_2081) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L3), .B(SubCellInst_SboxInst_6_T2), .Z(
        SubCellInst_SboxInst_6_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2080), 
        .B(new_AGEMA_signal_1970), .Z(new_AGEMA_signal_2308) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2081), 
        .B(new_AGEMA_signal_1971), .Z(new_AGEMA_signal_2309) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3635), 
        .B(SubCellInst_SboxInst_6_T2), .Z(SubCellInst_SboxInst_6_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3637), 
        .B(new_AGEMA_signal_1970), .Z(new_AGEMA_signal_2204) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3639), 
        .B(new_AGEMA_signal_1971), .Z(new_AGEMA_signal_2205) );
  INV_X1 SubCellInst_SboxInst_7_U3_U1 ( .A(SubCellInst_SboxInst_7_YY_1_), .ZN(
        ShiftRowsOutput[23]) );
  INV_X1 SubCellInst_SboxInst_7_U2_U1 ( .A(SubCellInst_SboxInst_7_YY_0_), .ZN(
        ShiftRowsOutput[22]) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U37 ( .A(new_AGEMA_signal_1828), .B(
        Fresh[44]), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U36 ( .A(Fresh[43]), .B(
        SubCellInst_SboxInst_7_Q1), .Z(
        SubCellInst_SboxInst_7_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U35 ( .A(new_AGEMA_signal_1829), .B(
        Fresh[44]), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U34 ( .A(Fresh[42]), .B(
        SubCellInst_SboxInst_7_Q1), .Z(
        SubCellInst_SboxInst_7_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U33 ( .A(Fresh[43]), .B(
        new_AGEMA_signal_1829), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U32 ( .A(new_AGEMA_signal_1828), .B(
        Fresh[42]), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U25 ( .A1(Ciphertext_s2[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U24 ( .A1(Ciphertext_s2[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U23 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND1_U1_U22 ( .A(Fresh[44]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U21 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND1_U1_U19 ( .A(Fresh[43]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND1_U1_U17 ( .A(Fresh[42]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U16 ( .A1(new_AGEMA_signal_1829), 
        .A2(Ciphertext_s2[30]), .ZN(SubCellInst_SboxInst_7_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U15 ( .A1(new_AGEMA_signal_1828), 
        .A2(Ciphertext_s1[30]), .ZN(SubCellInst_SboxInst_7_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_7_Q1), 
        .A2(SubCellInst_SboxInst_7_n3), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND1_U1_n33), .Z(new_AGEMA_signal_1975) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n32), .B(
        SubCellInst_SboxInst_7_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_7_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND1_U1_n30), .Z(new_AGEMA_signal_1974) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n29), .B(
        SubCellInst_SboxInst_7_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_7_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND1_U1_n27), .Z(SubCellInst_SboxInst_7_T0) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n26), .B(
        SubCellInst_SboxInst_7_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_7_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3641), 
        .B(SubCellInst_SboxInst_7_T0), .Z(SubCellInst_SboxInst_7_Q2) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3643), 
        .B(new_AGEMA_signal_1974), .Z(new_AGEMA_signal_2084) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3645), 
        .B(new_AGEMA_signal_1975), .Z(new_AGEMA_signal_2085) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U37 ( .A(new_AGEMA_signal_1830), .B(
        Fresh[47]), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U36 ( .A(Fresh[46]), .B(
        SubCellInst_SboxInst_7_Q4), .Z(
        SubCellInst_SboxInst_7_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U35 ( .A(new_AGEMA_signal_1831), .B(
        Fresh[47]), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U34 ( .A(Fresh[45]), .B(
        SubCellInst_SboxInst_7_Q4), .Z(
        SubCellInst_SboxInst_7_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U33 ( .A(Fresh[46]), .B(
        new_AGEMA_signal_1831), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U32 ( .A(new_AGEMA_signal_1830), .B(
        Fresh[45]), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U25 ( .A1(Ciphertext_s2[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U24 ( .A1(Ciphertext_s2[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U23 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND3_U1_U22 ( .A(Fresh[47]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U21 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND3_U1_U19 ( .A(Fresh[46]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND3_U1_U17 ( .A(Fresh[45]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U16 ( .A1(new_AGEMA_signal_1831), 
        .A2(Ciphertext_s2[30]), .ZN(SubCellInst_SboxInst_7_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U15 ( .A1(new_AGEMA_signal_1830), 
        .A2(Ciphertext_s1[30]), .ZN(SubCellInst_SboxInst_7_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_7_Q4), 
        .A2(SubCellInst_SboxInst_7_n3), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND3_U1_n33), .Z(new_AGEMA_signal_1977) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n32), .B(
        SubCellInst_SboxInst_7_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_7_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND3_U1_n30), .Z(new_AGEMA_signal_1976) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n29), .B(
        SubCellInst_SboxInst_7_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_7_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND3_U1_n27), .Z(SubCellInst_SboxInst_7_T2) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n26), .B(
        SubCellInst_SboxInst_7_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_7_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3647), 
        .B(SubCellInst_SboxInst_7_T2), .Z(SubCellInst_SboxInst_7_Q7) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3649), 
        .B(new_AGEMA_signal_1976), .Z(new_AGEMA_signal_2086) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3651), 
        .B(new_AGEMA_signal_1977), .Z(new_AGEMA_signal_2087) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3653), 
        .B(SubCellInst_SboxInst_7_T0), .Z(SubCellInst_SboxInst_7_L3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3655), 
        .B(new_AGEMA_signal_1974), .Z(new_AGEMA_signal_2088) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3657), 
        .B(new_AGEMA_signal_1975), .Z(new_AGEMA_signal_2089) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L3), .B(SubCellInst_SboxInst_7_T2), .Z(
        SubCellInst_SboxInst_7_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2088), 
        .B(new_AGEMA_signal_1976), .Z(new_AGEMA_signal_2312) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2089), 
        .B(new_AGEMA_signal_1977), .Z(new_AGEMA_signal_2313) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3659), 
        .B(SubCellInst_SboxInst_7_T2), .Z(SubCellInst_SboxInst_7_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3661), 
        .B(new_AGEMA_signal_1976), .Z(new_AGEMA_signal_2212) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3663), 
        .B(new_AGEMA_signal_1977), .Z(new_AGEMA_signal_2213) );
  INV_X1 SubCellInst_SboxInst_8_U3_U1 ( .A(SubCellInst_SboxInst_8_YY_1_), .ZN(
        AddRoundConstantOutput[35]) );
  INV_X1 SubCellInst_SboxInst_8_U2_U1 ( .A(SubCellInst_SboxInst_8_YY_0_), .ZN(
        AddRoundConstantOutput[34]) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U37 ( .A(new_AGEMA_signal_1840), .B(
        Fresh[50]), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U36 ( .A(Fresh[49]), .B(
        SubCellInst_SboxInst_8_Q1), .Z(
        SubCellInst_SboxInst_8_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U35 ( .A(new_AGEMA_signal_1841), .B(
        Fresh[50]), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U34 ( .A(Fresh[48]), .B(
        SubCellInst_SboxInst_8_Q1), .Z(
        SubCellInst_SboxInst_8_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U33 ( .A(Fresh[49]), .B(
        new_AGEMA_signal_1841), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U32 ( .A(new_AGEMA_signal_1840), .B(
        Fresh[48]), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U25 ( .A1(Ciphertext_s2[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U24 ( .A1(Ciphertext_s2[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U23 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND1_U1_U22 ( .A(Fresh[50]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U21 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND1_U1_U19 ( .A(Fresh[49]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND1_U1_U17 ( .A(Fresh[48]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U16 ( .A1(new_AGEMA_signal_1841), 
        .A2(Ciphertext_s2[34]), .ZN(SubCellInst_SboxInst_8_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U15 ( .A1(new_AGEMA_signal_1840), 
        .A2(Ciphertext_s1[34]), .ZN(SubCellInst_SboxInst_8_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_8_Q1), 
        .A2(SubCellInst_SboxInst_8_n3), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND1_U1_n33), .Z(new_AGEMA_signal_1981) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n32), .B(
        SubCellInst_SboxInst_8_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_8_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND1_U1_n30), .Z(new_AGEMA_signal_1980) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n29), .B(
        SubCellInst_SboxInst_8_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_8_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND1_U1_n27), .Z(SubCellInst_SboxInst_8_T0) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n26), .B(
        SubCellInst_SboxInst_8_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_8_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3665), 
        .B(SubCellInst_SboxInst_8_T0), .Z(SubCellInst_SboxInst_8_Q2) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3667), 
        .B(new_AGEMA_signal_1980), .Z(new_AGEMA_signal_2092) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3669), 
        .B(new_AGEMA_signal_1981), .Z(new_AGEMA_signal_2093) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U37 ( .A(new_AGEMA_signal_1842), .B(
        Fresh[53]), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U36 ( .A(Fresh[52]), .B(
        SubCellInst_SboxInst_8_Q4), .Z(
        SubCellInst_SboxInst_8_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U35 ( .A(new_AGEMA_signal_1843), .B(
        Fresh[53]), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U34 ( .A(Fresh[51]), .B(
        SubCellInst_SboxInst_8_Q4), .Z(
        SubCellInst_SboxInst_8_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U33 ( .A(Fresh[52]), .B(
        new_AGEMA_signal_1843), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U32 ( .A(new_AGEMA_signal_1842), .B(
        Fresh[51]), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U25 ( .A1(Ciphertext_s2[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U24 ( .A1(Ciphertext_s2[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U23 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND3_U1_U22 ( .A(Fresh[53]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U21 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND3_U1_U19 ( .A(Fresh[52]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND3_U1_U17 ( .A(Fresh[51]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U16 ( .A1(new_AGEMA_signal_1843), 
        .A2(Ciphertext_s2[34]), .ZN(SubCellInst_SboxInst_8_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U15 ( .A1(new_AGEMA_signal_1842), 
        .A2(Ciphertext_s1[34]), .ZN(SubCellInst_SboxInst_8_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_8_Q4), 
        .A2(SubCellInst_SboxInst_8_n3), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND3_U1_n33), .Z(new_AGEMA_signal_1983) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n32), .B(
        SubCellInst_SboxInst_8_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_8_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND3_U1_n30), .Z(new_AGEMA_signal_1982) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n29), .B(
        SubCellInst_SboxInst_8_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_8_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND3_U1_n27), .Z(SubCellInst_SboxInst_8_T2) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n26), .B(
        SubCellInst_SboxInst_8_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_8_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3671), 
        .B(SubCellInst_SboxInst_8_T2), .Z(SubCellInst_SboxInst_8_Q7) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3673), 
        .B(new_AGEMA_signal_1982), .Z(new_AGEMA_signal_2094) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3675), 
        .B(new_AGEMA_signal_1983), .Z(new_AGEMA_signal_2095) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3677), 
        .B(SubCellInst_SboxInst_8_T0), .Z(SubCellInst_SboxInst_8_L3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3679), 
        .B(new_AGEMA_signal_1980), .Z(new_AGEMA_signal_2096) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3681), 
        .B(new_AGEMA_signal_1981), .Z(new_AGEMA_signal_2097) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L3), .B(SubCellInst_SboxInst_8_T2), .Z(
        SubCellInst_SboxInst_8_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2096), 
        .B(new_AGEMA_signal_1982), .Z(new_AGEMA_signal_2316) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2097), 
        .B(new_AGEMA_signal_1983), .Z(new_AGEMA_signal_2317) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3683), 
        .B(SubCellInst_SboxInst_8_T2), .Z(SubCellInst_SboxInst_8_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3685), 
        .B(new_AGEMA_signal_1982), .Z(new_AGEMA_signal_2220) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3687), 
        .B(new_AGEMA_signal_1983), .Z(new_AGEMA_signal_2221) );
  INV_X1 SubCellInst_SboxInst_9_U3_U1 ( .A(SubCellInst_SboxInst_9_YY_1_), .ZN(
        AddRoundConstantOutput[39]) );
  INV_X1 SubCellInst_SboxInst_9_U2_U1 ( .A(SubCellInst_SboxInst_9_YY_0_), .ZN(
        AddRoundConstantOutput[38]) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U37 ( .A(new_AGEMA_signal_1852), .B(
        Fresh[56]), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U36 ( .A(Fresh[55]), .B(
        SubCellInst_SboxInst_9_Q1), .Z(
        SubCellInst_SboxInst_9_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U35 ( .A(new_AGEMA_signal_1853), .B(
        Fresh[56]), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U34 ( .A(Fresh[54]), .B(
        SubCellInst_SboxInst_9_Q1), .Z(
        SubCellInst_SboxInst_9_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U33 ( .A(Fresh[55]), .B(
        new_AGEMA_signal_1853), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U32 ( .A(new_AGEMA_signal_1852), .B(
        Fresh[54]), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U25 ( .A1(Ciphertext_s2[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U24 ( .A1(Ciphertext_s2[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U23 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND1_U1_U22 ( .A(Fresh[56]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U21 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND1_U1_U19 ( .A(Fresh[55]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND1_U1_U17 ( .A(Fresh[54]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U16 ( .A1(new_AGEMA_signal_1853), 
        .A2(Ciphertext_s2[38]), .ZN(SubCellInst_SboxInst_9_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U15 ( .A1(new_AGEMA_signal_1852), 
        .A2(Ciphertext_s1[38]), .ZN(SubCellInst_SboxInst_9_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_9_Q1), 
        .A2(SubCellInst_SboxInst_9_n3), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND1_U1_n33), .Z(new_AGEMA_signal_1987) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n32), .B(
        SubCellInst_SboxInst_9_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_9_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND1_U1_n30), .Z(new_AGEMA_signal_1986) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n29), .B(
        SubCellInst_SboxInst_9_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_9_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND1_U1_n27), .Z(SubCellInst_SboxInst_9_T0) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n26), .B(
        SubCellInst_SboxInst_9_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_9_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3689), 
        .B(SubCellInst_SboxInst_9_T0), .Z(SubCellInst_SboxInst_9_Q2) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3691), 
        .B(new_AGEMA_signal_1986), .Z(new_AGEMA_signal_2100) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3693), 
        .B(new_AGEMA_signal_1987), .Z(new_AGEMA_signal_2101) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U37 ( .A(new_AGEMA_signal_1854), .B(
        Fresh[59]), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U36 ( .A(Fresh[58]), .B(
        SubCellInst_SboxInst_9_Q4), .Z(
        SubCellInst_SboxInst_9_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U35 ( .A(new_AGEMA_signal_1855), .B(
        Fresh[59]), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U34 ( .A(Fresh[57]), .B(
        SubCellInst_SboxInst_9_Q4), .Z(
        SubCellInst_SboxInst_9_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U33 ( .A(Fresh[58]), .B(
        new_AGEMA_signal_1855), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U32 ( .A(new_AGEMA_signal_1854), .B(
        Fresh[57]), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U25 ( .A1(Ciphertext_s2[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U24 ( .A1(Ciphertext_s2[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U23 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND3_U1_U22 ( .A(Fresh[59]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U21 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND3_U1_U19 ( .A(Fresh[58]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND3_U1_U17 ( .A(Fresh[57]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U16 ( .A1(new_AGEMA_signal_1855), 
        .A2(Ciphertext_s2[38]), .ZN(SubCellInst_SboxInst_9_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U15 ( .A1(new_AGEMA_signal_1854), 
        .A2(Ciphertext_s1[38]), .ZN(SubCellInst_SboxInst_9_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_9_Q4), 
        .A2(SubCellInst_SboxInst_9_n3), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND3_U1_n33), .Z(new_AGEMA_signal_1989) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n32), .B(
        SubCellInst_SboxInst_9_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_9_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND3_U1_n30), .Z(new_AGEMA_signal_1988) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n29), .B(
        SubCellInst_SboxInst_9_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_9_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND3_U1_n27), .Z(SubCellInst_SboxInst_9_T2) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n26), .B(
        SubCellInst_SboxInst_9_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_9_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3695), 
        .B(SubCellInst_SboxInst_9_T2), .Z(SubCellInst_SboxInst_9_Q7) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3697), 
        .B(new_AGEMA_signal_1988), .Z(new_AGEMA_signal_2102) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3699), 
        .B(new_AGEMA_signal_1989), .Z(new_AGEMA_signal_2103) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3701), 
        .B(SubCellInst_SboxInst_9_T0), .Z(SubCellInst_SboxInst_9_L3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3703), 
        .B(new_AGEMA_signal_1986), .Z(new_AGEMA_signal_2104) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3705), 
        .B(new_AGEMA_signal_1987), .Z(new_AGEMA_signal_2105) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L3), .B(SubCellInst_SboxInst_9_T2), .Z(
        SubCellInst_SboxInst_9_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2104), 
        .B(new_AGEMA_signal_1988), .Z(new_AGEMA_signal_2320) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2105), 
        .B(new_AGEMA_signal_1989), .Z(new_AGEMA_signal_2321) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3707), 
        .B(SubCellInst_SboxInst_9_T2), .Z(SubCellInst_SboxInst_9_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3709), 
        .B(new_AGEMA_signal_1988), .Z(new_AGEMA_signal_2228) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3711), 
        .B(new_AGEMA_signal_1989), .Z(new_AGEMA_signal_2229) );
  INV_X1 SubCellInst_SboxInst_10_U3_U1 ( .A(SubCellInst_SboxInst_10_YY_1_), 
        .ZN(AddRoundConstantOutput[43]) );
  INV_X1 SubCellInst_SboxInst_10_U2_U1 ( .A(SubCellInst_SboxInst_10_YY_0_), 
        .ZN(AddRoundConstantOutput[42]) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U37 ( .A(new_AGEMA_signal_1864), .B(
        Fresh[62]), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U36 ( .A(Fresh[61]), .B(
        SubCellInst_SboxInst_10_Q1), .Z(
        SubCellInst_SboxInst_10_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U35 ( .A(new_AGEMA_signal_1865), .B(
        Fresh[62]), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U34 ( .A(Fresh[60]), .B(
        SubCellInst_SboxInst_10_Q1), .Z(
        SubCellInst_SboxInst_10_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U33 ( .A(Fresh[61]), .B(
        new_AGEMA_signal_1865), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U32 ( .A(new_AGEMA_signal_1864), .B(
        Fresh[60]), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U25 ( .A1(Ciphertext_s2[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U24 ( .A1(Ciphertext_s2[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U23 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND1_U1_U22 ( .A(Fresh[62]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U21 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_10_n3), .A2(SubCellInst_SboxInst_10_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND1_U1_U19 ( .A(Fresh[61]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_10_n3), .A2(SubCellInst_SboxInst_10_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND1_U1_U17 ( .A(Fresh[60]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U16 ( .A1(new_AGEMA_signal_1865), 
        .A2(Ciphertext_s2[42]), .ZN(SubCellInst_SboxInst_10_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U15 ( .A1(new_AGEMA_signal_1864), 
        .A2(Ciphertext_s1[42]), .ZN(SubCellInst_SboxInst_10_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_10_Q1), .A2(SubCellInst_SboxInst_10_n3), .ZN(SubCellInst_SboxInst_10_AND1_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND1_U1_n33), .Z(new_AGEMA_signal_1993) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n32), .B(
        SubCellInst_SboxInst_10_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_10_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND1_U1_n30), .Z(new_AGEMA_signal_1992) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n29), .B(
        SubCellInst_SboxInst_10_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_10_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND1_U1_n27), .Z(SubCellInst_SboxInst_10_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n26), .B(
        SubCellInst_SboxInst_10_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_10_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3713), 
        .B(SubCellInst_SboxInst_10_T0), .Z(SubCellInst_SboxInst_10_Q2) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3715), 
        .B(new_AGEMA_signal_1992), .Z(new_AGEMA_signal_2108) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3717), 
        .B(new_AGEMA_signal_1993), .Z(new_AGEMA_signal_2109) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U37 ( .A(new_AGEMA_signal_1866), .B(
        Fresh[65]), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U36 ( .A(Fresh[64]), .B(
        SubCellInst_SboxInst_10_Q4), .Z(
        SubCellInst_SboxInst_10_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U35 ( .A(new_AGEMA_signal_1867), .B(
        Fresh[65]), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U34 ( .A(Fresh[63]), .B(
        SubCellInst_SboxInst_10_Q4), .Z(
        SubCellInst_SboxInst_10_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U33 ( .A(Fresh[64]), .B(
        new_AGEMA_signal_1867), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U32 ( .A(new_AGEMA_signal_1866), .B(
        Fresh[63]), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U25 ( .A1(Ciphertext_s2[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U24 ( .A1(Ciphertext_s2[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U23 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND3_U1_U22 ( .A(Fresh[65]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U21 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_10_n3), .A2(SubCellInst_SboxInst_10_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND3_U1_U19 ( .A(Fresh[64]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_10_n3), .A2(SubCellInst_SboxInst_10_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND3_U1_U17 ( .A(Fresh[63]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U16 ( .A1(new_AGEMA_signal_1867), 
        .A2(Ciphertext_s2[42]), .ZN(SubCellInst_SboxInst_10_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U15 ( .A1(new_AGEMA_signal_1866), 
        .A2(Ciphertext_s1[42]), .ZN(SubCellInst_SboxInst_10_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_10_Q4), .A2(SubCellInst_SboxInst_10_n3), .ZN(SubCellInst_SboxInst_10_AND3_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND3_U1_n33), .Z(new_AGEMA_signal_1995) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n32), .B(
        SubCellInst_SboxInst_10_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_10_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND3_U1_n30), .Z(new_AGEMA_signal_1994) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n29), .B(
        SubCellInst_SboxInst_10_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_10_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND3_U1_n27), .Z(SubCellInst_SboxInst_10_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n26), .B(
        SubCellInst_SboxInst_10_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_10_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3719), 
        .B(SubCellInst_SboxInst_10_T2), .Z(SubCellInst_SboxInst_10_Q7) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3721), 
        .B(new_AGEMA_signal_1994), .Z(new_AGEMA_signal_2110) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3723), 
        .B(new_AGEMA_signal_1995), .Z(new_AGEMA_signal_2111) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3725), .B(SubCellInst_SboxInst_10_T0), .Z(SubCellInst_SboxInst_10_L3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3727), .B(new_AGEMA_signal_1992), .Z(new_AGEMA_signal_2112) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3729), .B(new_AGEMA_signal_1993), .Z(new_AGEMA_signal_2113) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L3), .B(SubCellInst_SboxInst_10_T2), .Z(
        SubCellInst_SboxInst_10_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2112), .B(new_AGEMA_signal_1994), .Z(new_AGEMA_signal_2324) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2113), .B(new_AGEMA_signal_1995), .Z(new_AGEMA_signal_2325) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3731), .B(SubCellInst_SboxInst_10_T2), .Z(SubCellInst_SboxInst_10_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3733), .B(new_AGEMA_signal_1994), .Z(new_AGEMA_signal_2236) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3735), .B(new_AGEMA_signal_1995), .Z(new_AGEMA_signal_2237) );
  INV_X1 SubCellInst_SboxInst_11_U3_U1 ( .A(SubCellInst_SboxInst_11_YY_1_), 
        .ZN(SubCellOutput_47) );
  INV_X1 SubCellInst_SboxInst_11_U2_U1 ( .A(SubCellInst_SboxInst_11_YY_0_), 
        .ZN(SubCellOutput_46) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U37 ( .A(new_AGEMA_signal_1876), .B(
        Fresh[68]), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U36 ( .A(Fresh[67]), .B(
        SubCellInst_SboxInst_11_Q1), .Z(
        SubCellInst_SboxInst_11_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U35 ( .A(new_AGEMA_signal_1877), .B(
        Fresh[68]), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U34 ( .A(Fresh[66]), .B(
        SubCellInst_SboxInst_11_Q1), .Z(
        SubCellInst_SboxInst_11_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U33 ( .A(Fresh[67]), .B(
        new_AGEMA_signal_1877), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U32 ( .A(new_AGEMA_signal_1876), .B(
        Fresh[66]), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U25 ( .A1(Ciphertext_s2[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U24 ( .A1(Ciphertext_s2[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U23 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND1_U1_U22 ( .A(Fresh[68]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U21 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_11_n3), .A2(SubCellInst_SboxInst_11_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND1_U1_U19 ( .A(Fresh[67]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_11_n3), .A2(SubCellInst_SboxInst_11_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND1_U1_U17 ( .A(Fresh[66]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U16 ( .A1(new_AGEMA_signal_1877), 
        .A2(Ciphertext_s2[46]), .ZN(SubCellInst_SboxInst_11_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U15 ( .A1(new_AGEMA_signal_1876), 
        .A2(Ciphertext_s1[46]), .ZN(SubCellInst_SboxInst_11_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_11_Q1), .A2(SubCellInst_SboxInst_11_n3), .ZN(SubCellInst_SboxInst_11_AND1_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND1_U1_n33), .Z(new_AGEMA_signal_1999) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n32), .B(
        SubCellInst_SboxInst_11_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_11_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND1_U1_n30), .Z(new_AGEMA_signal_1998) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n29), .B(
        SubCellInst_SboxInst_11_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_11_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND1_U1_n27), .Z(SubCellInst_SboxInst_11_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n26), .B(
        SubCellInst_SboxInst_11_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_11_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3737), 
        .B(SubCellInst_SboxInst_11_T0), .Z(SubCellInst_SboxInst_11_Q2) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3739), 
        .B(new_AGEMA_signal_1998), .Z(new_AGEMA_signal_2116) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3741), 
        .B(new_AGEMA_signal_1999), .Z(new_AGEMA_signal_2117) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U37 ( .A(new_AGEMA_signal_1878), .B(
        Fresh[71]), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U36 ( .A(Fresh[70]), .B(
        SubCellInst_SboxInst_11_Q4), .Z(
        SubCellInst_SboxInst_11_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U35 ( .A(new_AGEMA_signal_1879), .B(
        Fresh[71]), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U34 ( .A(Fresh[69]), .B(
        SubCellInst_SboxInst_11_Q4), .Z(
        SubCellInst_SboxInst_11_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U33 ( .A(Fresh[70]), .B(
        new_AGEMA_signal_1879), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U32 ( .A(new_AGEMA_signal_1878), .B(
        Fresh[69]), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U25 ( .A1(Ciphertext_s2[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U24 ( .A1(Ciphertext_s2[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U23 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND3_U1_U22 ( .A(Fresh[71]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U21 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_11_n3), .A2(SubCellInst_SboxInst_11_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND3_U1_U19 ( .A(Fresh[70]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_11_n3), .A2(SubCellInst_SboxInst_11_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND3_U1_U17 ( .A(Fresh[69]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U16 ( .A1(new_AGEMA_signal_1879), 
        .A2(Ciphertext_s2[46]), .ZN(SubCellInst_SboxInst_11_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U15 ( .A1(new_AGEMA_signal_1878), 
        .A2(Ciphertext_s1[46]), .ZN(SubCellInst_SboxInst_11_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_11_Q4), .A2(SubCellInst_SboxInst_11_n3), .ZN(SubCellInst_SboxInst_11_AND3_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND3_U1_n33), .Z(new_AGEMA_signal_2001) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n32), .B(
        SubCellInst_SboxInst_11_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_11_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND3_U1_n30), .Z(new_AGEMA_signal_2000) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n29), .B(
        SubCellInst_SboxInst_11_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_11_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND3_U1_n27), .Z(SubCellInst_SboxInst_11_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n26), .B(
        SubCellInst_SboxInst_11_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_11_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3743), 
        .B(SubCellInst_SboxInst_11_T2), .Z(SubCellInst_SboxInst_11_Q7) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3745), 
        .B(new_AGEMA_signal_2000), .Z(new_AGEMA_signal_2118) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3747), 
        .B(new_AGEMA_signal_2001), .Z(new_AGEMA_signal_2119) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3749), .B(SubCellInst_SboxInst_11_T0), .Z(SubCellInst_SboxInst_11_L3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3751), .B(new_AGEMA_signal_1998), .Z(new_AGEMA_signal_2120) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3753), .B(new_AGEMA_signal_1999), .Z(new_AGEMA_signal_2121) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L3), .B(SubCellInst_SboxInst_11_T2), .Z(
        SubCellInst_SboxInst_11_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2120), .B(new_AGEMA_signal_2000), .Z(new_AGEMA_signal_2328) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2121), .B(new_AGEMA_signal_2001), .Z(new_AGEMA_signal_2329) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3755), .B(SubCellInst_SboxInst_11_T2), .Z(SubCellInst_SboxInst_11_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3757), .B(new_AGEMA_signal_2000), .Z(new_AGEMA_signal_2244) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3759), .B(new_AGEMA_signal_2001), .Z(new_AGEMA_signal_2245) );
  INV_X1 SubCellInst_SboxInst_12_U3_U1 ( .A(SubCellInst_SboxInst_12_YY_1_), 
        .ZN(AddRoundConstantOutput[51]) );
  INV_X1 SubCellInst_SboxInst_12_U2_U1 ( .A(SubCellInst_SboxInst_12_YY_0_), 
        .ZN(AddRoundConstantOutput[50]) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U37 ( .A(new_AGEMA_signal_1888), .B(
        Fresh[74]), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U36 ( .A(Fresh[73]), .B(
        SubCellInst_SboxInst_12_Q1), .Z(
        SubCellInst_SboxInst_12_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U35 ( .A(new_AGEMA_signal_1889), .B(
        Fresh[74]), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U34 ( .A(Fresh[72]), .B(
        SubCellInst_SboxInst_12_Q1), .Z(
        SubCellInst_SboxInst_12_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U33 ( .A(Fresh[73]), .B(
        new_AGEMA_signal_1889), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U32 ( .A(new_AGEMA_signal_1888), .B(
        Fresh[72]), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U25 ( .A1(Ciphertext_s2[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U24 ( .A1(Ciphertext_s2[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U23 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND1_U1_U22 ( .A(Fresh[74]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U21 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_12_n3), .A2(SubCellInst_SboxInst_12_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND1_U1_U19 ( .A(Fresh[73]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_12_n3), .A2(SubCellInst_SboxInst_12_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND1_U1_U17 ( .A(Fresh[72]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U16 ( .A1(new_AGEMA_signal_1889), 
        .A2(Ciphertext_s2[50]), .ZN(SubCellInst_SboxInst_12_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U15 ( .A1(new_AGEMA_signal_1888), 
        .A2(Ciphertext_s1[50]), .ZN(SubCellInst_SboxInst_12_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_12_Q1), .A2(SubCellInst_SboxInst_12_n3), .ZN(SubCellInst_SboxInst_12_AND1_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND1_U1_n33), .Z(new_AGEMA_signal_2005) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n32), .B(
        SubCellInst_SboxInst_12_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_12_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND1_U1_n30), .Z(new_AGEMA_signal_2004) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n29), .B(
        SubCellInst_SboxInst_12_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_12_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND1_U1_n27), .Z(SubCellInst_SboxInst_12_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n26), .B(
        SubCellInst_SboxInst_12_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_12_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3761), 
        .B(SubCellInst_SboxInst_12_T0), .Z(SubCellInst_SboxInst_12_Q2) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3763), 
        .B(new_AGEMA_signal_2004), .Z(new_AGEMA_signal_2124) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3765), 
        .B(new_AGEMA_signal_2005), .Z(new_AGEMA_signal_2125) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U37 ( .A(new_AGEMA_signal_1890), .B(
        Fresh[77]), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U36 ( .A(Fresh[76]), .B(
        SubCellInst_SboxInst_12_Q4), .Z(
        SubCellInst_SboxInst_12_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U35 ( .A(new_AGEMA_signal_1891), .B(
        Fresh[77]), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U34 ( .A(Fresh[75]), .B(
        SubCellInst_SboxInst_12_Q4), .Z(
        SubCellInst_SboxInst_12_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U33 ( .A(Fresh[76]), .B(
        new_AGEMA_signal_1891), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U32 ( .A(new_AGEMA_signal_1890), .B(
        Fresh[75]), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U25 ( .A1(Ciphertext_s2[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U24 ( .A1(Ciphertext_s2[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U23 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND3_U1_U22 ( .A(Fresh[77]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U21 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_12_n3), .A2(SubCellInst_SboxInst_12_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND3_U1_U19 ( .A(Fresh[76]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_12_n3), .A2(SubCellInst_SboxInst_12_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND3_U1_U17 ( .A(Fresh[75]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U16 ( .A1(new_AGEMA_signal_1891), 
        .A2(Ciphertext_s2[50]), .ZN(SubCellInst_SboxInst_12_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U15 ( .A1(new_AGEMA_signal_1890), 
        .A2(Ciphertext_s1[50]), .ZN(SubCellInst_SboxInst_12_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_12_Q4), .A2(SubCellInst_SboxInst_12_n3), .ZN(SubCellInst_SboxInst_12_AND3_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND3_U1_n33), .Z(new_AGEMA_signal_2007) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n32), .B(
        SubCellInst_SboxInst_12_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_12_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND3_U1_n30), .Z(new_AGEMA_signal_2006) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n29), .B(
        SubCellInst_SboxInst_12_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_12_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND3_U1_n27), .Z(SubCellInst_SboxInst_12_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n26), .B(
        SubCellInst_SboxInst_12_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_12_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3767), 
        .B(SubCellInst_SboxInst_12_T2), .Z(SubCellInst_SboxInst_12_Q7) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3769), 
        .B(new_AGEMA_signal_2006), .Z(new_AGEMA_signal_2126) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3771), 
        .B(new_AGEMA_signal_2007), .Z(new_AGEMA_signal_2127) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3773), .B(SubCellInst_SboxInst_12_T0), .Z(SubCellInst_SboxInst_12_L3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3775), .B(new_AGEMA_signal_2004), .Z(new_AGEMA_signal_2128) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3777), .B(new_AGEMA_signal_2005), .Z(new_AGEMA_signal_2129) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L3), .B(SubCellInst_SboxInst_12_T2), .Z(
        SubCellInst_SboxInst_12_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2128), .B(new_AGEMA_signal_2006), .Z(new_AGEMA_signal_2332) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2129), .B(new_AGEMA_signal_2007), .Z(new_AGEMA_signal_2333) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3779), .B(SubCellInst_SboxInst_12_T2), .Z(SubCellInst_SboxInst_12_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3781), .B(new_AGEMA_signal_2006), .Z(new_AGEMA_signal_2252) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3783), .B(new_AGEMA_signal_2007), .Z(new_AGEMA_signal_2253) );
  INV_X1 SubCellInst_SboxInst_13_U3_U1 ( .A(SubCellInst_SboxInst_13_YY_1_), 
        .ZN(AddRoundConstantOutput[55]) );
  INV_X1 SubCellInst_SboxInst_13_U2_U1 ( .A(SubCellInst_SboxInst_13_YY_0_), 
        .ZN(AddRoundConstantOutput[54]) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U37 ( .A(new_AGEMA_signal_1900), .B(
        Fresh[80]), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U36 ( .A(Fresh[79]), .B(
        SubCellInst_SboxInst_13_Q1), .Z(
        SubCellInst_SboxInst_13_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U35 ( .A(new_AGEMA_signal_1901), .B(
        Fresh[80]), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U34 ( .A(Fresh[78]), .B(
        SubCellInst_SboxInst_13_Q1), .Z(
        SubCellInst_SboxInst_13_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U33 ( .A(Fresh[79]), .B(
        new_AGEMA_signal_1901), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U32 ( .A(new_AGEMA_signal_1900), .B(
        Fresh[78]), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U25 ( .A1(Ciphertext_s2[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U24 ( .A1(Ciphertext_s2[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U23 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND1_U1_U22 ( .A(Fresh[80]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U21 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_13_n3), .A2(SubCellInst_SboxInst_13_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND1_U1_U19 ( .A(Fresh[79]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_13_n3), .A2(SubCellInst_SboxInst_13_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND1_U1_U17 ( .A(Fresh[78]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U16 ( .A1(new_AGEMA_signal_1901), 
        .A2(Ciphertext_s2[54]), .ZN(SubCellInst_SboxInst_13_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U15 ( .A1(new_AGEMA_signal_1900), 
        .A2(Ciphertext_s1[54]), .ZN(SubCellInst_SboxInst_13_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_13_Q1), .A2(SubCellInst_SboxInst_13_n3), .ZN(SubCellInst_SboxInst_13_AND1_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND1_U1_n33), .Z(new_AGEMA_signal_2011) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n32), .B(
        SubCellInst_SboxInst_13_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_13_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND1_U1_n30), .Z(new_AGEMA_signal_2010) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n29), .B(
        SubCellInst_SboxInst_13_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_13_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND1_U1_n27), .Z(SubCellInst_SboxInst_13_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n26), .B(
        SubCellInst_SboxInst_13_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_13_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3785), 
        .B(SubCellInst_SboxInst_13_T0), .Z(SubCellInst_SboxInst_13_Q2) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3787), 
        .B(new_AGEMA_signal_2010), .Z(new_AGEMA_signal_2132) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3789), 
        .B(new_AGEMA_signal_2011), .Z(new_AGEMA_signal_2133) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U37 ( .A(new_AGEMA_signal_1902), .B(
        Fresh[83]), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U36 ( .A(Fresh[82]), .B(
        SubCellInst_SboxInst_13_Q4), .Z(
        SubCellInst_SboxInst_13_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U35 ( .A(new_AGEMA_signal_1903), .B(
        Fresh[83]), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U34 ( .A(Fresh[81]), .B(
        SubCellInst_SboxInst_13_Q4), .Z(
        SubCellInst_SboxInst_13_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U33 ( .A(Fresh[82]), .B(
        new_AGEMA_signal_1903), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U32 ( .A(new_AGEMA_signal_1902), .B(
        Fresh[81]), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U25 ( .A1(Ciphertext_s2[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U24 ( .A1(Ciphertext_s2[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U23 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND3_U1_U22 ( .A(Fresh[83]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U21 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_13_n3), .A2(SubCellInst_SboxInst_13_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND3_U1_U19 ( .A(Fresh[82]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_13_n3), .A2(SubCellInst_SboxInst_13_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND3_U1_U17 ( .A(Fresh[81]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U16 ( .A1(new_AGEMA_signal_1903), 
        .A2(Ciphertext_s2[54]), .ZN(SubCellInst_SboxInst_13_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U15 ( .A1(new_AGEMA_signal_1902), 
        .A2(Ciphertext_s1[54]), .ZN(SubCellInst_SboxInst_13_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_13_Q4), .A2(SubCellInst_SboxInst_13_n3), .ZN(SubCellInst_SboxInst_13_AND3_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND3_U1_n33), .Z(new_AGEMA_signal_2013) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n32), .B(
        SubCellInst_SboxInst_13_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_13_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND3_U1_n30), .Z(new_AGEMA_signal_2012) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n29), .B(
        SubCellInst_SboxInst_13_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_13_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND3_U1_n27), .Z(SubCellInst_SboxInst_13_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n26), .B(
        SubCellInst_SboxInst_13_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_13_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3791), 
        .B(SubCellInst_SboxInst_13_T2), .Z(SubCellInst_SboxInst_13_Q7) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3793), 
        .B(new_AGEMA_signal_2012), .Z(new_AGEMA_signal_2134) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3795), 
        .B(new_AGEMA_signal_2013), .Z(new_AGEMA_signal_2135) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3797), .B(SubCellInst_SboxInst_13_T0), .Z(SubCellInst_SboxInst_13_L3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3799), .B(new_AGEMA_signal_2010), .Z(new_AGEMA_signal_2136) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3801), .B(new_AGEMA_signal_2011), .Z(new_AGEMA_signal_2137) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L3), .B(SubCellInst_SboxInst_13_T2), .Z(
        SubCellInst_SboxInst_13_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2136), .B(new_AGEMA_signal_2012), .Z(new_AGEMA_signal_2336) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2137), .B(new_AGEMA_signal_2013), .Z(new_AGEMA_signal_2337) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3803), .B(SubCellInst_SboxInst_13_T2), .Z(SubCellInst_SboxInst_13_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3805), .B(new_AGEMA_signal_2012), .Z(new_AGEMA_signal_2260) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3807), .B(new_AGEMA_signal_2013), .Z(new_AGEMA_signal_2261) );
  INV_X1 SubCellInst_SboxInst_14_U3_U1 ( .A(SubCellInst_SboxInst_14_YY_1_), 
        .ZN(AddRoundConstantOutput[59]) );
  INV_X1 SubCellInst_SboxInst_14_U2_U1 ( .A(SubCellInst_SboxInst_14_YY_0_), 
        .ZN(AddRoundConstantOutput[58]) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U37 ( .A(new_AGEMA_signal_1912), .B(
        Fresh[86]), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U36 ( .A(Fresh[85]), .B(
        SubCellInst_SboxInst_14_Q1), .Z(
        SubCellInst_SboxInst_14_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U35 ( .A(new_AGEMA_signal_1913), .B(
        Fresh[86]), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U34 ( .A(Fresh[84]), .B(
        SubCellInst_SboxInst_14_Q1), .Z(
        SubCellInst_SboxInst_14_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U33 ( .A(Fresh[85]), .B(
        new_AGEMA_signal_1913), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U32 ( .A(new_AGEMA_signal_1912), .B(
        Fresh[84]), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U25 ( .A1(Ciphertext_s2[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U24 ( .A1(Ciphertext_s2[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U23 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND1_U1_U22 ( .A(Fresh[86]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U21 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_14_n3), .A2(SubCellInst_SboxInst_14_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND1_U1_U19 ( .A(Fresh[85]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_14_n3), .A2(SubCellInst_SboxInst_14_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND1_U1_U17 ( .A(Fresh[84]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U16 ( .A1(new_AGEMA_signal_1913), 
        .A2(Ciphertext_s2[58]), .ZN(SubCellInst_SboxInst_14_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U15 ( .A1(new_AGEMA_signal_1912), 
        .A2(Ciphertext_s1[58]), .ZN(SubCellInst_SboxInst_14_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_14_Q1), .A2(SubCellInst_SboxInst_14_n3), .ZN(SubCellInst_SboxInst_14_AND1_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND1_U1_n33), .Z(new_AGEMA_signal_2017) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n32), .B(
        SubCellInst_SboxInst_14_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_14_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND1_U1_n30), .Z(new_AGEMA_signal_2016) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n29), .B(
        SubCellInst_SboxInst_14_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_14_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND1_U1_n27), .Z(SubCellInst_SboxInst_14_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n26), .B(
        SubCellInst_SboxInst_14_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_14_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3809), 
        .B(SubCellInst_SboxInst_14_T0), .Z(SubCellInst_SboxInst_14_Q2) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3811), 
        .B(new_AGEMA_signal_2016), .Z(new_AGEMA_signal_2140) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3813), 
        .B(new_AGEMA_signal_2017), .Z(new_AGEMA_signal_2141) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U37 ( .A(new_AGEMA_signal_1914), .B(
        Fresh[89]), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U36 ( .A(Fresh[88]), .B(
        SubCellInst_SboxInst_14_Q4), .Z(
        SubCellInst_SboxInst_14_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U35 ( .A(new_AGEMA_signal_1915), .B(
        Fresh[89]), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U34 ( .A(Fresh[87]), .B(
        SubCellInst_SboxInst_14_Q4), .Z(
        SubCellInst_SboxInst_14_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U33 ( .A(Fresh[88]), .B(
        new_AGEMA_signal_1915), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U32 ( .A(new_AGEMA_signal_1914), .B(
        Fresh[87]), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U25 ( .A1(Ciphertext_s2[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U24 ( .A1(Ciphertext_s2[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U23 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND3_U1_U22 ( .A(Fresh[89]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U21 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_14_n3), .A2(SubCellInst_SboxInst_14_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND3_U1_U19 ( .A(Fresh[88]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_14_n3), .A2(SubCellInst_SboxInst_14_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND3_U1_U17 ( .A(Fresh[87]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U16 ( .A1(new_AGEMA_signal_1915), 
        .A2(Ciphertext_s2[58]), .ZN(SubCellInst_SboxInst_14_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U15 ( .A1(new_AGEMA_signal_1914), 
        .A2(Ciphertext_s1[58]), .ZN(SubCellInst_SboxInst_14_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_14_Q4), .A2(SubCellInst_SboxInst_14_n3), .ZN(SubCellInst_SboxInst_14_AND3_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND3_U1_n33), .Z(new_AGEMA_signal_2019) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n32), .B(
        SubCellInst_SboxInst_14_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_14_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND3_U1_n30), .Z(new_AGEMA_signal_2018) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n29), .B(
        SubCellInst_SboxInst_14_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_14_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND3_U1_n27), .Z(SubCellInst_SboxInst_14_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n26), .B(
        SubCellInst_SboxInst_14_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_14_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3815), 
        .B(SubCellInst_SboxInst_14_T2), .Z(SubCellInst_SboxInst_14_Q7) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3817), 
        .B(new_AGEMA_signal_2018), .Z(new_AGEMA_signal_2142) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3819), 
        .B(new_AGEMA_signal_2019), .Z(new_AGEMA_signal_2143) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3821), .B(SubCellInst_SboxInst_14_T0), .Z(SubCellInst_SboxInst_14_L3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3823), .B(new_AGEMA_signal_2016), .Z(new_AGEMA_signal_2144) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3825), .B(new_AGEMA_signal_2017), .Z(new_AGEMA_signal_2145) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L3), .B(SubCellInst_SboxInst_14_T2), .Z(
        SubCellInst_SboxInst_14_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2144), .B(new_AGEMA_signal_2018), .Z(new_AGEMA_signal_2340) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2145), .B(new_AGEMA_signal_2019), .Z(new_AGEMA_signal_2341) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3827), .B(SubCellInst_SboxInst_14_T2), .Z(SubCellInst_SboxInst_14_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3829), .B(new_AGEMA_signal_2018), .Z(new_AGEMA_signal_2268) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3831), .B(new_AGEMA_signal_2019), .Z(new_AGEMA_signal_2269) );
  INV_X1 SubCellInst_SboxInst_15_U3_U1 ( .A(SubCellInst_SboxInst_15_YY_1_), 
        .ZN(SubCellOutput[63]) );
  INV_X1 SubCellInst_SboxInst_15_U2_U1 ( .A(SubCellInst_SboxInst_15_YY_0_), 
        .ZN(SubCellOutput[62]) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U37 ( .A(new_AGEMA_signal_1924), .B(
        Fresh[92]), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U36 ( .A(Fresh[91]), .B(
        SubCellInst_SboxInst_15_Q1), .Z(
        SubCellInst_SboxInst_15_AND1_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U35 ( .A(new_AGEMA_signal_1925), .B(
        Fresh[92]), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U34 ( .A(Fresh[90]), .B(
        SubCellInst_SboxInst_15_Q1), .Z(
        SubCellInst_SboxInst_15_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U33 ( .A(Fresh[91]), .B(
        new_AGEMA_signal_1925), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U32 ( .A(new_AGEMA_signal_1924), .B(
        Fresh[90]), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U31 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U30 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U29 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U28 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U27 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U26 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U25 ( .A1(Ciphertext_s2[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U24 ( .A1(Ciphertext_s2[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U23 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n36), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND1_U1_U22 ( .A(Fresh[92]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U21 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U20 ( .A1(SubCellInst_SboxInst_15_n3), .A2(SubCellInst_SboxInst_15_AND1_U1_n35), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND1_U1_U19 ( .A(Fresh[91]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U18 ( .A1(SubCellInst_SboxInst_15_n3), .A2(SubCellInst_SboxInst_15_AND1_U1_n34), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND1_U1_U17 ( .A(Fresh[90]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U16 ( .A1(new_AGEMA_signal_1925), 
        .A2(Ciphertext_s2[62]), .ZN(SubCellInst_SboxInst_15_AND1_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U15 ( .A1(new_AGEMA_signal_1924), 
        .A2(Ciphertext_s1[62]), .ZN(SubCellInst_SboxInst_15_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U14 ( .A1(SubCellInst_SboxInst_15_Q1), .A2(SubCellInst_SboxInst_15_n3), .ZN(SubCellInst_SboxInst_15_AND1_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U13 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND1_U1_n33), .Z(new_AGEMA_signal_2023) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U12 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n32), .B(
        SubCellInst_SboxInst_15_AND1_U1_n31), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U11 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND1_U1_z[2]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U10 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_15_AND1_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U9 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND1_U1_n30), .Z(new_AGEMA_signal_2022) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U8 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n29), .B(
        SubCellInst_SboxInst_15_AND1_U1_n28), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U7 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND1_U1_z[1]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U6 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_15_AND1_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND1_U1_n27), .Z(SubCellInst_SboxInst_15_T0)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n26), .B(
        SubCellInst_SboxInst_15_AND1_U1_n25), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND1_U1_z[0]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_15_AND1_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR2_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3833), 
        .B(SubCellInst_SboxInst_15_T0), .Z(SubCellInst_SboxInst_15_Q2) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3835), 
        .B(new_AGEMA_signal_2022), .Z(new_AGEMA_signal_2148) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR2_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3837), 
        .B(new_AGEMA_signal_2023), .Z(new_AGEMA_signal_2149) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U37 ( .A(new_AGEMA_signal_1926), .B(
        Fresh[95]), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U36 ( .A(Fresh[94]), .B(
        SubCellInst_SboxInst_15_Q4), .Z(
        SubCellInst_SboxInst_15_AND3_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U35 ( .A(new_AGEMA_signal_1927), .B(
        Fresh[95]), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U34 ( .A(Fresh[93]), .B(
        SubCellInst_SboxInst_15_Q4), .Z(
        SubCellInst_SboxInst_15_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U33 ( .A(Fresh[94]), .B(
        new_AGEMA_signal_1927), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U32 ( .A(new_AGEMA_signal_1926), .B(
        Fresh[93]), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U31 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U30 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U29 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U28 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U27 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U26 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U25 ( .A1(Ciphertext_s2[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U24 ( .A1(Ciphertext_s2[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U23 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n36), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND3_U1_U22 ( .A(Fresh[95]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U21 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U20 ( .A1(SubCellInst_SboxInst_15_n3), .A2(SubCellInst_SboxInst_15_AND3_U1_n35), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND3_U1_U19 ( .A(Fresh[94]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U18 ( .A1(SubCellInst_SboxInst_15_n3), .A2(SubCellInst_SboxInst_15_AND3_U1_n34), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND3_U1_U17 ( .A(Fresh[93]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U16 ( .A1(new_AGEMA_signal_1927), 
        .A2(Ciphertext_s2[62]), .ZN(SubCellInst_SboxInst_15_AND3_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U15 ( .A1(new_AGEMA_signal_1926), 
        .A2(Ciphertext_s1[62]), .ZN(SubCellInst_SboxInst_15_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U14 ( .A1(SubCellInst_SboxInst_15_Q4), .A2(SubCellInst_SboxInst_15_n3), .ZN(SubCellInst_SboxInst_15_AND3_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U13 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND3_U1_n33), .Z(new_AGEMA_signal_2025) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U12 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n32), .B(
        SubCellInst_SboxInst_15_AND3_U1_n31), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U11 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND3_U1_z[2]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U10 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_15_AND3_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U9 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND3_U1_n30), .Z(new_AGEMA_signal_2024) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U8 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n29), .B(
        SubCellInst_SboxInst_15_AND3_U1_n28), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U7 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND3_U1_z[1]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U6 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_15_AND3_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND3_U1_n27), .Z(SubCellInst_SboxInst_15_T2)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n26), .B(
        SubCellInst_SboxInst_15_AND3_U1_n25), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND3_U1_z[0]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_15_AND3_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_a_i_2_s_current_state_reg ( .D(
        Ciphertext_s2[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR7_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3839), 
        .B(SubCellInst_SboxInst_15_T2), .Z(SubCellInst_SboxInst_15_Q7) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3841), 
        .B(new_AGEMA_signal_2024), .Z(new_AGEMA_signal_2150) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR7_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3843), 
        .B(new_AGEMA_signal_2025), .Z(new_AGEMA_signal_2151) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR11_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3845), .B(SubCellInst_SboxInst_15_T0), .Z(SubCellInst_SboxInst_15_L3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3847), .B(new_AGEMA_signal_2022), .Z(new_AGEMA_signal_2152) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR11_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3849), .B(new_AGEMA_signal_2023), .Z(new_AGEMA_signal_2153) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L3), .B(SubCellInst_SboxInst_15_T2), .Z(
        SubCellInst_SboxInst_15_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2152), .B(new_AGEMA_signal_2024), .Z(new_AGEMA_signal_2344) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2153), .B(new_AGEMA_signal_2025), .Z(new_AGEMA_signal_2345) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR13_U1_Ins_0_U1 ( .A(new_AGEMA_signal_3851), .B(SubCellInst_SboxInst_15_T2), .Z(SubCellInst_SboxInst_15_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3853), .B(new_AGEMA_signal_2024), .Z(new_AGEMA_signal_2276) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3855), .B(new_AGEMA_signal_2025), .Z(new_AGEMA_signal_2277) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_2_n1), .B(new_AGEMA_signal_3857), 
        .ZN(AddRoundConstantOutput[62]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2348), .B(1'b0), .Z(new_AGEMA_signal_2436) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2349), .B(1'b0), .Z(new_AGEMA_signal_2437) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[62]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_2_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2276), .Z(new_AGEMA_signal_2348) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2277), .Z(new_AGEMA_signal_2349) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_3_n1), .B(new_AGEMA_signal_3859), 
        .ZN(AddRoundConstantOutput[63]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2438), .B(1'b0), .Z(new_AGEMA_signal_2522) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2439), .B(1'b0), .Z(new_AGEMA_signal_2523) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[63]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_3_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2344), .Z(new_AGEMA_signal_2438) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2345), .Z(new_AGEMA_signal_2439) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_2_n1), .B(1'b0), .ZN(
        AddRoundConstantOutput[46]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2350), .B(1'b0), .Z(new_AGEMA_signal_2440) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2351), .B(1'b0), .Z(new_AGEMA_signal_2441) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_46), .ZN(AddConstXOR_AddConstXOR_XORInst_1_2_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2244), .Z(new_AGEMA_signal_2350) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2245), .Z(new_AGEMA_signal_2351) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_3_n1), .B(1'b0), .ZN(
        AddRoundConstantOutput[47]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2442), .B(1'b0), .Z(new_AGEMA_signal_2526) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2443), .B(1'b0), .Z(new_AGEMA_signal_2527) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_47), .ZN(AddConstXOR_AddConstXOR_XORInst_1_3_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2328), .Z(new_AGEMA_signal_2442) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2329), .Z(new_AGEMA_signal_2443) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_2_n1), .B(new_AGEMA_signal_3861), .ZN(
        ShiftRowsOutput[46]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2352), .B(new_AGEMA_signal_3863), .Z(
        new_AGEMA_signal_2444) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2353), .B(new_AGEMA_signal_3865), .Z(
        new_AGEMA_signal_2445) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[34]), .ZN(AddRoundTweakeyXOR_XORInst_0_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2220), .Z(new_AGEMA_signal_2352) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2221), .Z(new_AGEMA_signal_2353) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_3_n1), .B(new_AGEMA_signal_3867), .ZN(
        ShiftRowsOutput[47]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2446), .B(new_AGEMA_signal_3869), .Z(
        new_AGEMA_signal_2530) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2447), .B(new_AGEMA_signal_3871), .Z(
        new_AGEMA_signal_2531) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[35]), .ZN(AddRoundTweakeyXOR_XORInst_0_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2316), .Z(new_AGEMA_signal_2446) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2317), .Z(new_AGEMA_signal_2447) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_2_n1), .B(new_AGEMA_signal_3873), .ZN(
        ShiftRowsOutput[34]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2354), .B(new_AGEMA_signal_3875), .Z(
        new_AGEMA_signal_2448) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2355), .B(new_AGEMA_signal_3877), .Z(
        new_AGEMA_signal_2449) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[38]), .ZN(AddRoundTweakeyXOR_XORInst_1_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2228), .Z(new_AGEMA_signal_2354) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2229), .Z(new_AGEMA_signal_2355) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_3_n1), .B(new_AGEMA_signal_3879), .ZN(
        ShiftRowsOutput[35]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2450), .B(new_AGEMA_signal_3881), .Z(
        new_AGEMA_signal_2534) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2451), .B(new_AGEMA_signal_3883), .Z(
        new_AGEMA_signal_2535) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[39]), .ZN(AddRoundTweakeyXOR_XORInst_1_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2320), .Z(new_AGEMA_signal_2450) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2321), .Z(new_AGEMA_signal_2451) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_2_n1), .B(new_AGEMA_signal_3885), .ZN(
        ShiftRowsOutput[38]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2356), .B(new_AGEMA_signal_3887), .Z(
        new_AGEMA_signal_2452) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2357), .B(new_AGEMA_signal_3889), .Z(
        new_AGEMA_signal_2453) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[42]), .ZN(AddRoundTweakeyXOR_XORInst_2_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2236), .Z(new_AGEMA_signal_2356) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2237), .Z(new_AGEMA_signal_2357) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_3_n1), .B(new_AGEMA_signal_3891), .ZN(
        ShiftRowsOutput[39]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2454), .B(new_AGEMA_signal_3893), .Z(
        new_AGEMA_signal_2538) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2455), .B(new_AGEMA_signal_3895), .Z(
        new_AGEMA_signal_2539) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[43]), .ZN(AddRoundTweakeyXOR_XORInst_2_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2324), .Z(new_AGEMA_signal_2454) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2325), .Z(new_AGEMA_signal_2455) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_2_n1), .B(new_AGEMA_signal_3897), .ZN(
        ShiftRowsOutput[42]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2540), .B(new_AGEMA_signal_3899), .Z(
        new_AGEMA_signal_2616) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2541), .B(new_AGEMA_signal_3901), .Z(
        new_AGEMA_signal_2617) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[46]), .ZN(AddRoundTweakeyXOR_XORInst_3_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2440), .Z(new_AGEMA_signal_2540) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2441), .Z(new_AGEMA_signal_2541) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_3_n1), .B(new_AGEMA_signal_3903), .ZN(
        ShiftRowsOutput[43]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2618), .B(new_AGEMA_signal_3905), .Z(
        new_AGEMA_signal_2742) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2619), .B(new_AGEMA_signal_3907), .Z(
        new_AGEMA_signal_2743) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[47]), .ZN(AddRoundTweakeyXOR_XORInst_3_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2526), .Z(new_AGEMA_signal_2618) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2527), .Z(new_AGEMA_signal_2619) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_2_n1), .B(new_AGEMA_signal_3909), .ZN(
        MCOutput[34]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2358), .B(new_AGEMA_signal_3911), .Z(
        new_AGEMA_signal_2456) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2359), .B(new_AGEMA_signal_3913), .Z(
        new_AGEMA_signal_2457) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[50]), .ZN(AddRoundTweakeyXOR_XORInst_4_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2252), .Z(new_AGEMA_signal_2358) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2253), .Z(new_AGEMA_signal_2359) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_3_n1), .B(new_AGEMA_signal_3915), .ZN(
        MCOutput[35]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2458), .B(new_AGEMA_signal_3917), .Z(
        new_AGEMA_signal_2544) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2459), .B(new_AGEMA_signal_3919), .Z(
        new_AGEMA_signal_2545) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[51]), .ZN(AddRoundTweakeyXOR_XORInst_4_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2332), .Z(new_AGEMA_signal_2458) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2333), .Z(new_AGEMA_signal_2459) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_2_n1), .B(new_AGEMA_signal_3921), .ZN(
        MCOutput[38]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2360), .B(new_AGEMA_signal_3923), .Z(
        new_AGEMA_signal_2460) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2361), .B(new_AGEMA_signal_3925), .Z(
        new_AGEMA_signal_2461) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[54]), .ZN(AddRoundTweakeyXOR_XORInst_5_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2260), .Z(new_AGEMA_signal_2360) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2261), .Z(new_AGEMA_signal_2361) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_3_n1), .B(new_AGEMA_signal_3927), .ZN(
        MCOutput[39]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2462), .B(new_AGEMA_signal_3929), .Z(
        new_AGEMA_signal_2548) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2463), .B(new_AGEMA_signal_3931), .Z(
        new_AGEMA_signal_2549) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[55]), .ZN(AddRoundTweakeyXOR_XORInst_5_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2336), .Z(new_AGEMA_signal_2462) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2337), .Z(new_AGEMA_signal_2463) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_2_n1), .B(new_AGEMA_signal_3933), .ZN(
        MCOutput[42]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2362), .B(new_AGEMA_signal_3935), .Z(
        new_AGEMA_signal_2464) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2363), .B(new_AGEMA_signal_3937), .Z(
        new_AGEMA_signal_2465) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[58]), .ZN(AddRoundTweakeyXOR_XORInst_6_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2268), .Z(new_AGEMA_signal_2362) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2269), .Z(new_AGEMA_signal_2363) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_3_n1), .B(new_AGEMA_signal_3939), .ZN(
        MCOutput[43]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2466), .B(new_AGEMA_signal_3941), .Z(
        new_AGEMA_signal_2552) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2467), .B(new_AGEMA_signal_3943), .Z(
        new_AGEMA_signal_2553) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[59]), .ZN(AddRoundTweakeyXOR_XORInst_6_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2340), .Z(new_AGEMA_signal_2466) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2341), .Z(new_AGEMA_signal_2467) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_2_n1), .B(new_AGEMA_signal_3945), .ZN(
        MCOutput[46]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2554), .B(new_AGEMA_signal_3947), .Z(
        new_AGEMA_signal_2632) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2555), .B(new_AGEMA_signal_3949), .Z(
        new_AGEMA_signal_2633) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[62]), .ZN(AddRoundTweakeyXOR_XORInst_7_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2436), .Z(new_AGEMA_signal_2554) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2437), .Z(new_AGEMA_signal_2555) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_3_n1), .B(new_AGEMA_signal_3951), .ZN(
        MCOutput[47]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2634), .B(new_AGEMA_signal_3953), .Z(
        new_AGEMA_signal_2752) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2635), .B(new_AGEMA_signal_3955), .Z(
        new_AGEMA_signal_2753) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[63]), .ZN(AddRoundTweakeyXOR_XORInst_7_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2522), .Z(new_AGEMA_signal_2634) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2523), .Z(new_AGEMA_signal_2635) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_2_n2), 
        .B(MCInst_MCR0_XORInst_0_2_n1), .ZN(MCOutput[50]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2558), .B(
        new_AGEMA_signal_2364), .Z(new_AGEMA_signal_2638) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2559), .B(
        new_AGEMA_signal_2365), .Z(new_AGEMA_signal_2639) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[18]), .B(
        ShiftRowsOutput[2]), .ZN(MCInst_MCR0_XORInst_0_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2204), .B(
        new_AGEMA_signal_2180), .Z(new_AGEMA_signal_2364) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2205), .B(
        new_AGEMA_signal_2181), .Z(new_AGEMA_signal_2365) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[34]), 
        .Z(MCInst_MCR0_XORInst_0_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2456), .Z(new_AGEMA_signal_2558) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2457), .Z(new_AGEMA_signal_2559) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_3_n2), 
        .B(MCInst_MCR0_XORInst_0_3_n1), .ZN(MCOutput[51]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2640), .B(
        new_AGEMA_signal_2468), .Z(new_AGEMA_signal_2756) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2641), .B(
        new_AGEMA_signal_2469), .Z(new_AGEMA_signal_2757) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[19]), .B(
        ShiftRowsOutput[3]), .ZN(MCInst_MCR0_XORInst_0_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2308), .B(
        new_AGEMA_signal_2296), .Z(new_AGEMA_signal_2468) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2309), .B(
        new_AGEMA_signal_2297), .Z(new_AGEMA_signal_2469) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[35]), 
        .Z(MCInst_MCR0_XORInst_0_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2544), .Z(new_AGEMA_signal_2640) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2545), .Z(new_AGEMA_signal_2641) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_2_n2), 
        .B(MCInst_MCR0_XORInst_1_2_n1), .ZN(MCOutput[54]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2562), .B(
        new_AGEMA_signal_2366), .Z(new_AGEMA_signal_2642) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2563), .B(
        new_AGEMA_signal_2367), .Z(new_AGEMA_signal_2643) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[22]), .B(
        ShiftRowsOutput[6]), .ZN(MCInst_MCR0_XORInst_1_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2212), .B(
        new_AGEMA_signal_2156), .Z(new_AGEMA_signal_2366) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2213), .B(
        new_AGEMA_signal_2157), .Z(new_AGEMA_signal_2367) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[38]), 
        .Z(MCInst_MCR0_XORInst_1_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2460), .Z(new_AGEMA_signal_2562) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2461), .Z(new_AGEMA_signal_2563) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_3_n2), 
        .B(MCInst_MCR0_XORInst_1_3_n1), .ZN(MCOutput[55]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2644), .B(
        new_AGEMA_signal_2470), .Z(new_AGEMA_signal_2762) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2645), .B(
        new_AGEMA_signal_2471), .Z(new_AGEMA_signal_2763) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[23]), .B(
        ShiftRowsOutput[7]), .ZN(MCInst_MCR0_XORInst_1_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2312), .B(
        new_AGEMA_signal_2284), .Z(new_AGEMA_signal_2470) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2313), .B(
        new_AGEMA_signal_2285), .Z(new_AGEMA_signal_2471) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[39]), 
        .Z(MCInst_MCR0_XORInst_1_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2548), .Z(new_AGEMA_signal_2644) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2549), .Z(new_AGEMA_signal_2645) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_2_n2), 
        .B(MCInst_MCR0_XORInst_2_2_n1), .ZN(MCOutput[58]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2566), .B(
        new_AGEMA_signal_2368), .Z(new_AGEMA_signal_2648) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2567), .B(
        new_AGEMA_signal_2369), .Z(new_AGEMA_signal_2649) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[26]), .B(
        ShiftRowsOutput[10]), .ZN(MCInst_MCR0_XORInst_2_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2188), .B(
        new_AGEMA_signal_2164), .Z(new_AGEMA_signal_2368) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2189), .B(
        new_AGEMA_signal_2165), .Z(new_AGEMA_signal_2369) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[42]), 
        .Z(MCInst_MCR0_XORInst_2_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2464), .Z(new_AGEMA_signal_2566) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2465), .Z(new_AGEMA_signal_2567) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_3_n2), 
        .B(MCInst_MCR0_XORInst_2_3_n1), .ZN(MCOutput[59]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2650), .B(
        new_AGEMA_signal_2472), .Z(new_AGEMA_signal_2766) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2651), .B(
        new_AGEMA_signal_2473), .Z(new_AGEMA_signal_2767) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[27]), .B(
        ShiftRowsOutput[11]), .ZN(MCInst_MCR0_XORInst_2_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2300), .B(
        new_AGEMA_signal_2288), .Z(new_AGEMA_signal_2472) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2301), .B(
        new_AGEMA_signal_2289), .Z(new_AGEMA_signal_2473) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[43]), 
        .Z(MCInst_MCR0_XORInst_2_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2552), .Z(new_AGEMA_signal_2650) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2553), .Z(new_AGEMA_signal_2651) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_2_n2), 
        .B(MCInst_MCR0_XORInst_3_2_n1), .ZN(MCOutput[62]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2768), .B(
        new_AGEMA_signal_2370), .Z(new_AGEMA_signal_2870) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2769), .B(
        new_AGEMA_signal_2371), .Z(new_AGEMA_signal_2871) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[30]), .B(
        ShiftRowsOutput[14]), .ZN(MCInst_MCR0_XORInst_3_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2196), .B(
        new_AGEMA_signal_2172), .Z(new_AGEMA_signal_2370) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2197), .B(
        new_AGEMA_signal_2173), .Z(new_AGEMA_signal_2371) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[46]), 
        .Z(MCInst_MCR0_XORInst_3_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2632), .Z(new_AGEMA_signal_2768) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2633), .Z(new_AGEMA_signal_2769) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_3_n2), 
        .B(MCInst_MCR0_XORInst_3_3_n1), .ZN(MCOutput[63]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2872), .B(
        new_AGEMA_signal_2474), .Z(new_AGEMA_signal_2970) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2873), .B(
        new_AGEMA_signal_2475), .Z(new_AGEMA_signal_2971) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[31]), .B(
        ShiftRowsOutput[15]), .ZN(MCInst_MCR0_XORInst_3_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2304), .B(
        new_AGEMA_signal_2292), .Z(new_AGEMA_signal_2474) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2305), .B(
        new_AGEMA_signal_2293), .Z(new_AGEMA_signal_2475) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[47]), 
        .Z(MCInst_MCR0_XORInst_3_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2752), .Z(new_AGEMA_signal_2872) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2753), .Z(new_AGEMA_signal_2873) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_2_n1), 
        .B(ShiftRowsOutput[18]), .ZN(MCOutput[18]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2570), .B(
        new_AGEMA_signal_2204), .Z(new_AGEMA_signal_2654) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2571), .B(
        new_AGEMA_signal_2205), .Z(new_AGEMA_signal_2655) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[34]), .ZN(MCInst_MCR2_XORInst_0_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2448), .Z(new_AGEMA_signal_2570) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2449), .Z(new_AGEMA_signal_2571) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_3_n1), 
        .B(ShiftRowsOutput[19]), .ZN(MCOutput[19]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2656), .B(
        new_AGEMA_signal_2308), .Z(new_AGEMA_signal_2772) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2657), .B(
        new_AGEMA_signal_2309), .Z(new_AGEMA_signal_2773) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[35]), .ZN(MCInst_MCR2_XORInst_0_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2534), .Z(new_AGEMA_signal_2656) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2535), .Z(new_AGEMA_signal_2657) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_2_n1), 
        .B(ShiftRowsOutput[22]), .ZN(MCOutput[22]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2572), .B(
        new_AGEMA_signal_2212), .Z(new_AGEMA_signal_2658) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2573), .B(
        new_AGEMA_signal_2213), .Z(new_AGEMA_signal_2659) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[38]), .ZN(MCInst_MCR2_XORInst_1_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2452), .Z(new_AGEMA_signal_2572) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2453), .Z(new_AGEMA_signal_2573) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_3_n1), 
        .B(ShiftRowsOutput[23]), .ZN(MCOutput[23]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2660), .B(
        new_AGEMA_signal_2312), .Z(new_AGEMA_signal_2776) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2661), .B(
        new_AGEMA_signal_2313), .Z(new_AGEMA_signal_2777) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[39]), .ZN(MCInst_MCR2_XORInst_1_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2538), .Z(new_AGEMA_signal_2660) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2539), .Z(new_AGEMA_signal_2661) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_2_n1), 
        .B(ShiftRowsOutput[26]), .ZN(MCOutput[26]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2778), .B(
        new_AGEMA_signal_2188), .Z(new_AGEMA_signal_2882) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2779), .B(
        new_AGEMA_signal_2189), .Z(new_AGEMA_signal_2883) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[42]), .ZN(MCInst_MCR2_XORInst_2_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2616), .Z(new_AGEMA_signal_2778) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2617), .Z(new_AGEMA_signal_2779) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_3_n1), 
        .B(ShiftRowsOutput[27]), .ZN(MCOutput[27]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2884), .B(
        new_AGEMA_signal_2300), .Z(new_AGEMA_signal_2978) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2885), .B(
        new_AGEMA_signal_2301), .Z(new_AGEMA_signal_2979) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[43]), .ZN(MCInst_MCR2_XORInst_2_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2742), .Z(new_AGEMA_signal_2884) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2743), .Z(new_AGEMA_signal_2885) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_2_n1), 
        .B(ShiftRowsOutput[30]), .ZN(MCOutput[30]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2574), .B(
        new_AGEMA_signal_2196), .Z(new_AGEMA_signal_2662) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2575), .B(
        new_AGEMA_signal_2197), .Z(new_AGEMA_signal_2663) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[46]), .ZN(MCInst_MCR2_XORInst_3_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2444), .Z(new_AGEMA_signal_2574) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2445), .Z(new_AGEMA_signal_2575) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_3_n1), 
        .B(ShiftRowsOutput[31]), .ZN(MCOutput[31]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2664), .B(
        new_AGEMA_signal_2304), .Z(new_AGEMA_signal_2782) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2665), .B(
        new_AGEMA_signal_2305), .Z(new_AGEMA_signal_2783) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[47]), .ZN(MCInst_MCR2_XORInst_3_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2530), .Z(new_AGEMA_signal_2664) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2531), .Z(new_AGEMA_signal_2665) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_2_n1), 
        .B(ShiftRowsOutput[18]), .ZN(MCOutput[2]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2576), .B(
        new_AGEMA_signal_2204), .Z(new_AGEMA_signal_2666) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2577), .B(
        new_AGEMA_signal_2205), .Z(new_AGEMA_signal_2667) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[34]), 
        .ZN(MCInst_MCR3_XORInst_0_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2456), .Z(new_AGEMA_signal_2576) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2457), .Z(new_AGEMA_signal_2577) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_3_n1), 
        .B(ShiftRowsOutput[19]), .ZN(MCOutput[3]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2668), .B(
        new_AGEMA_signal_2308), .Z(new_AGEMA_signal_2786) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2669), .B(
        new_AGEMA_signal_2309), .Z(new_AGEMA_signal_2787) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[35]), 
        .ZN(MCInst_MCR3_XORInst_0_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2544), .Z(new_AGEMA_signal_2668) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2545), .Z(new_AGEMA_signal_2669) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_2_n1), 
        .B(ShiftRowsOutput[22]), .ZN(MCOutput[6]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2578), .B(
        new_AGEMA_signal_2212), .Z(new_AGEMA_signal_2670) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2579), .B(
        new_AGEMA_signal_2213), .Z(new_AGEMA_signal_2671) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[38]), 
        .ZN(MCInst_MCR3_XORInst_1_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2460), .Z(new_AGEMA_signal_2578) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2461), .Z(new_AGEMA_signal_2579) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_3_n1), 
        .B(ShiftRowsOutput[23]), .ZN(MCOutput[7]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2672), .B(
        new_AGEMA_signal_2312), .Z(new_AGEMA_signal_2790) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2673), .B(
        new_AGEMA_signal_2313), .Z(new_AGEMA_signal_2791) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[39]), 
        .ZN(MCInst_MCR3_XORInst_1_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2548), .Z(new_AGEMA_signal_2672) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2549), .Z(new_AGEMA_signal_2673) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_2_n1), 
        .B(ShiftRowsOutput[26]), .ZN(MCOutput[10]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2580), .B(
        new_AGEMA_signal_2188), .Z(new_AGEMA_signal_2674) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2581), .B(
        new_AGEMA_signal_2189), .Z(new_AGEMA_signal_2675) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[42]), 
        .ZN(MCInst_MCR3_XORInst_2_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2464), .Z(new_AGEMA_signal_2580) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2465), .Z(new_AGEMA_signal_2581) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_3_n1), 
        .B(ShiftRowsOutput[27]), .ZN(MCOutput[11]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2676), .B(
        new_AGEMA_signal_2300), .Z(new_AGEMA_signal_2794) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2677), .B(
        new_AGEMA_signal_2301), .Z(new_AGEMA_signal_2795) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[43]), 
        .ZN(MCInst_MCR3_XORInst_2_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2552), .Z(new_AGEMA_signal_2676) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2553), .Z(new_AGEMA_signal_2677) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_2_n1), 
        .B(ShiftRowsOutput[30]), .ZN(MCOutput[14]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2796), .B(
        new_AGEMA_signal_2196), .Z(new_AGEMA_signal_2902) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2797), .B(
        new_AGEMA_signal_2197), .Z(new_AGEMA_signal_2903) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[46]), 
        .ZN(MCInst_MCR3_XORInst_3_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2632), .Z(new_AGEMA_signal_2796) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2633), .Z(new_AGEMA_signal_2797) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_3_n1), 
        .B(ShiftRowsOutput[31]), .ZN(MCOutput[15]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2904), .B(
        new_AGEMA_signal_2304), .Z(new_AGEMA_signal_2990) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2905), .B(
        new_AGEMA_signal_2305), .Z(new_AGEMA_signal_2991) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[47]), 
        .ZN(MCInst_MCR3_XORInst_3_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2752), .Z(new_AGEMA_signal_2904) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2753), .Z(new_AGEMA_signal_2905) );
  DFF_X1 new_AGEMA_reg_buffer_1001_s_current_state_reg ( .D(
        new_AGEMA_signal_3278), .CK(clk), .Q(new_AGEMA_signal_3279), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1003_s_current_state_reg ( .D(
        new_AGEMA_signal_3280), .CK(clk), .Q(new_AGEMA_signal_3281), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1005_s_current_state_reg ( .D(
        new_AGEMA_signal_3282), .CK(clk), .Q(new_AGEMA_signal_3283), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1007_s_current_state_reg ( .D(
        new_AGEMA_signal_3284), .CK(clk), .Q(new_AGEMA_signal_3285), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1009_s_current_state_reg ( .D(
        new_AGEMA_signal_3286), .CK(clk), .Q(new_AGEMA_signal_3287), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1011_s_current_state_reg ( .D(
        new_AGEMA_signal_3288), .CK(clk), .Q(new_AGEMA_signal_3289), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1013_s_current_state_reg ( .D(
        new_AGEMA_signal_3290), .CK(clk), .Q(new_AGEMA_signal_3291), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1015_s_current_state_reg ( .D(
        new_AGEMA_signal_3292), .CK(clk), .Q(new_AGEMA_signal_3293), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1017_s_current_state_reg ( .D(
        new_AGEMA_signal_3294), .CK(clk), .Q(new_AGEMA_signal_3295), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1019_s_current_state_reg ( .D(
        new_AGEMA_signal_3296), .CK(clk), .Q(new_AGEMA_signal_3297), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1021_s_current_state_reg ( .D(
        new_AGEMA_signal_3298), .CK(clk), .Q(new_AGEMA_signal_3299), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1023_s_current_state_reg ( .D(
        new_AGEMA_signal_3300), .CK(clk), .Q(new_AGEMA_signal_3301), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1025_s_current_state_reg ( .D(
        new_AGEMA_signal_3302), .CK(clk), .Q(new_AGEMA_signal_3303), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1027_s_current_state_reg ( .D(
        new_AGEMA_signal_3304), .CK(clk), .Q(new_AGEMA_signal_3305), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1029_s_current_state_reg ( .D(
        new_AGEMA_signal_3306), .CK(clk), .Q(new_AGEMA_signal_3307), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1031_s_current_state_reg ( .D(
        new_AGEMA_signal_3308), .CK(clk), .Q(new_AGEMA_signal_3309), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1033_s_current_state_reg ( .D(
        new_AGEMA_signal_3310), .CK(clk), .Q(new_AGEMA_signal_3311), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1035_s_current_state_reg ( .D(
        new_AGEMA_signal_3312), .CK(clk), .Q(new_AGEMA_signal_3313), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1037_s_current_state_reg ( .D(
        new_AGEMA_signal_3314), .CK(clk), .Q(new_AGEMA_signal_3315), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1039_s_current_state_reg ( .D(
        new_AGEMA_signal_3316), .CK(clk), .Q(new_AGEMA_signal_3317), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1041_s_current_state_reg ( .D(
        new_AGEMA_signal_3318), .CK(clk), .Q(new_AGEMA_signal_3319), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1043_s_current_state_reg ( .D(
        new_AGEMA_signal_3320), .CK(clk), .Q(new_AGEMA_signal_3321), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1045_s_current_state_reg ( .D(
        new_AGEMA_signal_3322), .CK(clk), .Q(new_AGEMA_signal_3323), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1047_s_current_state_reg ( .D(
        new_AGEMA_signal_3324), .CK(clk), .Q(new_AGEMA_signal_3325), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1049_s_current_state_reg ( .D(
        new_AGEMA_signal_3326), .CK(clk), .Q(new_AGEMA_signal_3327), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1051_s_current_state_reg ( .D(
        new_AGEMA_signal_3328), .CK(clk), .Q(new_AGEMA_signal_3329), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1053_s_current_state_reg ( .D(
        new_AGEMA_signal_3330), .CK(clk), .Q(new_AGEMA_signal_3331), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1055_s_current_state_reg ( .D(
        new_AGEMA_signal_3332), .CK(clk), .Q(new_AGEMA_signal_3333), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1057_s_current_state_reg ( .D(
        new_AGEMA_signal_3334), .CK(clk), .Q(new_AGEMA_signal_3335), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1059_s_current_state_reg ( .D(
        new_AGEMA_signal_3336), .CK(clk), .Q(new_AGEMA_signal_3337), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1061_s_current_state_reg ( .D(
        new_AGEMA_signal_3338), .CK(clk), .Q(new_AGEMA_signal_3339), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1063_s_current_state_reg ( .D(
        new_AGEMA_signal_3340), .CK(clk), .Q(new_AGEMA_signal_3341), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1065_s_current_state_reg ( .D(
        new_AGEMA_signal_3342), .CK(clk), .Q(new_AGEMA_signal_3343), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1067_s_current_state_reg ( .D(
        new_AGEMA_signal_3344), .CK(clk), .Q(new_AGEMA_signal_3345), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1069_s_current_state_reg ( .D(
        new_AGEMA_signal_3346), .CK(clk), .Q(new_AGEMA_signal_3347), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1071_s_current_state_reg ( .D(
        new_AGEMA_signal_3348), .CK(clk), .Q(new_AGEMA_signal_3349), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1073_s_current_state_reg ( .D(
        new_AGEMA_signal_3350), .CK(clk), .Q(new_AGEMA_signal_3351), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1075_s_current_state_reg ( .D(
        new_AGEMA_signal_3352), .CK(clk), .Q(new_AGEMA_signal_3353), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1077_s_current_state_reg ( .D(
        new_AGEMA_signal_3354), .CK(clk), .Q(new_AGEMA_signal_3355), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1079_s_current_state_reg ( .D(
        new_AGEMA_signal_3356), .CK(clk), .Q(new_AGEMA_signal_3357), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1081_s_current_state_reg ( .D(
        new_AGEMA_signal_3358), .CK(clk), .Q(new_AGEMA_signal_3359), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1083_s_current_state_reg ( .D(
        new_AGEMA_signal_3360), .CK(clk), .Q(new_AGEMA_signal_3361), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1085_s_current_state_reg ( .D(
        new_AGEMA_signal_3362), .CK(clk), .Q(new_AGEMA_signal_3363), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1087_s_current_state_reg ( .D(
        new_AGEMA_signal_3364), .CK(clk), .Q(new_AGEMA_signal_3365), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1089_s_current_state_reg ( .D(
        new_AGEMA_signal_3366), .CK(clk), .Q(new_AGEMA_signal_3367), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1091_s_current_state_reg ( .D(
        new_AGEMA_signal_3368), .CK(clk), .Q(new_AGEMA_signal_3369), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1093_s_current_state_reg ( .D(
        new_AGEMA_signal_3370), .CK(clk), .Q(new_AGEMA_signal_3371), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1095_s_current_state_reg ( .D(
        new_AGEMA_signal_3372), .CK(clk), .Q(new_AGEMA_signal_3373), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1097_s_current_state_reg ( .D(
        new_AGEMA_signal_3374), .CK(clk), .Q(new_AGEMA_signal_3375), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1099_s_current_state_reg ( .D(
        new_AGEMA_signal_3376), .CK(clk), .Q(new_AGEMA_signal_3377), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1101_s_current_state_reg ( .D(
        new_AGEMA_signal_3378), .CK(clk), .Q(new_AGEMA_signal_3379), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1103_s_current_state_reg ( .D(
        new_AGEMA_signal_3380), .CK(clk), .Q(new_AGEMA_signal_3381), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1105_s_current_state_reg ( .D(
        new_AGEMA_signal_3382), .CK(clk), .Q(new_AGEMA_signal_3383), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1107_s_current_state_reg ( .D(
        new_AGEMA_signal_3384), .CK(clk), .Q(new_AGEMA_signal_3385), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1109_s_current_state_reg ( .D(
        new_AGEMA_signal_3386), .CK(clk), .Q(new_AGEMA_signal_3387), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1111_s_current_state_reg ( .D(
        new_AGEMA_signal_3388), .CK(clk), .Q(new_AGEMA_signal_3389), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1113_s_current_state_reg ( .D(
        new_AGEMA_signal_3390), .CK(clk), .Q(new_AGEMA_signal_3391), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1115_s_current_state_reg ( .D(
        new_AGEMA_signal_3392), .CK(clk), .Q(new_AGEMA_signal_3393), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1117_s_current_state_reg ( .D(
        new_AGEMA_signal_3394), .CK(clk), .Q(new_AGEMA_signal_3395), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1119_s_current_state_reg ( .D(
        new_AGEMA_signal_3396), .CK(clk), .Q(new_AGEMA_signal_3397), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1121_s_current_state_reg ( .D(
        new_AGEMA_signal_3398), .CK(clk), .Q(new_AGEMA_signal_3399), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1123_s_current_state_reg ( .D(
        new_AGEMA_signal_3400), .CK(clk), .Q(new_AGEMA_signal_3401), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1125_s_current_state_reg ( .D(
        new_AGEMA_signal_3402), .CK(clk), .Q(new_AGEMA_signal_3403), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1127_s_current_state_reg ( .D(
        new_AGEMA_signal_3404), .CK(clk), .Q(new_AGEMA_signal_3405), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1129_s_current_state_reg ( .D(
        new_AGEMA_signal_3406), .CK(clk), .Q(new_AGEMA_signal_3407), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1131_s_current_state_reg ( .D(
        new_AGEMA_signal_3408), .CK(clk), .Q(new_AGEMA_signal_3409), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1133_s_current_state_reg ( .D(
        new_AGEMA_signal_3410), .CK(clk), .Q(new_AGEMA_signal_3411), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1135_s_current_state_reg ( .D(
        new_AGEMA_signal_3412), .CK(clk), .Q(new_AGEMA_signal_3413), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1137_s_current_state_reg ( .D(
        new_AGEMA_signal_3414), .CK(clk), .Q(new_AGEMA_signal_3415), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1139_s_current_state_reg ( .D(
        new_AGEMA_signal_3416), .CK(clk), .Q(new_AGEMA_signal_3417), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1141_s_current_state_reg ( .D(
        new_AGEMA_signal_3418), .CK(clk), .Q(new_AGEMA_signal_3419), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1143_s_current_state_reg ( .D(
        new_AGEMA_signal_3420), .CK(clk), .Q(new_AGEMA_signal_3421), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1145_s_current_state_reg ( .D(
        new_AGEMA_signal_3422), .CK(clk), .Q(new_AGEMA_signal_3423), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1147_s_current_state_reg ( .D(
        new_AGEMA_signal_3424), .CK(clk), .Q(new_AGEMA_signal_3425), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1149_s_current_state_reg ( .D(
        new_AGEMA_signal_3426), .CK(clk), .Q(new_AGEMA_signal_3427), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1151_s_current_state_reg ( .D(
        new_AGEMA_signal_3428), .CK(clk), .Q(new_AGEMA_signal_3429), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1153_s_current_state_reg ( .D(
        new_AGEMA_signal_3430), .CK(clk), .Q(new_AGEMA_signal_3431), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1155_s_current_state_reg ( .D(
        new_AGEMA_signal_3432), .CK(clk), .Q(new_AGEMA_signal_3433), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1157_s_current_state_reg ( .D(
        new_AGEMA_signal_3434), .CK(clk), .Q(new_AGEMA_signal_3435), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1159_s_current_state_reg ( .D(
        new_AGEMA_signal_3436), .CK(clk), .Q(new_AGEMA_signal_3437), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1161_s_current_state_reg ( .D(
        new_AGEMA_signal_3438), .CK(clk), .Q(new_AGEMA_signal_3439), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1163_s_current_state_reg ( .D(
        new_AGEMA_signal_3440), .CK(clk), .Q(new_AGEMA_signal_3441), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1165_s_current_state_reg ( .D(
        new_AGEMA_signal_3442), .CK(clk), .Q(new_AGEMA_signal_3443), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1167_s_current_state_reg ( .D(
        new_AGEMA_signal_3444), .CK(clk), .Q(new_AGEMA_signal_3445), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1169_s_current_state_reg ( .D(
        new_AGEMA_signal_3446), .CK(clk), .Q(new_AGEMA_signal_3447), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1171_s_current_state_reg ( .D(
        new_AGEMA_signal_3448), .CK(clk), .Q(new_AGEMA_signal_3449), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1173_s_current_state_reg ( .D(
        new_AGEMA_signal_3450), .CK(clk), .Q(new_AGEMA_signal_3451), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1175_s_current_state_reg ( .D(
        new_AGEMA_signal_3452), .CK(clk), .Q(new_AGEMA_signal_3453), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1177_s_current_state_reg ( .D(
        new_AGEMA_signal_3454), .CK(clk), .Q(new_AGEMA_signal_3455), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1179_s_current_state_reg ( .D(
        new_AGEMA_signal_3456), .CK(clk), .Q(new_AGEMA_signal_3457), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1181_s_current_state_reg ( .D(
        new_AGEMA_signal_3458), .CK(clk), .Q(new_AGEMA_signal_3459), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1183_s_current_state_reg ( .D(
        new_AGEMA_signal_3460), .CK(clk), .Q(new_AGEMA_signal_3461), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1185_s_current_state_reg ( .D(
        new_AGEMA_signal_3462), .CK(clk), .Q(new_AGEMA_signal_3463), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1187_s_current_state_reg ( .D(
        new_AGEMA_signal_3464), .CK(clk), .Q(new_AGEMA_signal_3465), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1189_s_current_state_reg ( .D(
        new_AGEMA_signal_3466), .CK(clk), .Q(new_AGEMA_signal_3467), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1191_s_current_state_reg ( .D(
        new_AGEMA_signal_3468), .CK(clk), .Q(new_AGEMA_signal_3469), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1193_s_current_state_reg ( .D(
        new_AGEMA_signal_3470), .CK(clk), .Q(new_AGEMA_signal_3471), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1195_s_current_state_reg ( .D(
        new_AGEMA_signal_3472), .CK(clk), .Q(new_AGEMA_signal_3473), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1197_s_current_state_reg ( .D(
        new_AGEMA_signal_3474), .CK(clk), .Q(new_AGEMA_signal_3475), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1199_s_current_state_reg ( .D(
        new_AGEMA_signal_3476), .CK(clk), .Q(new_AGEMA_signal_3477), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1201_s_current_state_reg ( .D(
        new_AGEMA_signal_3478), .CK(clk), .Q(new_AGEMA_signal_3479), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1203_s_current_state_reg ( .D(
        new_AGEMA_signal_3480), .CK(clk), .Q(new_AGEMA_signal_3481), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1205_s_current_state_reg ( .D(
        new_AGEMA_signal_3482), .CK(clk), .Q(new_AGEMA_signal_3483), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1207_s_current_state_reg ( .D(
        new_AGEMA_signal_3484), .CK(clk), .Q(new_AGEMA_signal_3485), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1209_s_current_state_reg ( .D(
        new_AGEMA_signal_3486), .CK(clk), .Q(new_AGEMA_signal_3487), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1211_s_current_state_reg ( .D(
        new_AGEMA_signal_3488), .CK(clk), .Q(new_AGEMA_signal_3489), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1213_s_current_state_reg ( .D(
        new_AGEMA_signal_3490), .CK(clk), .Q(new_AGEMA_signal_3491), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1215_s_current_state_reg ( .D(
        new_AGEMA_signal_3492), .CK(clk), .Q(new_AGEMA_signal_3493), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1217_s_current_state_reg ( .D(
        new_AGEMA_signal_3494), .CK(clk), .Q(new_AGEMA_signal_3495), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1219_s_current_state_reg ( .D(
        new_AGEMA_signal_3496), .CK(clk), .Q(new_AGEMA_signal_3497), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1221_s_current_state_reg ( .D(
        new_AGEMA_signal_3498), .CK(clk), .Q(new_AGEMA_signal_3499), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1223_s_current_state_reg ( .D(
        new_AGEMA_signal_3500), .CK(clk), .Q(new_AGEMA_signal_3501), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1225_s_current_state_reg ( .D(
        new_AGEMA_signal_3502), .CK(clk), .Q(new_AGEMA_signal_3503), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1227_s_current_state_reg ( .D(
        new_AGEMA_signal_3504), .CK(clk), .Q(new_AGEMA_signal_3505), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1229_s_current_state_reg ( .D(
        new_AGEMA_signal_3506), .CK(clk), .Q(new_AGEMA_signal_3507), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1231_s_current_state_reg ( .D(
        new_AGEMA_signal_3508), .CK(clk), .Q(new_AGEMA_signal_3509), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1233_s_current_state_reg ( .D(
        new_AGEMA_signal_3510), .CK(clk), .Q(new_AGEMA_signal_3511), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1235_s_current_state_reg ( .D(
        new_AGEMA_signal_3512), .CK(clk), .Q(new_AGEMA_signal_3513), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1237_s_current_state_reg ( .D(
        new_AGEMA_signal_3514), .CK(clk), .Q(new_AGEMA_signal_3515), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1239_s_current_state_reg ( .D(
        new_AGEMA_signal_3516), .CK(clk), .Q(new_AGEMA_signal_3517), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1241_s_current_state_reg ( .D(
        new_AGEMA_signal_3518), .CK(clk), .Q(new_AGEMA_signal_3519), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1243_s_current_state_reg ( .D(
        new_AGEMA_signal_3520), .CK(clk), .Q(new_AGEMA_signal_3521), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1245_s_current_state_reg ( .D(
        new_AGEMA_signal_3522), .CK(clk), .Q(new_AGEMA_signal_3523), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1247_s_current_state_reg ( .D(
        new_AGEMA_signal_3524), .CK(clk), .Q(new_AGEMA_signal_3525), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1249_s_current_state_reg ( .D(
        new_AGEMA_signal_3526), .CK(clk), .Q(new_AGEMA_signal_3527), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1251_s_current_state_reg ( .D(
        new_AGEMA_signal_3528), .CK(clk), .Q(new_AGEMA_signal_3529), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1253_s_current_state_reg ( .D(
        new_AGEMA_signal_3530), .CK(clk), .Q(new_AGEMA_signal_3531), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1255_s_current_state_reg ( .D(
        new_AGEMA_signal_3532), .CK(clk), .Q(new_AGEMA_signal_3533), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1257_s_current_state_reg ( .D(
        new_AGEMA_signal_3534), .CK(clk), .Q(new_AGEMA_signal_3535), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1259_s_current_state_reg ( .D(
        new_AGEMA_signal_3536), .CK(clk), .Q(new_AGEMA_signal_3537), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1261_s_current_state_reg ( .D(
        new_AGEMA_signal_3538), .CK(clk), .Q(new_AGEMA_signal_3539), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1263_s_current_state_reg ( .D(
        new_AGEMA_signal_3540), .CK(clk), .Q(new_AGEMA_signal_3541), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1265_s_current_state_reg ( .D(
        new_AGEMA_signal_3542), .CK(clk), .Q(new_AGEMA_signal_3543), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1267_s_current_state_reg ( .D(
        new_AGEMA_signal_3544), .CK(clk), .Q(new_AGEMA_signal_3545), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1269_s_current_state_reg ( .D(
        new_AGEMA_signal_3546), .CK(clk), .Q(new_AGEMA_signal_3547), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1271_s_current_state_reg ( .D(
        new_AGEMA_signal_3548), .CK(clk), .Q(new_AGEMA_signal_3549), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1273_s_current_state_reg ( .D(
        new_AGEMA_signal_3550), .CK(clk), .Q(new_AGEMA_signal_3551), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1275_s_current_state_reg ( .D(
        new_AGEMA_signal_3552), .CK(clk), .Q(new_AGEMA_signal_3553), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1277_s_current_state_reg ( .D(
        new_AGEMA_signal_3554), .CK(clk), .Q(new_AGEMA_signal_3555), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1279_s_current_state_reg ( .D(
        new_AGEMA_signal_3556), .CK(clk), .Q(new_AGEMA_signal_3557), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1281_s_current_state_reg ( .D(
        new_AGEMA_signal_3558), .CK(clk), .Q(new_AGEMA_signal_3559), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1283_s_current_state_reg ( .D(
        new_AGEMA_signal_3560), .CK(clk), .Q(new_AGEMA_signal_3561), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1285_s_current_state_reg ( .D(
        new_AGEMA_signal_3562), .CK(clk), .Q(new_AGEMA_signal_3563), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1287_s_current_state_reg ( .D(
        new_AGEMA_signal_3564), .CK(clk), .Q(new_AGEMA_signal_3565), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1289_s_current_state_reg ( .D(
        new_AGEMA_signal_3566), .CK(clk), .Q(new_AGEMA_signal_3567), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1291_s_current_state_reg ( .D(
        new_AGEMA_signal_3568), .CK(clk), .Q(new_AGEMA_signal_3569), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1293_s_current_state_reg ( .D(
        new_AGEMA_signal_3570), .CK(clk), .Q(new_AGEMA_signal_3571), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1295_s_current_state_reg ( .D(
        new_AGEMA_signal_3572), .CK(clk), .Q(new_AGEMA_signal_3573), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1297_s_current_state_reg ( .D(
        new_AGEMA_signal_3574), .CK(clk), .Q(new_AGEMA_signal_3575), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1299_s_current_state_reg ( .D(
        new_AGEMA_signal_3576), .CK(clk), .Q(new_AGEMA_signal_3577), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1301_s_current_state_reg ( .D(
        new_AGEMA_signal_3578), .CK(clk), .Q(new_AGEMA_signal_3579), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1303_s_current_state_reg ( .D(
        new_AGEMA_signal_3580), .CK(clk), .Q(new_AGEMA_signal_3581), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1305_s_current_state_reg ( .D(
        new_AGEMA_signal_3582), .CK(clk), .Q(new_AGEMA_signal_3583), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1307_s_current_state_reg ( .D(
        new_AGEMA_signal_3584), .CK(clk), .Q(new_AGEMA_signal_3585), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1309_s_current_state_reg ( .D(
        new_AGEMA_signal_3586), .CK(clk), .Q(new_AGEMA_signal_3587), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1311_s_current_state_reg ( .D(
        new_AGEMA_signal_3588), .CK(clk), .Q(new_AGEMA_signal_3589), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1313_s_current_state_reg ( .D(
        new_AGEMA_signal_3590), .CK(clk), .Q(new_AGEMA_signal_3591), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1315_s_current_state_reg ( .D(
        new_AGEMA_signal_3592), .CK(clk), .Q(new_AGEMA_signal_3593), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1317_s_current_state_reg ( .D(
        new_AGEMA_signal_3594), .CK(clk), .Q(new_AGEMA_signal_3595), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1319_s_current_state_reg ( .D(
        new_AGEMA_signal_3596), .CK(clk), .Q(new_AGEMA_signal_3597), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1321_s_current_state_reg ( .D(
        new_AGEMA_signal_3598), .CK(clk), .Q(new_AGEMA_signal_3599), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1323_s_current_state_reg ( .D(
        new_AGEMA_signal_3600), .CK(clk), .Q(new_AGEMA_signal_3601), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1325_s_current_state_reg ( .D(
        new_AGEMA_signal_3602), .CK(clk), .Q(new_AGEMA_signal_3603), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1327_s_current_state_reg ( .D(
        new_AGEMA_signal_3604), .CK(clk), .Q(new_AGEMA_signal_3605), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1329_s_current_state_reg ( .D(
        new_AGEMA_signal_3606), .CK(clk), .Q(new_AGEMA_signal_3607), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1331_s_current_state_reg ( .D(
        new_AGEMA_signal_3608), .CK(clk), .Q(new_AGEMA_signal_3609), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1333_s_current_state_reg ( .D(
        new_AGEMA_signal_3610), .CK(clk), .Q(new_AGEMA_signal_3611), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1335_s_current_state_reg ( .D(
        new_AGEMA_signal_3612), .CK(clk), .Q(new_AGEMA_signal_3613), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1337_s_current_state_reg ( .D(
        new_AGEMA_signal_3614), .CK(clk), .Q(new_AGEMA_signal_3615), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1339_s_current_state_reg ( .D(
        new_AGEMA_signal_3616), .CK(clk), .Q(new_AGEMA_signal_3617), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1341_s_current_state_reg ( .D(
        new_AGEMA_signal_3618), .CK(clk), .Q(new_AGEMA_signal_3619), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1343_s_current_state_reg ( .D(
        new_AGEMA_signal_3620), .CK(clk), .Q(new_AGEMA_signal_3621), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1345_s_current_state_reg ( .D(
        new_AGEMA_signal_3622), .CK(clk), .Q(new_AGEMA_signal_3623), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1347_s_current_state_reg ( .D(
        new_AGEMA_signal_3624), .CK(clk), .Q(new_AGEMA_signal_3625), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1349_s_current_state_reg ( .D(
        new_AGEMA_signal_3626), .CK(clk), .Q(new_AGEMA_signal_3627), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1351_s_current_state_reg ( .D(
        new_AGEMA_signal_3628), .CK(clk), .Q(new_AGEMA_signal_3629), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1353_s_current_state_reg ( .D(
        new_AGEMA_signal_3630), .CK(clk), .Q(new_AGEMA_signal_3631), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1355_s_current_state_reg ( .D(
        new_AGEMA_signal_3632), .CK(clk), .Q(new_AGEMA_signal_3633), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1357_s_current_state_reg ( .D(
        new_AGEMA_signal_3634), .CK(clk), .Q(new_AGEMA_signal_3635), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1359_s_current_state_reg ( .D(
        new_AGEMA_signal_3636), .CK(clk), .Q(new_AGEMA_signal_3637), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1361_s_current_state_reg ( .D(
        new_AGEMA_signal_3638), .CK(clk), .Q(new_AGEMA_signal_3639), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1363_s_current_state_reg ( .D(
        new_AGEMA_signal_3640), .CK(clk), .Q(new_AGEMA_signal_3641), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1365_s_current_state_reg ( .D(
        new_AGEMA_signal_3642), .CK(clk), .Q(new_AGEMA_signal_3643), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1367_s_current_state_reg ( .D(
        new_AGEMA_signal_3644), .CK(clk), .Q(new_AGEMA_signal_3645), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1369_s_current_state_reg ( .D(
        new_AGEMA_signal_3646), .CK(clk), .Q(new_AGEMA_signal_3647), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1371_s_current_state_reg ( .D(
        new_AGEMA_signal_3648), .CK(clk), .Q(new_AGEMA_signal_3649), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1373_s_current_state_reg ( .D(
        new_AGEMA_signal_3650), .CK(clk), .Q(new_AGEMA_signal_3651), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1375_s_current_state_reg ( .D(
        new_AGEMA_signal_3652), .CK(clk), .Q(new_AGEMA_signal_3653), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1377_s_current_state_reg ( .D(
        new_AGEMA_signal_3654), .CK(clk), .Q(new_AGEMA_signal_3655), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1379_s_current_state_reg ( .D(
        new_AGEMA_signal_3656), .CK(clk), .Q(new_AGEMA_signal_3657), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1381_s_current_state_reg ( .D(
        new_AGEMA_signal_3658), .CK(clk), .Q(new_AGEMA_signal_3659), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1383_s_current_state_reg ( .D(
        new_AGEMA_signal_3660), .CK(clk), .Q(new_AGEMA_signal_3661), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1385_s_current_state_reg ( .D(
        new_AGEMA_signal_3662), .CK(clk), .Q(new_AGEMA_signal_3663), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1387_s_current_state_reg ( .D(
        new_AGEMA_signal_3664), .CK(clk), .Q(new_AGEMA_signal_3665), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1389_s_current_state_reg ( .D(
        new_AGEMA_signal_3666), .CK(clk), .Q(new_AGEMA_signal_3667), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1391_s_current_state_reg ( .D(
        new_AGEMA_signal_3668), .CK(clk), .Q(new_AGEMA_signal_3669), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1393_s_current_state_reg ( .D(
        new_AGEMA_signal_3670), .CK(clk), .Q(new_AGEMA_signal_3671), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1395_s_current_state_reg ( .D(
        new_AGEMA_signal_3672), .CK(clk), .Q(new_AGEMA_signal_3673), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1397_s_current_state_reg ( .D(
        new_AGEMA_signal_3674), .CK(clk), .Q(new_AGEMA_signal_3675), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1399_s_current_state_reg ( .D(
        new_AGEMA_signal_3676), .CK(clk), .Q(new_AGEMA_signal_3677), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1401_s_current_state_reg ( .D(
        new_AGEMA_signal_3678), .CK(clk), .Q(new_AGEMA_signal_3679), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1403_s_current_state_reg ( .D(
        new_AGEMA_signal_3680), .CK(clk), .Q(new_AGEMA_signal_3681), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1405_s_current_state_reg ( .D(
        new_AGEMA_signal_3682), .CK(clk), .Q(new_AGEMA_signal_3683), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1407_s_current_state_reg ( .D(
        new_AGEMA_signal_3684), .CK(clk), .Q(new_AGEMA_signal_3685), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1409_s_current_state_reg ( .D(
        new_AGEMA_signal_3686), .CK(clk), .Q(new_AGEMA_signal_3687), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1411_s_current_state_reg ( .D(
        new_AGEMA_signal_3688), .CK(clk), .Q(new_AGEMA_signal_3689), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1413_s_current_state_reg ( .D(
        new_AGEMA_signal_3690), .CK(clk), .Q(new_AGEMA_signal_3691), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1415_s_current_state_reg ( .D(
        new_AGEMA_signal_3692), .CK(clk), .Q(new_AGEMA_signal_3693), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1417_s_current_state_reg ( .D(
        new_AGEMA_signal_3694), .CK(clk), .Q(new_AGEMA_signal_3695), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1419_s_current_state_reg ( .D(
        new_AGEMA_signal_3696), .CK(clk), .Q(new_AGEMA_signal_3697), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1421_s_current_state_reg ( .D(
        new_AGEMA_signal_3698), .CK(clk), .Q(new_AGEMA_signal_3699), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1423_s_current_state_reg ( .D(
        new_AGEMA_signal_3700), .CK(clk), .Q(new_AGEMA_signal_3701), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1425_s_current_state_reg ( .D(
        new_AGEMA_signal_3702), .CK(clk), .Q(new_AGEMA_signal_3703), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1427_s_current_state_reg ( .D(
        new_AGEMA_signal_3704), .CK(clk), .Q(new_AGEMA_signal_3705), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1429_s_current_state_reg ( .D(
        new_AGEMA_signal_3706), .CK(clk), .Q(new_AGEMA_signal_3707), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1431_s_current_state_reg ( .D(
        new_AGEMA_signal_3708), .CK(clk), .Q(new_AGEMA_signal_3709), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1433_s_current_state_reg ( .D(
        new_AGEMA_signal_3710), .CK(clk), .Q(new_AGEMA_signal_3711), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1435_s_current_state_reg ( .D(
        new_AGEMA_signal_3712), .CK(clk), .Q(new_AGEMA_signal_3713), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1437_s_current_state_reg ( .D(
        new_AGEMA_signal_3714), .CK(clk), .Q(new_AGEMA_signal_3715), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1439_s_current_state_reg ( .D(
        new_AGEMA_signal_3716), .CK(clk), .Q(new_AGEMA_signal_3717), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1441_s_current_state_reg ( .D(
        new_AGEMA_signal_3718), .CK(clk), .Q(new_AGEMA_signal_3719), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1443_s_current_state_reg ( .D(
        new_AGEMA_signal_3720), .CK(clk), .Q(new_AGEMA_signal_3721), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1445_s_current_state_reg ( .D(
        new_AGEMA_signal_3722), .CK(clk), .Q(new_AGEMA_signal_3723), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1447_s_current_state_reg ( .D(
        new_AGEMA_signal_3724), .CK(clk), .Q(new_AGEMA_signal_3725), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1449_s_current_state_reg ( .D(
        new_AGEMA_signal_3726), .CK(clk), .Q(new_AGEMA_signal_3727), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1451_s_current_state_reg ( .D(
        new_AGEMA_signal_3728), .CK(clk), .Q(new_AGEMA_signal_3729), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1453_s_current_state_reg ( .D(
        new_AGEMA_signal_3730), .CK(clk), .Q(new_AGEMA_signal_3731), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1455_s_current_state_reg ( .D(
        new_AGEMA_signal_3732), .CK(clk), .Q(new_AGEMA_signal_3733), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1457_s_current_state_reg ( .D(
        new_AGEMA_signal_3734), .CK(clk), .Q(new_AGEMA_signal_3735), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1459_s_current_state_reg ( .D(
        new_AGEMA_signal_3736), .CK(clk), .Q(new_AGEMA_signal_3737), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1461_s_current_state_reg ( .D(
        new_AGEMA_signal_3738), .CK(clk), .Q(new_AGEMA_signal_3739), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1463_s_current_state_reg ( .D(
        new_AGEMA_signal_3740), .CK(clk), .Q(new_AGEMA_signal_3741), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1465_s_current_state_reg ( .D(
        new_AGEMA_signal_3742), .CK(clk), .Q(new_AGEMA_signal_3743), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1467_s_current_state_reg ( .D(
        new_AGEMA_signal_3744), .CK(clk), .Q(new_AGEMA_signal_3745), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1469_s_current_state_reg ( .D(
        new_AGEMA_signal_3746), .CK(clk), .Q(new_AGEMA_signal_3747), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1471_s_current_state_reg ( .D(
        new_AGEMA_signal_3748), .CK(clk), .Q(new_AGEMA_signal_3749), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1473_s_current_state_reg ( .D(
        new_AGEMA_signal_3750), .CK(clk), .Q(new_AGEMA_signal_3751), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1475_s_current_state_reg ( .D(
        new_AGEMA_signal_3752), .CK(clk), .Q(new_AGEMA_signal_3753), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1477_s_current_state_reg ( .D(
        new_AGEMA_signal_3754), .CK(clk), .Q(new_AGEMA_signal_3755), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1479_s_current_state_reg ( .D(
        new_AGEMA_signal_3756), .CK(clk), .Q(new_AGEMA_signal_3757), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1481_s_current_state_reg ( .D(
        new_AGEMA_signal_3758), .CK(clk), .Q(new_AGEMA_signal_3759), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1483_s_current_state_reg ( .D(
        new_AGEMA_signal_3760), .CK(clk), .Q(new_AGEMA_signal_3761), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1485_s_current_state_reg ( .D(
        new_AGEMA_signal_3762), .CK(clk), .Q(new_AGEMA_signal_3763), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1487_s_current_state_reg ( .D(
        new_AGEMA_signal_3764), .CK(clk), .Q(new_AGEMA_signal_3765), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1489_s_current_state_reg ( .D(
        new_AGEMA_signal_3766), .CK(clk), .Q(new_AGEMA_signal_3767), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1491_s_current_state_reg ( .D(
        new_AGEMA_signal_3768), .CK(clk), .Q(new_AGEMA_signal_3769), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1493_s_current_state_reg ( .D(
        new_AGEMA_signal_3770), .CK(clk), .Q(new_AGEMA_signal_3771), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1495_s_current_state_reg ( .D(
        new_AGEMA_signal_3772), .CK(clk), .Q(new_AGEMA_signal_3773), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1497_s_current_state_reg ( .D(
        new_AGEMA_signal_3774), .CK(clk), .Q(new_AGEMA_signal_3775), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1499_s_current_state_reg ( .D(
        new_AGEMA_signal_3776), .CK(clk), .Q(new_AGEMA_signal_3777), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1501_s_current_state_reg ( .D(
        new_AGEMA_signal_3778), .CK(clk), .Q(new_AGEMA_signal_3779), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1503_s_current_state_reg ( .D(
        new_AGEMA_signal_3780), .CK(clk), .Q(new_AGEMA_signal_3781), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1505_s_current_state_reg ( .D(
        new_AGEMA_signal_3782), .CK(clk), .Q(new_AGEMA_signal_3783), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1507_s_current_state_reg ( .D(
        new_AGEMA_signal_3784), .CK(clk), .Q(new_AGEMA_signal_3785), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1509_s_current_state_reg ( .D(
        new_AGEMA_signal_3786), .CK(clk), .Q(new_AGEMA_signal_3787), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1511_s_current_state_reg ( .D(
        new_AGEMA_signal_3788), .CK(clk), .Q(new_AGEMA_signal_3789), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1513_s_current_state_reg ( .D(
        new_AGEMA_signal_3790), .CK(clk), .Q(new_AGEMA_signal_3791), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1515_s_current_state_reg ( .D(
        new_AGEMA_signal_3792), .CK(clk), .Q(new_AGEMA_signal_3793), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1517_s_current_state_reg ( .D(
        new_AGEMA_signal_3794), .CK(clk), .Q(new_AGEMA_signal_3795), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1519_s_current_state_reg ( .D(
        new_AGEMA_signal_3796), .CK(clk), .Q(new_AGEMA_signal_3797), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1521_s_current_state_reg ( .D(
        new_AGEMA_signal_3798), .CK(clk), .Q(new_AGEMA_signal_3799), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1523_s_current_state_reg ( .D(
        new_AGEMA_signal_3800), .CK(clk), .Q(new_AGEMA_signal_3801), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1525_s_current_state_reg ( .D(
        new_AGEMA_signal_3802), .CK(clk), .Q(new_AGEMA_signal_3803), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1527_s_current_state_reg ( .D(
        new_AGEMA_signal_3804), .CK(clk), .Q(new_AGEMA_signal_3805), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1529_s_current_state_reg ( .D(
        new_AGEMA_signal_3806), .CK(clk), .Q(new_AGEMA_signal_3807), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1531_s_current_state_reg ( .D(
        new_AGEMA_signal_3808), .CK(clk), .Q(new_AGEMA_signal_3809), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1533_s_current_state_reg ( .D(
        new_AGEMA_signal_3810), .CK(clk), .Q(new_AGEMA_signal_3811), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1535_s_current_state_reg ( .D(
        new_AGEMA_signal_3812), .CK(clk), .Q(new_AGEMA_signal_3813), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1537_s_current_state_reg ( .D(
        new_AGEMA_signal_3814), .CK(clk), .Q(new_AGEMA_signal_3815), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1539_s_current_state_reg ( .D(
        new_AGEMA_signal_3816), .CK(clk), .Q(new_AGEMA_signal_3817), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1541_s_current_state_reg ( .D(
        new_AGEMA_signal_3818), .CK(clk), .Q(new_AGEMA_signal_3819), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1543_s_current_state_reg ( .D(
        new_AGEMA_signal_3820), .CK(clk), .Q(new_AGEMA_signal_3821), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1545_s_current_state_reg ( .D(
        new_AGEMA_signal_3822), .CK(clk), .Q(new_AGEMA_signal_3823), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1547_s_current_state_reg ( .D(
        new_AGEMA_signal_3824), .CK(clk), .Q(new_AGEMA_signal_3825), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1549_s_current_state_reg ( .D(
        new_AGEMA_signal_3826), .CK(clk), .Q(new_AGEMA_signal_3827), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1551_s_current_state_reg ( .D(
        new_AGEMA_signal_3828), .CK(clk), .Q(new_AGEMA_signal_3829), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1553_s_current_state_reg ( .D(
        new_AGEMA_signal_3830), .CK(clk), .Q(new_AGEMA_signal_3831), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1555_s_current_state_reg ( .D(
        new_AGEMA_signal_3832), .CK(clk), .Q(new_AGEMA_signal_3833), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1557_s_current_state_reg ( .D(
        new_AGEMA_signal_3834), .CK(clk), .Q(new_AGEMA_signal_3835), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1559_s_current_state_reg ( .D(
        new_AGEMA_signal_3836), .CK(clk), .Q(new_AGEMA_signal_3837), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1561_s_current_state_reg ( .D(
        new_AGEMA_signal_3838), .CK(clk), .Q(new_AGEMA_signal_3839), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1563_s_current_state_reg ( .D(
        new_AGEMA_signal_3840), .CK(clk), .Q(new_AGEMA_signal_3841), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1565_s_current_state_reg ( .D(
        new_AGEMA_signal_3842), .CK(clk), .Q(new_AGEMA_signal_3843), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1567_s_current_state_reg ( .D(
        new_AGEMA_signal_3844), .CK(clk), .Q(new_AGEMA_signal_3845), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1569_s_current_state_reg ( .D(
        new_AGEMA_signal_3846), .CK(clk), .Q(new_AGEMA_signal_3847), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1571_s_current_state_reg ( .D(
        new_AGEMA_signal_3848), .CK(clk), .Q(new_AGEMA_signal_3849), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1573_s_current_state_reg ( .D(
        new_AGEMA_signal_3850), .CK(clk), .Q(new_AGEMA_signal_3851), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1575_s_current_state_reg ( .D(
        new_AGEMA_signal_3852), .CK(clk), .Q(new_AGEMA_signal_3853), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1577_s_current_state_reg ( .D(
        new_AGEMA_signal_3854), .CK(clk), .Q(new_AGEMA_signal_3855), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1579_s_current_state_reg ( .D(
        new_AGEMA_signal_3856), .CK(clk), .Q(new_AGEMA_signal_3857), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1581_s_current_state_reg ( .D(
        new_AGEMA_signal_3858), .CK(clk), .Q(new_AGEMA_signal_3859), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1583_s_current_state_reg ( .D(
        new_AGEMA_signal_3860), .CK(clk), .Q(new_AGEMA_signal_3861), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1585_s_current_state_reg ( .D(
        new_AGEMA_signal_3862), .CK(clk), .Q(new_AGEMA_signal_3863), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1587_s_current_state_reg ( .D(
        new_AGEMA_signal_3864), .CK(clk), .Q(new_AGEMA_signal_3865), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1589_s_current_state_reg ( .D(
        new_AGEMA_signal_3866), .CK(clk), .Q(new_AGEMA_signal_3867), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1591_s_current_state_reg ( .D(
        new_AGEMA_signal_3868), .CK(clk), .Q(new_AGEMA_signal_3869), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1593_s_current_state_reg ( .D(
        new_AGEMA_signal_3870), .CK(clk), .Q(new_AGEMA_signal_3871), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1595_s_current_state_reg ( .D(
        new_AGEMA_signal_3872), .CK(clk), .Q(new_AGEMA_signal_3873), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1597_s_current_state_reg ( .D(
        new_AGEMA_signal_3874), .CK(clk), .Q(new_AGEMA_signal_3875), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1599_s_current_state_reg ( .D(
        new_AGEMA_signal_3876), .CK(clk), .Q(new_AGEMA_signal_3877), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1601_s_current_state_reg ( .D(
        new_AGEMA_signal_3878), .CK(clk), .Q(new_AGEMA_signal_3879), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1603_s_current_state_reg ( .D(
        new_AGEMA_signal_3880), .CK(clk), .Q(new_AGEMA_signal_3881), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1605_s_current_state_reg ( .D(
        new_AGEMA_signal_3882), .CK(clk), .Q(new_AGEMA_signal_3883), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1607_s_current_state_reg ( .D(
        new_AGEMA_signal_3884), .CK(clk), .Q(new_AGEMA_signal_3885), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1609_s_current_state_reg ( .D(
        new_AGEMA_signal_3886), .CK(clk), .Q(new_AGEMA_signal_3887), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1611_s_current_state_reg ( .D(
        new_AGEMA_signal_3888), .CK(clk), .Q(new_AGEMA_signal_3889), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1613_s_current_state_reg ( .D(
        new_AGEMA_signal_3890), .CK(clk), .Q(new_AGEMA_signal_3891), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1615_s_current_state_reg ( .D(
        new_AGEMA_signal_3892), .CK(clk), .Q(new_AGEMA_signal_3893), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1617_s_current_state_reg ( .D(
        new_AGEMA_signal_3894), .CK(clk), .Q(new_AGEMA_signal_3895), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1619_s_current_state_reg ( .D(
        new_AGEMA_signal_3896), .CK(clk), .Q(new_AGEMA_signal_3897), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1621_s_current_state_reg ( .D(
        new_AGEMA_signal_3898), .CK(clk), .Q(new_AGEMA_signal_3899), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1623_s_current_state_reg ( .D(
        new_AGEMA_signal_3900), .CK(clk), .Q(new_AGEMA_signal_3901), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1625_s_current_state_reg ( .D(
        new_AGEMA_signal_3902), .CK(clk), .Q(new_AGEMA_signal_3903), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1627_s_current_state_reg ( .D(
        new_AGEMA_signal_3904), .CK(clk), .Q(new_AGEMA_signal_3905), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1629_s_current_state_reg ( .D(
        new_AGEMA_signal_3906), .CK(clk), .Q(new_AGEMA_signal_3907), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1631_s_current_state_reg ( .D(
        new_AGEMA_signal_3908), .CK(clk), .Q(new_AGEMA_signal_3909), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1633_s_current_state_reg ( .D(
        new_AGEMA_signal_3910), .CK(clk), .Q(new_AGEMA_signal_3911), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1635_s_current_state_reg ( .D(
        new_AGEMA_signal_3912), .CK(clk), .Q(new_AGEMA_signal_3913), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1637_s_current_state_reg ( .D(
        new_AGEMA_signal_3914), .CK(clk), .Q(new_AGEMA_signal_3915), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1639_s_current_state_reg ( .D(
        new_AGEMA_signal_3916), .CK(clk), .Q(new_AGEMA_signal_3917), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1641_s_current_state_reg ( .D(
        new_AGEMA_signal_3918), .CK(clk), .Q(new_AGEMA_signal_3919), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1643_s_current_state_reg ( .D(
        new_AGEMA_signal_3920), .CK(clk), .Q(new_AGEMA_signal_3921), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1645_s_current_state_reg ( .D(
        new_AGEMA_signal_3922), .CK(clk), .Q(new_AGEMA_signal_3923), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1647_s_current_state_reg ( .D(
        new_AGEMA_signal_3924), .CK(clk), .Q(new_AGEMA_signal_3925), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1649_s_current_state_reg ( .D(
        new_AGEMA_signal_3926), .CK(clk), .Q(new_AGEMA_signal_3927), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1651_s_current_state_reg ( .D(
        new_AGEMA_signal_3928), .CK(clk), .Q(new_AGEMA_signal_3929), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1653_s_current_state_reg ( .D(
        new_AGEMA_signal_3930), .CK(clk), .Q(new_AGEMA_signal_3931), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1655_s_current_state_reg ( .D(
        new_AGEMA_signal_3932), .CK(clk), .Q(new_AGEMA_signal_3933), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1657_s_current_state_reg ( .D(
        new_AGEMA_signal_3934), .CK(clk), .Q(new_AGEMA_signal_3935), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1659_s_current_state_reg ( .D(
        new_AGEMA_signal_3936), .CK(clk), .Q(new_AGEMA_signal_3937), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1661_s_current_state_reg ( .D(
        new_AGEMA_signal_3938), .CK(clk), .Q(new_AGEMA_signal_3939), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1663_s_current_state_reg ( .D(
        new_AGEMA_signal_3940), .CK(clk), .Q(new_AGEMA_signal_3941), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1665_s_current_state_reg ( .D(
        new_AGEMA_signal_3942), .CK(clk), .Q(new_AGEMA_signal_3943), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1667_s_current_state_reg ( .D(
        new_AGEMA_signal_3944), .CK(clk), .Q(new_AGEMA_signal_3945), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1669_s_current_state_reg ( .D(
        new_AGEMA_signal_3946), .CK(clk), .Q(new_AGEMA_signal_3947), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1671_s_current_state_reg ( .D(
        new_AGEMA_signal_3948), .CK(clk), .Q(new_AGEMA_signal_3949), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1673_s_current_state_reg ( .D(
        new_AGEMA_signal_3950), .CK(clk), .Q(new_AGEMA_signal_3951), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1675_s_current_state_reg ( .D(
        new_AGEMA_signal_3952), .CK(clk), .Q(new_AGEMA_signal_3953), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1677_s_current_state_reg ( .D(
        new_AGEMA_signal_3954), .CK(clk), .Q(new_AGEMA_signal_3955), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1681_s_current_state_reg ( .D(
        new_AGEMA_signal_3958), .CK(clk), .Q(new_AGEMA_signal_3959), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1685_s_current_state_reg ( .D(
        new_AGEMA_signal_3962), .CK(clk), .Q(new_AGEMA_signal_3963), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1689_s_current_state_reg ( .D(
        new_AGEMA_signal_3966), .CK(clk), .Q(new_AGEMA_signal_3967), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1693_s_current_state_reg ( .D(
        new_AGEMA_signal_3970), .CK(clk), .Q(new_AGEMA_signal_3971), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1697_s_current_state_reg ( .D(
        new_AGEMA_signal_3974), .CK(clk), .Q(new_AGEMA_signal_3975), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1701_s_current_state_reg ( .D(
        new_AGEMA_signal_3978), .CK(clk), .Q(new_AGEMA_signal_3979), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1705_s_current_state_reg ( .D(
        new_AGEMA_signal_3982), .CK(clk), .Q(new_AGEMA_signal_3983), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1709_s_current_state_reg ( .D(
        new_AGEMA_signal_3986), .CK(clk), .Q(new_AGEMA_signal_3987), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1713_s_current_state_reg ( .D(
        new_AGEMA_signal_3990), .CK(clk), .Q(new_AGEMA_signal_3991), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1717_s_current_state_reg ( .D(
        new_AGEMA_signal_3994), .CK(clk), .Q(new_AGEMA_signal_3995), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1721_s_current_state_reg ( .D(
        new_AGEMA_signal_3998), .CK(clk), .Q(new_AGEMA_signal_3999), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1725_s_current_state_reg ( .D(
        new_AGEMA_signal_4002), .CK(clk), .Q(new_AGEMA_signal_4003), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1729_s_current_state_reg ( .D(
        new_AGEMA_signal_4006), .CK(clk), .Q(new_AGEMA_signal_4007), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1733_s_current_state_reg ( .D(
        new_AGEMA_signal_4010), .CK(clk), .Q(new_AGEMA_signal_4011), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1737_s_current_state_reg ( .D(
        new_AGEMA_signal_4014), .CK(clk), .Q(new_AGEMA_signal_4015), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1741_s_current_state_reg ( .D(
        new_AGEMA_signal_4018), .CK(clk), .Q(new_AGEMA_signal_4019), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1745_s_current_state_reg ( .D(
        new_AGEMA_signal_4022), .CK(clk), .Q(new_AGEMA_signal_4023), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1749_s_current_state_reg ( .D(
        new_AGEMA_signal_4026), .CK(clk), .Q(new_AGEMA_signal_4027), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1753_s_current_state_reg ( .D(
        new_AGEMA_signal_4030), .CK(clk), .Q(new_AGEMA_signal_4031), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1757_s_current_state_reg ( .D(
        new_AGEMA_signal_4034), .CK(clk), .Q(new_AGEMA_signal_4035), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1761_s_current_state_reg ( .D(
        new_AGEMA_signal_4038), .CK(clk), .Q(new_AGEMA_signal_4039), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1765_s_current_state_reg ( .D(
        new_AGEMA_signal_4042), .CK(clk), .Q(new_AGEMA_signal_4043), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1769_s_current_state_reg ( .D(
        new_AGEMA_signal_4046), .CK(clk), .Q(new_AGEMA_signal_4047), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1773_s_current_state_reg ( .D(
        new_AGEMA_signal_4050), .CK(clk), .Q(new_AGEMA_signal_4051), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1777_s_current_state_reg ( .D(
        new_AGEMA_signal_4054), .CK(clk), .Q(new_AGEMA_signal_4055), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1781_s_current_state_reg ( .D(
        new_AGEMA_signal_4058), .CK(clk), .Q(new_AGEMA_signal_4059), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1785_s_current_state_reg ( .D(
        new_AGEMA_signal_4062), .CK(clk), .Q(new_AGEMA_signal_4063), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1789_s_current_state_reg ( .D(
        new_AGEMA_signal_4066), .CK(clk), .Q(new_AGEMA_signal_4067), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1793_s_current_state_reg ( .D(
        new_AGEMA_signal_4070), .CK(clk), .Q(new_AGEMA_signal_4071), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1797_s_current_state_reg ( .D(
        new_AGEMA_signal_4074), .CK(clk), .Q(new_AGEMA_signal_4075), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1801_s_current_state_reg ( .D(
        new_AGEMA_signal_4078), .CK(clk), .Q(new_AGEMA_signal_4079), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1805_s_current_state_reg ( .D(
        new_AGEMA_signal_4082), .CK(clk), .Q(new_AGEMA_signal_4083), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1809_s_current_state_reg ( .D(
        new_AGEMA_signal_4086), .CK(clk), .Q(new_AGEMA_signal_4087), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1813_s_current_state_reg ( .D(
        new_AGEMA_signal_4090), .CK(clk), .Q(new_AGEMA_signal_4091), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1817_s_current_state_reg ( .D(
        new_AGEMA_signal_4094), .CK(clk), .Q(new_AGEMA_signal_4095), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1821_s_current_state_reg ( .D(
        new_AGEMA_signal_4098), .CK(clk), .Q(new_AGEMA_signal_4099), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1825_s_current_state_reg ( .D(
        new_AGEMA_signal_4102), .CK(clk), .Q(new_AGEMA_signal_4103), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1829_s_current_state_reg ( .D(
        new_AGEMA_signal_4106), .CK(clk), .Q(new_AGEMA_signal_4107), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1833_s_current_state_reg ( .D(
        new_AGEMA_signal_4110), .CK(clk), .Q(new_AGEMA_signal_4111), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1837_s_current_state_reg ( .D(
        new_AGEMA_signal_4114), .CK(clk), .Q(new_AGEMA_signal_4115), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1841_s_current_state_reg ( .D(
        new_AGEMA_signal_4118), .CK(clk), .Q(new_AGEMA_signal_4119), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1845_s_current_state_reg ( .D(
        new_AGEMA_signal_4122), .CK(clk), .Q(new_AGEMA_signal_4123), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1849_s_current_state_reg ( .D(
        new_AGEMA_signal_4126), .CK(clk), .Q(new_AGEMA_signal_4127), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1853_s_current_state_reg ( .D(
        new_AGEMA_signal_4130), .CK(clk), .Q(new_AGEMA_signal_4131), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1857_s_current_state_reg ( .D(
        new_AGEMA_signal_4134), .CK(clk), .Q(new_AGEMA_signal_4135), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1861_s_current_state_reg ( .D(
        new_AGEMA_signal_4138), .CK(clk), .Q(new_AGEMA_signal_4139), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1865_s_current_state_reg ( .D(
        new_AGEMA_signal_4142), .CK(clk), .Q(new_AGEMA_signal_4143), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1869_s_current_state_reg ( .D(
        new_AGEMA_signal_4146), .CK(clk), .Q(new_AGEMA_signal_4147), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1873_s_current_state_reg ( .D(
        new_AGEMA_signal_4150), .CK(clk), .Q(new_AGEMA_signal_4151), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1877_s_current_state_reg ( .D(
        new_AGEMA_signal_4154), .CK(clk), .Q(new_AGEMA_signal_4155), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1881_s_current_state_reg ( .D(
        new_AGEMA_signal_4158), .CK(clk), .Q(new_AGEMA_signal_4159), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1885_s_current_state_reg ( .D(
        new_AGEMA_signal_4162), .CK(clk), .Q(new_AGEMA_signal_4163), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1889_s_current_state_reg ( .D(
        new_AGEMA_signal_4166), .CK(clk), .Q(new_AGEMA_signal_4167), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1893_s_current_state_reg ( .D(
        new_AGEMA_signal_4170), .CK(clk), .Q(new_AGEMA_signal_4171), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1897_s_current_state_reg ( .D(
        new_AGEMA_signal_4174), .CK(clk), .Q(new_AGEMA_signal_4175), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1901_s_current_state_reg ( .D(
        new_AGEMA_signal_4178), .CK(clk), .Q(new_AGEMA_signal_4179), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1905_s_current_state_reg ( .D(
        new_AGEMA_signal_4182), .CK(clk), .Q(new_AGEMA_signal_4183), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1909_s_current_state_reg ( .D(
        new_AGEMA_signal_4186), .CK(clk), .Q(new_AGEMA_signal_4187), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1913_s_current_state_reg ( .D(
        new_AGEMA_signal_4190), .CK(clk), .Q(new_AGEMA_signal_4191), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1917_s_current_state_reg ( .D(
        new_AGEMA_signal_4194), .CK(clk), .Q(new_AGEMA_signal_4195), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1921_s_current_state_reg ( .D(
        new_AGEMA_signal_4198), .CK(clk), .Q(new_AGEMA_signal_4199), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1925_s_current_state_reg ( .D(
        new_AGEMA_signal_4202), .CK(clk), .Q(new_AGEMA_signal_4203), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1929_s_current_state_reg ( .D(
        new_AGEMA_signal_4206), .CK(clk), .Q(new_AGEMA_signal_4207), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1933_s_current_state_reg ( .D(
        new_AGEMA_signal_4210), .CK(clk), .Q(new_AGEMA_signal_4211), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1937_s_current_state_reg ( .D(
        new_AGEMA_signal_4214), .CK(clk), .Q(new_AGEMA_signal_4215), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1941_s_current_state_reg ( .D(
        new_AGEMA_signal_4218), .CK(clk), .Q(new_AGEMA_signal_4219), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1945_s_current_state_reg ( .D(
        new_AGEMA_signal_4222), .CK(clk), .Q(new_AGEMA_signal_4223), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1949_s_current_state_reg ( .D(
        new_AGEMA_signal_4226), .CK(clk), .Q(new_AGEMA_signal_4227), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1953_s_current_state_reg ( .D(
        new_AGEMA_signal_4230), .CK(clk), .Q(new_AGEMA_signal_4231), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1957_s_current_state_reg ( .D(
        new_AGEMA_signal_4234), .CK(clk), .Q(new_AGEMA_signal_4235), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1961_s_current_state_reg ( .D(
        new_AGEMA_signal_4238), .CK(clk), .Q(new_AGEMA_signal_4239), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1965_s_current_state_reg ( .D(
        new_AGEMA_signal_4242), .CK(clk), .Q(new_AGEMA_signal_4243), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1969_s_current_state_reg ( .D(
        new_AGEMA_signal_4246), .CK(clk), .Q(new_AGEMA_signal_4247), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1973_s_current_state_reg ( .D(
        new_AGEMA_signal_4250), .CK(clk), .Q(new_AGEMA_signal_4251), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1977_s_current_state_reg ( .D(
        new_AGEMA_signal_4254), .CK(clk), .Q(new_AGEMA_signal_4255), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1981_s_current_state_reg ( .D(
        new_AGEMA_signal_4258), .CK(clk), .Q(new_AGEMA_signal_4259), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1985_s_current_state_reg ( .D(
        new_AGEMA_signal_4262), .CK(clk), .Q(new_AGEMA_signal_4263), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1989_s_current_state_reg ( .D(
        new_AGEMA_signal_4266), .CK(clk), .Q(new_AGEMA_signal_4267), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1993_s_current_state_reg ( .D(
        new_AGEMA_signal_4270), .CK(clk), .Q(new_AGEMA_signal_4271), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1997_s_current_state_reg ( .D(
        new_AGEMA_signal_4274), .CK(clk), .Q(new_AGEMA_signal_4275), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2001_s_current_state_reg ( .D(
        new_AGEMA_signal_4278), .CK(clk), .Q(new_AGEMA_signal_4279), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2005_s_current_state_reg ( .D(
        new_AGEMA_signal_4282), .CK(clk), .Q(new_AGEMA_signal_4283), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2009_s_current_state_reg ( .D(
        new_AGEMA_signal_4286), .CK(clk), .Q(new_AGEMA_signal_4287), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2013_s_current_state_reg ( .D(
        new_AGEMA_signal_4290), .CK(clk), .Q(new_AGEMA_signal_4291), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2017_s_current_state_reg ( .D(
        new_AGEMA_signal_4294), .CK(clk), .Q(new_AGEMA_signal_4295), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2021_s_current_state_reg ( .D(
        new_AGEMA_signal_4298), .CK(clk), .Q(new_AGEMA_signal_4299), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2025_s_current_state_reg ( .D(
        new_AGEMA_signal_4302), .CK(clk), .Q(new_AGEMA_signal_4303), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2029_s_current_state_reg ( .D(
        new_AGEMA_signal_4306), .CK(clk), .Q(new_AGEMA_signal_4307), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2033_s_current_state_reg ( .D(
        new_AGEMA_signal_4310), .CK(clk), .Q(new_AGEMA_signal_4311), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2037_s_current_state_reg ( .D(
        new_AGEMA_signal_4314), .CK(clk), .Q(new_AGEMA_signal_4315), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2041_s_current_state_reg ( .D(
        new_AGEMA_signal_4318), .CK(clk), .Q(new_AGEMA_signal_4319), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2045_s_current_state_reg ( .D(
        new_AGEMA_signal_4322), .CK(clk), .Q(new_AGEMA_signal_4323), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2049_s_current_state_reg ( .D(
        new_AGEMA_signal_4326), .CK(clk), .Q(new_AGEMA_signal_4327), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2053_s_current_state_reg ( .D(
        new_AGEMA_signal_4330), .CK(clk), .Q(new_AGEMA_signal_4331), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2057_s_current_state_reg ( .D(
        new_AGEMA_signal_4334), .CK(clk), .Q(new_AGEMA_signal_4335), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2061_s_current_state_reg ( .D(
        new_AGEMA_signal_4338), .CK(clk), .Q(new_AGEMA_signal_4339), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2065_s_current_state_reg ( .D(
        new_AGEMA_signal_4342), .CK(clk), .Q(new_AGEMA_signal_4343), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2067_s_current_state_reg ( .D(
        new_AGEMA_signal_4344), .CK(clk), .Q(new_AGEMA_signal_4345), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2069_s_current_state_reg ( .D(
        new_AGEMA_signal_4346), .CK(clk), .Q(new_AGEMA_signal_4347), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2077_s_current_state_reg ( .D(
        new_AGEMA_signal_4354), .CK(clk), .Q(new_AGEMA_signal_4355), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2079_s_current_state_reg ( .D(
        new_AGEMA_signal_4356), .CK(clk), .Q(new_AGEMA_signal_4357), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2081_s_current_state_reg ( .D(
        new_AGEMA_signal_4358), .CK(clk), .Q(new_AGEMA_signal_4359), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2083_s_current_state_reg ( .D(
        new_AGEMA_signal_4360), .CK(clk), .Q(new_AGEMA_signal_4361), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2087_s_current_state_reg ( .D(
        new_AGEMA_signal_4364), .CK(clk), .Q(new_AGEMA_signal_4365), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2091_s_current_state_reg ( .D(
        new_AGEMA_signal_4368), .CK(clk), .Q(new_AGEMA_signal_4369), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2101_s_current_state_reg ( .D(
        new_AGEMA_signal_4378), .CK(clk), .Q(new_AGEMA_signal_4379), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2103_s_current_state_reg ( .D(
        new_AGEMA_signal_4380), .CK(clk), .Q(new_AGEMA_signal_4381), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2105_s_current_state_reg ( .D(
        new_AGEMA_signal_4382), .CK(clk), .Q(new_AGEMA_signal_4383), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2113_s_current_state_reg ( .D(
        new_AGEMA_signal_4390), .CK(clk), .Q(new_AGEMA_signal_4391), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2115_s_current_state_reg ( .D(
        new_AGEMA_signal_4392), .CK(clk), .Q(new_AGEMA_signal_4393), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2117_s_current_state_reg ( .D(
        new_AGEMA_signal_4394), .CK(clk), .Q(new_AGEMA_signal_4395), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2119_s_current_state_reg ( .D(
        new_AGEMA_signal_4396), .CK(clk), .Q(new_AGEMA_signal_4397), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2123_s_current_state_reg ( .D(
        new_AGEMA_signal_4400), .CK(clk), .Q(new_AGEMA_signal_4401), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2127_s_current_state_reg ( .D(
        new_AGEMA_signal_4404), .CK(clk), .Q(new_AGEMA_signal_4405), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2137_s_current_state_reg ( .D(
        new_AGEMA_signal_4414), .CK(clk), .Q(new_AGEMA_signal_4415), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2139_s_current_state_reg ( .D(
        new_AGEMA_signal_4416), .CK(clk), .Q(new_AGEMA_signal_4417), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2141_s_current_state_reg ( .D(
        new_AGEMA_signal_4418), .CK(clk), .Q(new_AGEMA_signal_4419), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2149_s_current_state_reg ( .D(
        new_AGEMA_signal_4426), .CK(clk), .Q(new_AGEMA_signal_4427), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2151_s_current_state_reg ( .D(
        new_AGEMA_signal_4428), .CK(clk), .Q(new_AGEMA_signal_4429), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2153_s_current_state_reg ( .D(
        new_AGEMA_signal_4430), .CK(clk), .Q(new_AGEMA_signal_4431), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2155_s_current_state_reg ( .D(
        new_AGEMA_signal_4432), .CK(clk), .Q(new_AGEMA_signal_4433), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2159_s_current_state_reg ( .D(
        new_AGEMA_signal_4436), .CK(clk), .Q(new_AGEMA_signal_4437), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2163_s_current_state_reg ( .D(
        new_AGEMA_signal_4440), .CK(clk), .Q(new_AGEMA_signal_4441), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2173_s_current_state_reg ( .D(
        new_AGEMA_signal_4450), .CK(clk), .Q(new_AGEMA_signal_4451), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2175_s_current_state_reg ( .D(
        new_AGEMA_signal_4452), .CK(clk), .Q(new_AGEMA_signal_4453), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2177_s_current_state_reg ( .D(
        new_AGEMA_signal_4454), .CK(clk), .Q(new_AGEMA_signal_4455), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2185_s_current_state_reg ( .D(
        new_AGEMA_signal_4462), .CK(clk), .Q(new_AGEMA_signal_4463), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2187_s_current_state_reg ( .D(
        new_AGEMA_signal_4464), .CK(clk), .Q(new_AGEMA_signal_4465), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2189_s_current_state_reg ( .D(
        new_AGEMA_signal_4466), .CK(clk), .Q(new_AGEMA_signal_4467), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2191_s_current_state_reg ( .D(
        new_AGEMA_signal_4468), .CK(clk), .Q(new_AGEMA_signal_4469), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2195_s_current_state_reg ( .D(
        new_AGEMA_signal_4472), .CK(clk), .Q(new_AGEMA_signal_4473), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2199_s_current_state_reg ( .D(
        new_AGEMA_signal_4476), .CK(clk), .Q(new_AGEMA_signal_4477), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2209_s_current_state_reg ( .D(
        new_AGEMA_signal_4486), .CK(clk), .Q(new_AGEMA_signal_4487), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2211_s_current_state_reg ( .D(
        new_AGEMA_signal_4488), .CK(clk), .Q(new_AGEMA_signal_4489), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2213_s_current_state_reg ( .D(
        new_AGEMA_signal_4490), .CK(clk), .Q(new_AGEMA_signal_4491), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2221_s_current_state_reg ( .D(
        new_AGEMA_signal_4498), .CK(clk), .Q(new_AGEMA_signal_4499), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2223_s_current_state_reg ( .D(
        new_AGEMA_signal_4500), .CK(clk), .Q(new_AGEMA_signal_4501), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2225_s_current_state_reg ( .D(
        new_AGEMA_signal_4502), .CK(clk), .Q(new_AGEMA_signal_4503), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2227_s_current_state_reg ( .D(
        new_AGEMA_signal_4504), .CK(clk), .Q(new_AGEMA_signal_4505), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2231_s_current_state_reg ( .D(
        new_AGEMA_signal_4508), .CK(clk), .Q(new_AGEMA_signal_4509), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2235_s_current_state_reg ( .D(
        new_AGEMA_signal_4512), .CK(clk), .Q(new_AGEMA_signal_4513), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2245_s_current_state_reg ( .D(
        new_AGEMA_signal_4522), .CK(clk), .Q(new_AGEMA_signal_4523), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2247_s_current_state_reg ( .D(
        new_AGEMA_signal_4524), .CK(clk), .Q(new_AGEMA_signal_4525), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2249_s_current_state_reg ( .D(
        new_AGEMA_signal_4526), .CK(clk), .Q(new_AGEMA_signal_4527), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2257_s_current_state_reg ( .D(
        new_AGEMA_signal_4534), .CK(clk), .Q(new_AGEMA_signal_4535), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2259_s_current_state_reg ( .D(
        new_AGEMA_signal_4536), .CK(clk), .Q(new_AGEMA_signal_4537), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2261_s_current_state_reg ( .D(
        new_AGEMA_signal_4538), .CK(clk), .Q(new_AGEMA_signal_4539), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2263_s_current_state_reg ( .D(
        new_AGEMA_signal_4540), .CK(clk), .Q(new_AGEMA_signal_4541), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2267_s_current_state_reg ( .D(
        new_AGEMA_signal_4544), .CK(clk), .Q(new_AGEMA_signal_4545), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2271_s_current_state_reg ( .D(
        new_AGEMA_signal_4548), .CK(clk), .Q(new_AGEMA_signal_4549), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2281_s_current_state_reg ( .D(
        new_AGEMA_signal_4558), .CK(clk), .Q(new_AGEMA_signal_4559), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2283_s_current_state_reg ( .D(
        new_AGEMA_signal_4560), .CK(clk), .Q(new_AGEMA_signal_4561), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2285_s_current_state_reg ( .D(
        new_AGEMA_signal_4562), .CK(clk), .Q(new_AGEMA_signal_4563), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2293_s_current_state_reg ( .D(
        new_AGEMA_signal_4570), .CK(clk), .Q(new_AGEMA_signal_4571), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2295_s_current_state_reg ( .D(
        new_AGEMA_signal_4572), .CK(clk), .Q(new_AGEMA_signal_4573), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2297_s_current_state_reg ( .D(
        new_AGEMA_signal_4574), .CK(clk), .Q(new_AGEMA_signal_4575), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2299_s_current_state_reg ( .D(
        new_AGEMA_signal_4576), .CK(clk), .Q(new_AGEMA_signal_4577), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2303_s_current_state_reg ( .D(
        new_AGEMA_signal_4580), .CK(clk), .Q(new_AGEMA_signal_4581), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2307_s_current_state_reg ( .D(
        new_AGEMA_signal_4584), .CK(clk), .Q(new_AGEMA_signal_4585), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2317_s_current_state_reg ( .D(
        new_AGEMA_signal_4594), .CK(clk), .Q(new_AGEMA_signal_4595), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2319_s_current_state_reg ( .D(
        new_AGEMA_signal_4596), .CK(clk), .Q(new_AGEMA_signal_4597), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2321_s_current_state_reg ( .D(
        new_AGEMA_signal_4598), .CK(clk), .Q(new_AGEMA_signal_4599), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2329_s_current_state_reg ( .D(
        new_AGEMA_signal_4606), .CK(clk), .Q(new_AGEMA_signal_4607), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2331_s_current_state_reg ( .D(
        new_AGEMA_signal_4608), .CK(clk), .Q(new_AGEMA_signal_4609), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2333_s_current_state_reg ( .D(
        new_AGEMA_signal_4610), .CK(clk), .Q(new_AGEMA_signal_4611), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2335_s_current_state_reg ( .D(
        new_AGEMA_signal_4612), .CK(clk), .Q(new_AGEMA_signal_4613), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2339_s_current_state_reg ( .D(
        new_AGEMA_signal_4616), .CK(clk), .Q(new_AGEMA_signal_4617), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2343_s_current_state_reg ( .D(
        new_AGEMA_signal_4620), .CK(clk), .Q(new_AGEMA_signal_4621), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2353_s_current_state_reg ( .D(
        new_AGEMA_signal_4630), .CK(clk), .Q(new_AGEMA_signal_4631), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2355_s_current_state_reg ( .D(
        new_AGEMA_signal_4632), .CK(clk), .Q(new_AGEMA_signal_4633), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2357_s_current_state_reg ( .D(
        new_AGEMA_signal_4634), .CK(clk), .Q(new_AGEMA_signal_4635), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2365_s_current_state_reg ( .D(
        new_AGEMA_signal_4642), .CK(clk), .Q(new_AGEMA_signal_4643), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2367_s_current_state_reg ( .D(
        new_AGEMA_signal_4644), .CK(clk), .Q(new_AGEMA_signal_4645), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2369_s_current_state_reg ( .D(
        new_AGEMA_signal_4646), .CK(clk), .Q(new_AGEMA_signal_4647), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2371_s_current_state_reg ( .D(
        new_AGEMA_signal_4648), .CK(clk), .Q(new_AGEMA_signal_4649), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2375_s_current_state_reg ( .D(
        new_AGEMA_signal_4652), .CK(clk), .Q(new_AGEMA_signal_4653), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2379_s_current_state_reg ( .D(
        new_AGEMA_signal_4656), .CK(clk), .Q(new_AGEMA_signal_4657), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2389_s_current_state_reg ( .D(
        new_AGEMA_signal_4666), .CK(clk), .Q(new_AGEMA_signal_4667), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2391_s_current_state_reg ( .D(
        new_AGEMA_signal_4668), .CK(clk), .Q(new_AGEMA_signal_4669), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2393_s_current_state_reg ( .D(
        new_AGEMA_signal_4670), .CK(clk), .Q(new_AGEMA_signal_4671), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2401_s_current_state_reg ( .D(
        new_AGEMA_signal_4678), .CK(clk), .Q(new_AGEMA_signal_4679), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2403_s_current_state_reg ( .D(
        new_AGEMA_signal_4680), .CK(clk), .Q(new_AGEMA_signal_4681), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2405_s_current_state_reg ( .D(
        new_AGEMA_signal_4682), .CK(clk), .Q(new_AGEMA_signal_4683), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2407_s_current_state_reg ( .D(
        new_AGEMA_signal_4684), .CK(clk), .Q(new_AGEMA_signal_4685), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2411_s_current_state_reg ( .D(
        new_AGEMA_signal_4688), .CK(clk), .Q(new_AGEMA_signal_4689), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2415_s_current_state_reg ( .D(
        new_AGEMA_signal_4692), .CK(clk), .Q(new_AGEMA_signal_4693), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2425_s_current_state_reg ( .D(
        new_AGEMA_signal_4702), .CK(clk), .Q(new_AGEMA_signal_4703), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2427_s_current_state_reg ( .D(
        new_AGEMA_signal_4704), .CK(clk), .Q(new_AGEMA_signal_4705), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2429_s_current_state_reg ( .D(
        new_AGEMA_signal_4706), .CK(clk), .Q(new_AGEMA_signal_4707), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2437_s_current_state_reg ( .D(
        new_AGEMA_signal_4714), .CK(clk), .Q(new_AGEMA_signal_4715), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2439_s_current_state_reg ( .D(
        new_AGEMA_signal_4716), .CK(clk), .Q(new_AGEMA_signal_4717), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2441_s_current_state_reg ( .D(
        new_AGEMA_signal_4718), .CK(clk), .Q(new_AGEMA_signal_4719), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2443_s_current_state_reg ( .D(
        new_AGEMA_signal_4720), .CK(clk), .Q(new_AGEMA_signal_4721), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2447_s_current_state_reg ( .D(
        new_AGEMA_signal_4724), .CK(clk), .Q(new_AGEMA_signal_4725), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2451_s_current_state_reg ( .D(
        new_AGEMA_signal_4728), .CK(clk), .Q(new_AGEMA_signal_4729), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2461_s_current_state_reg ( .D(
        new_AGEMA_signal_4738), .CK(clk), .Q(new_AGEMA_signal_4739), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2463_s_current_state_reg ( .D(
        new_AGEMA_signal_4740), .CK(clk), .Q(new_AGEMA_signal_4741), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2465_s_current_state_reg ( .D(
        new_AGEMA_signal_4742), .CK(clk), .Q(new_AGEMA_signal_4743), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2473_s_current_state_reg ( .D(
        new_AGEMA_signal_4750), .CK(clk), .Q(new_AGEMA_signal_4751), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2475_s_current_state_reg ( .D(
        new_AGEMA_signal_4752), .CK(clk), .Q(new_AGEMA_signal_4753), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2477_s_current_state_reg ( .D(
        new_AGEMA_signal_4754), .CK(clk), .Q(new_AGEMA_signal_4755), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2479_s_current_state_reg ( .D(
        new_AGEMA_signal_4756), .CK(clk), .Q(new_AGEMA_signal_4757), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2483_s_current_state_reg ( .D(
        new_AGEMA_signal_4760), .CK(clk), .Q(new_AGEMA_signal_4761), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2487_s_current_state_reg ( .D(
        new_AGEMA_signal_4764), .CK(clk), .Q(new_AGEMA_signal_4765), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2497_s_current_state_reg ( .D(
        new_AGEMA_signal_4774), .CK(clk), .Q(new_AGEMA_signal_4775), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2499_s_current_state_reg ( .D(
        new_AGEMA_signal_4776), .CK(clk), .Q(new_AGEMA_signal_4777), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2501_s_current_state_reg ( .D(
        new_AGEMA_signal_4778), .CK(clk), .Q(new_AGEMA_signal_4779), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2509_s_current_state_reg ( .D(
        new_AGEMA_signal_4786), .CK(clk), .Q(new_AGEMA_signal_4787), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2511_s_current_state_reg ( .D(
        new_AGEMA_signal_4788), .CK(clk), .Q(new_AGEMA_signal_4789), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2513_s_current_state_reg ( .D(
        new_AGEMA_signal_4790), .CK(clk), .Q(new_AGEMA_signal_4791), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2515_s_current_state_reg ( .D(
        new_AGEMA_signal_4792), .CK(clk), .Q(new_AGEMA_signal_4793), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2519_s_current_state_reg ( .D(
        new_AGEMA_signal_4796), .CK(clk), .Q(new_AGEMA_signal_4797), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2523_s_current_state_reg ( .D(
        new_AGEMA_signal_4800), .CK(clk), .Q(new_AGEMA_signal_4801), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2533_s_current_state_reg ( .D(
        new_AGEMA_signal_4810), .CK(clk), .Q(new_AGEMA_signal_4811), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2535_s_current_state_reg ( .D(
        new_AGEMA_signal_4812), .CK(clk), .Q(new_AGEMA_signal_4813), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2537_s_current_state_reg ( .D(
        new_AGEMA_signal_4814), .CK(clk), .Q(new_AGEMA_signal_4815), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2545_s_current_state_reg ( .D(
        new_AGEMA_signal_4822), .CK(clk), .Q(new_AGEMA_signal_4823), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2547_s_current_state_reg ( .D(
        new_AGEMA_signal_4824), .CK(clk), .Q(new_AGEMA_signal_4825), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2549_s_current_state_reg ( .D(
        new_AGEMA_signal_4826), .CK(clk), .Q(new_AGEMA_signal_4827), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2551_s_current_state_reg ( .D(
        new_AGEMA_signal_4828), .CK(clk), .Q(new_AGEMA_signal_4829), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2555_s_current_state_reg ( .D(
        new_AGEMA_signal_4832), .CK(clk), .Q(new_AGEMA_signal_4833), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2559_s_current_state_reg ( .D(
        new_AGEMA_signal_4836), .CK(clk), .Q(new_AGEMA_signal_4837), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2569_s_current_state_reg ( .D(
        new_AGEMA_signal_4846), .CK(clk), .Q(new_AGEMA_signal_4847), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2571_s_current_state_reg ( .D(
        new_AGEMA_signal_4848), .CK(clk), .Q(new_AGEMA_signal_4849), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2573_s_current_state_reg ( .D(
        new_AGEMA_signal_4850), .CK(clk), .Q(new_AGEMA_signal_4851), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2581_s_current_state_reg ( .D(
        new_AGEMA_signal_4858), .CK(clk), .Q(new_AGEMA_signal_4859), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2583_s_current_state_reg ( .D(
        new_AGEMA_signal_4860), .CK(clk), .Q(new_AGEMA_signal_4861), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2585_s_current_state_reg ( .D(
        new_AGEMA_signal_4862), .CK(clk), .Q(new_AGEMA_signal_4863), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2587_s_current_state_reg ( .D(
        new_AGEMA_signal_4864), .CK(clk), .Q(new_AGEMA_signal_4865), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2591_s_current_state_reg ( .D(
        new_AGEMA_signal_4868), .CK(clk), .Q(new_AGEMA_signal_4869), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2595_s_current_state_reg ( .D(
        new_AGEMA_signal_4872), .CK(clk), .Q(new_AGEMA_signal_4873), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2605_s_current_state_reg ( .D(
        new_AGEMA_signal_4882), .CK(clk), .Q(new_AGEMA_signal_4883), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2607_s_current_state_reg ( .D(
        new_AGEMA_signal_4884), .CK(clk), .Q(new_AGEMA_signal_4885), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2609_s_current_state_reg ( .D(
        new_AGEMA_signal_4886), .CK(clk), .Q(new_AGEMA_signal_4887), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2617_s_current_state_reg ( .D(
        new_AGEMA_signal_4894), .CK(clk), .Q(new_AGEMA_signal_4895), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2619_s_current_state_reg ( .D(
        new_AGEMA_signal_4896), .CK(clk), .Q(new_AGEMA_signal_4897), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2621_s_current_state_reg ( .D(
        new_AGEMA_signal_4898), .CK(clk), .Q(new_AGEMA_signal_4899), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2623_s_current_state_reg ( .D(
        new_AGEMA_signal_4900), .CK(clk), .Q(new_AGEMA_signal_4901), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2627_s_current_state_reg ( .D(
        new_AGEMA_signal_4904), .CK(clk), .Q(new_AGEMA_signal_4905), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2631_s_current_state_reg ( .D(
        new_AGEMA_signal_4908), .CK(clk), .Q(new_AGEMA_signal_4909), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2641_s_current_state_reg ( .D(
        new_AGEMA_signal_4918), .CK(clk), .Q(new_AGEMA_signal_4919), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2645_s_current_state_reg ( .D(
        new_AGEMA_signal_4922), .CK(clk), .Q(new_AGEMA_signal_4923), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2649_s_current_state_reg ( .D(
        new_AGEMA_signal_4926), .CK(clk), .Q(new_AGEMA_signal_4927), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2653_s_current_state_reg ( .D(
        new_AGEMA_signal_4930), .CK(clk), .Q(new_AGEMA_signal_4931), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2657_s_current_state_reg ( .D(
        new_AGEMA_signal_4934), .CK(clk), .Q(new_AGEMA_signal_4935), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2661_s_current_state_reg ( .D(
        new_AGEMA_signal_4938), .CK(clk), .Q(new_AGEMA_signal_4939), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2665_s_current_state_reg ( .D(
        new_AGEMA_signal_4942), .CK(clk), .Q(new_AGEMA_signal_4943), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2669_s_current_state_reg ( .D(
        new_AGEMA_signal_4946), .CK(clk), .Q(new_AGEMA_signal_4947), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2673_s_current_state_reg ( .D(
        new_AGEMA_signal_4950), .CK(clk), .Q(new_AGEMA_signal_4951), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2677_s_current_state_reg ( .D(
        new_AGEMA_signal_4954), .CK(clk), .Q(new_AGEMA_signal_4955), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2681_s_current_state_reg ( .D(
        new_AGEMA_signal_4958), .CK(clk), .Q(new_AGEMA_signal_4959), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2685_s_current_state_reg ( .D(
        new_AGEMA_signal_4962), .CK(clk), .Q(new_AGEMA_signal_4963), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2689_s_current_state_reg ( .D(
        new_AGEMA_signal_4966), .CK(clk), .Q(new_AGEMA_signal_4967), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2693_s_current_state_reg ( .D(
        new_AGEMA_signal_4970), .CK(clk), .Q(new_AGEMA_signal_4971), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2697_s_current_state_reg ( .D(
        new_AGEMA_signal_4974), .CK(clk), .Q(new_AGEMA_signal_4975), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2701_s_current_state_reg ( .D(
        new_AGEMA_signal_4978), .CK(clk), .Q(new_AGEMA_signal_4979), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2705_s_current_state_reg ( .D(
        new_AGEMA_signal_4982), .CK(clk), .Q(new_AGEMA_signal_4983), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2709_s_current_state_reg ( .D(
        new_AGEMA_signal_4986), .CK(clk), .Q(new_AGEMA_signal_4987), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2713_s_current_state_reg ( .D(
        new_AGEMA_signal_4990), .CK(clk), .Q(new_AGEMA_signal_4991), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2717_s_current_state_reg ( .D(
        new_AGEMA_signal_4994), .CK(clk), .Q(new_AGEMA_signal_4995), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2721_s_current_state_reg ( .D(
        new_AGEMA_signal_4998), .CK(clk), .Q(new_AGEMA_signal_4999), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2725_s_current_state_reg ( .D(
        new_AGEMA_signal_5002), .CK(clk), .Q(new_AGEMA_signal_5003), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2729_s_current_state_reg ( .D(
        new_AGEMA_signal_5006), .CK(clk), .Q(new_AGEMA_signal_5007), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2733_s_current_state_reg ( .D(
        new_AGEMA_signal_5010), .CK(clk), .Q(new_AGEMA_signal_5011), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2737_s_current_state_reg ( .D(
        new_AGEMA_signal_5014), .CK(clk), .Q(new_AGEMA_signal_5015), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2741_s_current_state_reg ( .D(
        new_AGEMA_signal_5018), .CK(clk), .Q(new_AGEMA_signal_5019), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2745_s_current_state_reg ( .D(
        new_AGEMA_signal_5022), .CK(clk), .Q(new_AGEMA_signal_5023), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2749_s_current_state_reg ( .D(
        new_AGEMA_signal_5026), .CK(clk), .Q(new_AGEMA_signal_5027), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2753_s_current_state_reg ( .D(
        new_AGEMA_signal_5030), .CK(clk), .Q(new_AGEMA_signal_5031), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2757_s_current_state_reg ( .D(
        new_AGEMA_signal_5034), .CK(clk), .Q(new_AGEMA_signal_5035), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2761_s_current_state_reg ( .D(
        new_AGEMA_signal_5038), .CK(clk), .Q(new_AGEMA_signal_5039), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2765_s_current_state_reg ( .D(
        new_AGEMA_signal_5042), .CK(clk), .Q(new_AGEMA_signal_5043), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2769_s_current_state_reg ( .D(
        new_AGEMA_signal_5046), .CK(clk), .Q(new_AGEMA_signal_5047), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2773_s_current_state_reg ( .D(
        new_AGEMA_signal_5050), .CK(clk), .Q(new_AGEMA_signal_5051), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2777_s_current_state_reg ( .D(
        new_AGEMA_signal_5054), .CK(clk), .Q(new_AGEMA_signal_5055), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2781_s_current_state_reg ( .D(
        new_AGEMA_signal_5058), .CK(clk), .Q(new_AGEMA_signal_5059), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2785_s_current_state_reg ( .D(
        new_AGEMA_signal_5062), .CK(clk), .Q(new_AGEMA_signal_5063), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2789_s_current_state_reg ( .D(
        new_AGEMA_signal_5066), .CK(clk), .Q(new_AGEMA_signal_5067), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2793_s_current_state_reg ( .D(
        new_AGEMA_signal_5070), .CK(clk), .Q(new_AGEMA_signal_5071), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2797_s_current_state_reg ( .D(
        new_AGEMA_signal_5074), .CK(clk), .Q(new_AGEMA_signal_5075), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2801_s_current_state_reg ( .D(
        new_AGEMA_signal_5078), .CK(clk), .Q(new_AGEMA_signal_5079), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2805_s_current_state_reg ( .D(
        new_AGEMA_signal_5082), .CK(clk), .Q(new_AGEMA_signal_5083), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2809_s_current_state_reg ( .D(
        new_AGEMA_signal_5086), .CK(clk), .Q(new_AGEMA_signal_5087), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2813_s_current_state_reg ( .D(
        new_AGEMA_signal_5090), .CK(clk), .Q(new_AGEMA_signal_5091), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2817_s_current_state_reg ( .D(
        new_AGEMA_signal_5094), .CK(clk), .Q(new_AGEMA_signal_5095), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2821_s_current_state_reg ( .D(
        new_AGEMA_signal_5098), .CK(clk), .Q(new_AGEMA_signal_5099), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2825_s_current_state_reg ( .D(
        new_AGEMA_signal_5102), .CK(clk), .Q(new_AGEMA_signal_5103), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2829_s_current_state_reg ( .D(
        new_AGEMA_signal_5106), .CK(clk), .Q(new_AGEMA_signal_5107), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2833_s_current_state_reg ( .D(
        new_AGEMA_signal_5110), .CK(clk), .Q(new_AGEMA_signal_5111), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2837_s_current_state_reg ( .D(
        new_AGEMA_signal_5114), .CK(clk), .Q(new_AGEMA_signal_5115), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2841_s_current_state_reg ( .D(
        new_AGEMA_signal_5118), .CK(clk), .Q(new_AGEMA_signal_5119), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2845_s_current_state_reg ( .D(
        new_AGEMA_signal_5122), .CK(clk), .Q(new_AGEMA_signal_5123), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3041_s_current_state_reg ( .D(
        new_AGEMA_signal_5318), .CK(clk), .Q(new_AGEMA_signal_5319), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3045_s_current_state_reg ( .D(
        new_AGEMA_signal_5322), .CK(clk), .Q(new_AGEMA_signal_5323), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3049_s_current_state_reg ( .D(
        new_AGEMA_signal_5326), .CK(clk), .Q(new_AGEMA_signal_5327), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3053_s_current_state_reg ( .D(
        new_AGEMA_signal_5330), .CK(clk), .Q(new_AGEMA_signal_5331), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3057_s_current_state_reg ( .D(
        new_AGEMA_signal_5334), .CK(clk), .Q(new_AGEMA_signal_5335), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3061_s_current_state_reg ( .D(
        new_AGEMA_signal_5338), .CK(clk), .Q(new_AGEMA_signal_5339), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3065_s_current_state_reg ( .D(
        new_AGEMA_signal_5342), .CK(clk), .Q(new_AGEMA_signal_5343), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3069_s_current_state_reg ( .D(
        new_AGEMA_signal_5346), .CK(clk), .Q(new_AGEMA_signal_5347), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3073_s_current_state_reg ( .D(
        new_AGEMA_signal_5350), .CK(clk), .Q(new_AGEMA_signal_5351), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3077_s_current_state_reg ( .D(
        new_AGEMA_signal_5354), .CK(clk), .Q(new_AGEMA_signal_5355), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3081_s_current_state_reg ( .D(
        new_AGEMA_signal_5358), .CK(clk), .Q(new_AGEMA_signal_5359), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3085_s_current_state_reg ( .D(
        new_AGEMA_signal_5362), .CK(clk), .Q(new_AGEMA_signal_5363), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3089_s_current_state_reg ( .D(
        new_AGEMA_signal_5366), .CK(clk), .Q(new_AGEMA_signal_5367), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3093_s_current_state_reg ( .D(
        new_AGEMA_signal_5370), .CK(clk), .Q(new_AGEMA_signal_5371), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3097_s_current_state_reg ( .D(
        new_AGEMA_signal_5374), .CK(clk), .Q(new_AGEMA_signal_5375), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3101_s_current_state_reg ( .D(
        new_AGEMA_signal_5378), .CK(clk), .Q(new_AGEMA_signal_5379), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3105_s_current_state_reg ( .D(
        new_AGEMA_signal_5382), .CK(clk), .Q(new_AGEMA_signal_5383), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3109_s_current_state_reg ( .D(
        new_AGEMA_signal_5386), .CK(clk), .Q(new_AGEMA_signal_5387), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3113_s_current_state_reg ( .D(
        new_AGEMA_signal_5390), .CK(clk), .Q(new_AGEMA_signal_5391), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3117_s_current_state_reg ( .D(
        new_AGEMA_signal_5394), .CK(clk), .Q(new_AGEMA_signal_5395), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3121_s_current_state_reg ( .D(
        new_AGEMA_signal_5398), .CK(clk), .Q(new_AGEMA_signal_5399), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3125_s_current_state_reg ( .D(
        new_AGEMA_signal_5402), .CK(clk), .Q(new_AGEMA_signal_5403), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3129_s_current_state_reg ( .D(
        new_AGEMA_signal_5406), .CK(clk), .Q(new_AGEMA_signal_5407), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3133_s_current_state_reg ( .D(
        new_AGEMA_signal_5410), .CK(clk), .Q(new_AGEMA_signal_5411), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3137_s_current_state_reg ( .D(
        new_AGEMA_signal_5414), .CK(clk), .Q(new_AGEMA_signal_5415), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3141_s_current_state_reg ( .D(
        new_AGEMA_signal_5418), .CK(clk), .Q(new_AGEMA_signal_5419), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3145_s_current_state_reg ( .D(
        new_AGEMA_signal_5422), .CK(clk), .Q(new_AGEMA_signal_5423), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3149_s_current_state_reg ( .D(
        new_AGEMA_signal_5426), .CK(clk), .Q(new_AGEMA_signal_5427), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3153_s_current_state_reg ( .D(
        new_AGEMA_signal_5430), .CK(clk), .Q(new_AGEMA_signal_5431), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3157_s_current_state_reg ( .D(
        new_AGEMA_signal_5434), .CK(clk), .Q(new_AGEMA_signal_5435), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3161_s_current_state_reg ( .D(
        new_AGEMA_signal_5438), .CK(clk), .Q(new_AGEMA_signal_5439), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3165_s_current_state_reg ( .D(
        new_AGEMA_signal_5442), .CK(clk), .Q(new_AGEMA_signal_5443), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3169_s_current_state_reg ( .D(
        new_AGEMA_signal_5446), .CK(clk), .Q(new_AGEMA_signal_5447), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3173_s_current_state_reg ( .D(
        new_AGEMA_signal_5450), .CK(clk), .Q(new_AGEMA_signal_5451), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3177_s_current_state_reg ( .D(
        new_AGEMA_signal_5454), .CK(clk), .Q(new_AGEMA_signal_5455), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3181_s_current_state_reg ( .D(
        new_AGEMA_signal_5458), .CK(clk), .Q(new_AGEMA_signal_5459), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3185_s_current_state_reg ( .D(
        new_AGEMA_signal_5462), .CK(clk), .Q(new_AGEMA_signal_5463), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3189_s_current_state_reg ( .D(
        new_AGEMA_signal_5466), .CK(clk), .Q(new_AGEMA_signal_5467), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3193_s_current_state_reg ( .D(
        new_AGEMA_signal_5470), .CK(clk), .Q(new_AGEMA_signal_5471), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3197_s_current_state_reg ( .D(
        new_AGEMA_signal_5474), .CK(clk), .Q(new_AGEMA_signal_5475), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3201_s_current_state_reg ( .D(
        new_AGEMA_signal_5478), .CK(clk), .Q(new_AGEMA_signal_5479), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3205_s_current_state_reg ( .D(
        new_AGEMA_signal_5482), .CK(clk), .Q(new_AGEMA_signal_5483), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3209_s_current_state_reg ( .D(
        new_AGEMA_signal_5486), .CK(clk), .Q(new_AGEMA_signal_5487), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3213_s_current_state_reg ( .D(
        new_AGEMA_signal_5490), .CK(clk), .Q(new_AGEMA_signal_5491), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3217_s_current_state_reg ( .D(
        new_AGEMA_signal_5494), .CK(clk), .Q(new_AGEMA_signal_5495), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3221_s_current_state_reg ( .D(
        new_AGEMA_signal_5498), .CK(clk), .Q(new_AGEMA_signal_5499), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3225_s_current_state_reg ( .D(
        new_AGEMA_signal_5502), .CK(clk), .Q(new_AGEMA_signal_5503), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3229_s_current_state_reg ( .D(
        new_AGEMA_signal_5506), .CK(clk), .Q(new_AGEMA_signal_5507), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3233_s_current_state_reg ( .D(
        new_AGEMA_signal_5510), .CK(clk), .Q(new_AGEMA_signal_5511), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3237_s_current_state_reg ( .D(
        new_AGEMA_signal_5514), .CK(clk), .Q(new_AGEMA_signal_5515), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3241_s_current_state_reg ( .D(
        new_AGEMA_signal_5518), .CK(clk), .Q(new_AGEMA_signal_5519), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3245_s_current_state_reg ( .D(
        new_AGEMA_signal_5522), .CK(clk), .Q(new_AGEMA_signal_5523), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3249_s_current_state_reg ( .D(
        new_AGEMA_signal_5526), .CK(clk), .Q(new_AGEMA_signal_5527), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3253_s_current_state_reg ( .D(
        new_AGEMA_signal_5530), .CK(clk), .Q(new_AGEMA_signal_5531), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3257_s_current_state_reg ( .D(
        new_AGEMA_signal_5534), .CK(clk), .Q(new_AGEMA_signal_5535), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3261_s_current_state_reg ( .D(
        new_AGEMA_signal_5538), .CK(clk), .Q(new_AGEMA_signal_5539), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3265_s_current_state_reg ( .D(
        new_AGEMA_signal_5542), .CK(clk), .Q(new_AGEMA_signal_5543), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3269_s_current_state_reg ( .D(
        new_AGEMA_signal_5546), .CK(clk), .Q(new_AGEMA_signal_5547), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3273_s_current_state_reg ( .D(
        new_AGEMA_signal_5550), .CK(clk), .Q(new_AGEMA_signal_5551), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3277_s_current_state_reg ( .D(
        new_AGEMA_signal_5554), .CK(clk), .Q(new_AGEMA_signal_5555), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3281_s_current_state_reg ( .D(
        new_AGEMA_signal_5558), .CK(clk), .Q(new_AGEMA_signal_5559), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3285_s_current_state_reg ( .D(
        new_AGEMA_signal_5562), .CK(clk), .Q(new_AGEMA_signal_5563), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3289_s_current_state_reg ( .D(
        new_AGEMA_signal_5566), .CK(clk), .Q(new_AGEMA_signal_5567), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3293_s_current_state_reg ( .D(
        new_AGEMA_signal_5570), .CK(clk), .Q(new_AGEMA_signal_5571), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3297_s_current_state_reg ( .D(
        new_AGEMA_signal_5574), .CK(clk), .Q(new_AGEMA_signal_5575), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3301_s_current_state_reg ( .D(
        new_AGEMA_signal_5578), .CK(clk), .Q(new_AGEMA_signal_5579), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3305_s_current_state_reg ( .D(
        new_AGEMA_signal_5582), .CK(clk), .Q(new_AGEMA_signal_5583), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3309_s_current_state_reg ( .D(
        new_AGEMA_signal_5586), .CK(clk), .Q(new_AGEMA_signal_5587), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3313_s_current_state_reg ( .D(
        new_AGEMA_signal_5590), .CK(clk), .Q(new_AGEMA_signal_5591), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3317_s_current_state_reg ( .D(
        new_AGEMA_signal_5594), .CK(clk), .Q(new_AGEMA_signal_5595), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3321_s_current_state_reg ( .D(
        new_AGEMA_signal_5598), .CK(clk), .Q(new_AGEMA_signal_5599), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3325_s_current_state_reg ( .D(
        new_AGEMA_signal_5602), .CK(clk), .Q(new_AGEMA_signal_5603), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3329_s_current_state_reg ( .D(
        new_AGEMA_signal_5606), .CK(clk), .Q(new_AGEMA_signal_5607), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3333_s_current_state_reg ( .D(
        new_AGEMA_signal_5610), .CK(clk), .Q(new_AGEMA_signal_5611), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3337_s_current_state_reg ( .D(
        new_AGEMA_signal_5614), .CK(clk), .Q(new_AGEMA_signal_5615), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3341_s_current_state_reg ( .D(
        new_AGEMA_signal_5618), .CK(clk), .Q(new_AGEMA_signal_5619), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3345_s_current_state_reg ( .D(
        new_AGEMA_signal_5622), .CK(clk), .Q(new_AGEMA_signal_5623), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3349_s_current_state_reg ( .D(
        new_AGEMA_signal_5626), .CK(clk), .Q(new_AGEMA_signal_5627), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3353_s_current_state_reg ( .D(
        new_AGEMA_signal_5630), .CK(clk), .Q(new_AGEMA_signal_5631), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3357_s_current_state_reg ( .D(
        new_AGEMA_signal_5634), .CK(clk), .Q(new_AGEMA_signal_5635), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3361_s_current_state_reg ( .D(
        new_AGEMA_signal_5638), .CK(clk), .Q(new_AGEMA_signal_5639), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3365_s_current_state_reg ( .D(
        new_AGEMA_signal_5642), .CK(clk), .Q(new_AGEMA_signal_5643), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3369_s_current_state_reg ( .D(
        new_AGEMA_signal_5646), .CK(clk), .Q(new_AGEMA_signal_5647), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3373_s_current_state_reg ( .D(
        new_AGEMA_signal_5650), .CK(clk), .Q(new_AGEMA_signal_5651), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3377_s_current_state_reg ( .D(
        new_AGEMA_signal_5654), .CK(clk), .Q(new_AGEMA_signal_5655), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3381_s_current_state_reg ( .D(
        new_AGEMA_signal_5658), .CK(clk), .Q(new_AGEMA_signal_5659), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3385_s_current_state_reg ( .D(
        new_AGEMA_signal_5662), .CK(clk), .Q(new_AGEMA_signal_5663), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3389_s_current_state_reg ( .D(
        new_AGEMA_signal_5666), .CK(clk), .Q(new_AGEMA_signal_5667), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3393_s_current_state_reg ( .D(
        new_AGEMA_signal_5670), .CK(clk), .Q(new_AGEMA_signal_5671), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3397_s_current_state_reg ( .D(
        new_AGEMA_signal_5674), .CK(clk), .Q(new_AGEMA_signal_5675), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3401_s_current_state_reg ( .D(
        new_AGEMA_signal_5678), .CK(clk), .Q(new_AGEMA_signal_5679), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3405_s_current_state_reg ( .D(
        new_AGEMA_signal_5682), .CK(clk), .Q(new_AGEMA_signal_5683), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3409_s_current_state_reg ( .D(
        new_AGEMA_signal_5686), .CK(clk), .Q(new_AGEMA_signal_5687), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3413_s_current_state_reg ( .D(
        new_AGEMA_signal_5690), .CK(clk), .Q(new_AGEMA_signal_5691), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3417_s_current_state_reg ( .D(
        new_AGEMA_signal_5694), .CK(clk), .Q(new_AGEMA_signal_5695), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3421_s_current_state_reg ( .D(
        new_AGEMA_signal_5698), .CK(clk), .Q(new_AGEMA_signal_5699), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3425_s_current_state_reg ( .D(
        new_AGEMA_signal_5702), .CK(clk), .Q(new_AGEMA_signal_5703), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3429_s_current_state_reg ( .D(
        new_AGEMA_signal_5706), .CK(clk), .Q(new_AGEMA_signal_5707), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3433_s_current_state_reg ( .D(
        new_AGEMA_signal_5710), .CK(clk), .Q(new_AGEMA_signal_5711), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3437_s_current_state_reg ( .D(
        new_AGEMA_signal_5714), .CK(clk), .Q(new_AGEMA_signal_5715), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3441_s_current_state_reg ( .D(
        new_AGEMA_signal_5718), .CK(clk), .Q(new_AGEMA_signal_5719), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3445_s_current_state_reg ( .D(
        new_AGEMA_signal_5722), .CK(clk), .Q(new_AGEMA_signal_5723), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3449_s_current_state_reg ( .D(
        new_AGEMA_signal_5726), .CK(clk), .Q(new_AGEMA_signal_5727), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3453_s_current_state_reg ( .D(
        new_AGEMA_signal_5730), .CK(clk), .Q(new_AGEMA_signal_5731), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3457_s_current_state_reg ( .D(
        new_AGEMA_signal_5734), .CK(clk), .Q(new_AGEMA_signal_5735), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3461_s_current_state_reg ( .D(
        new_AGEMA_signal_5738), .CK(clk), .Q(new_AGEMA_signal_5739), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3465_s_current_state_reg ( .D(
        new_AGEMA_signal_5742), .CK(clk), .Q(new_AGEMA_signal_5743), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3469_s_current_state_reg ( .D(
        new_AGEMA_signal_5746), .CK(clk), .Q(new_AGEMA_signal_5747), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3473_s_current_state_reg ( .D(
        new_AGEMA_signal_5750), .CK(clk), .Q(new_AGEMA_signal_5751), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3477_s_current_state_reg ( .D(
        new_AGEMA_signal_5754), .CK(clk), .Q(new_AGEMA_signal_5755), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3481_s_current_state_reg ( .D(
        new_AGEMA_signal_5758), .CK(clk), .Q(new_AGEMA_signal_5759), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3485_s_current_state_reg ( .D(
        new_AGEMA_signal_5762), .CK(clk), .Q(new_AGEMA_signal_5763), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3489_s_current_state_reg ( .D(
        new_AGEMA_signal_5766), .CK(clk), .Q(new_AGEMA_signal_5767), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3493_s_current_state_reg ( .D(
        new_AGEMA_signal_5770), .CK(clk), .Q(new_AGEMA_signal_5771), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3497_s_current_state_reg ( .D(
        new_AGEMA_signal_5774), .CK(clk), .Q(new_AGEMA_signal_5775), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3501_s_current_state_reg ( .D(
        new_AGEMA_signal_5778), .CK(clk), .Q(new_AGEMA_signal_5779), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3505_s_current_state_reg ( .D(
        new_AGEMA_signal_5782), .CK(clk), .Q(new_AGEMA_signal_5783), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3509_s_current_state_reg ( .D(
        new_AGEMA_signal_5786), .CK(clk), .Q(new_AGEMA_signal_5787), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3513_s_current_state_reg ( .D(
        new_AGEMA_signal_5790), .CK(clk), .Q(new_AGEMA_signal_5791), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3517_s_current_state_reg ( .D(
        new_AGEMA_signal_5794), .CK(clk), .Q(new_AGEMA_signal_5795), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3521_s_current_state_reg ( .D(
        new_AGEMA_signal_5798), .CK(clk), .Q(new_AGEMA_signal_5799), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3525_s_current_state_reg ( .D(
        new_AGEMA_signal_5802), .CK(clk), .Q(new_AGEMA_signal_5803), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3529_s_current_state_reg ( .D(
        new_AGEMA_signal_5806), .CK(clk), .Q(new_AGEMA_signal_5807), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3533_s_current_state_reg ( .D(
        new_AGEMA_signal_5810), .CK(clk), .Q(new_AGEMA_signal_5811), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3537_s_current_state_reg ( .D(
        new_AGEMA_signal_5814), .CK(clk), .Q(new_AGEMA_signal_5815), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3541_s_current_state_reg ( .D(
        new_AGEMA_signal_5818), .CK(clk), .Q(new_AGEMA_signal_5819), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3545_s_current_state_reg ( .D(
        new_AGEMA_signal_5822), .CK(clk), .Q(new_AGEMA_signal_5823), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3549_s_current_state_reg ( .D(
        new_AGEMA_signal_5826), .CK(clk), .Q(new_AGEMA_signal_5827), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3553_s_current_state_reg ( .D(
        new_AGEMA_signal_5830), .CK(clk), .Q(new_AGEMA_signal_5831), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3557_s_current_state_reg ( .D(
        new_AGEMA_signal_5834), .CK(clk), .Q(new_AGEMA_signal_5835), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3561_s_current_state_reg ( .D(
        new_AGEMA_signal_5838), .CK(clk), .Q(new_AGEMA_signal_5839), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3565_s_current_state_reg ( .D(
        new_AGEMA_signal_5842), .CK(clk), .Q(new_AGEMA_signal_5843), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3569_s_current_state_reg ( .D(
        new_AGEMA_signal_5846), .CK(clk), .Q(new_AGEMA_signal_5847), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3573_s_current_state_reg ( .D(
        new_AGEMA_signal_5850), .CK(clk), .Q(new_AGEMA_signal_5851), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3577_s_current_state_reg ( .D(
        new_AGEMA_signal_5854), .CK(clk), .Q(new_AGEMA_signal_5855), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3581_s_current_state_reg ( .D(
        new_AGEMA_signal_5858), .CK(clk), .Q(new_AGEMA_signal_5859), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3585_s_current_state_reg ( .D(
        new_AGEMA_signal_5862), .CK(clk), .Q(new_AGEMA_signal_5863), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3589_s_current_state_reg ( .D(
        new_AGEMA_signal_5866), .CK(clk), .Q(new_AGEMA_signal_5867), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3593_s_current_state_reg ( .D(
        new_AGEMA_signal_5870), .CK(clk), .Q(new_AGEMA_signal_5871), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3597_s_current_state_reg ( .D(
        new_AGEMA_signal_5874), .CK(clk), .Q(new_AGEMA_signal_5875), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3601_s_current_state_reg ( .D(
        new_AGEMA_signal_5878), .CK(clk), .Q(new_AGEMA_signal_5879), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3605_s_current_state_reg ( .D(
        new_AGEMA_signal_5882), .CK(clk), .Q(new_AGEMA_signal_5883), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3609_s_current_state_reg ( .D(
        new_AGEMA_signal_5886), .CK(clk), .Q(new_AGEMA_signal_5887), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3613_s_current_state_reg ( .D(
        new_AGEMA_signal_5890), .CK(clk), .Q(new_AGEMA_signal_5891), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3617_s_current_state_reg ( .D(
        new_AGEMA_signal_5894), .CK(clk), .Q(new_AGEMA_signal_5895), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3621_s_current_state_reg ( .D(
        new_AGEMA_signal_5898), .CK(clk), .Q(new_AGEMA_signal_5899), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3625_s_current_state_reg ( .D(
        new_AGEMA_signal_5902), .CK(clk), .Q(new_AGEMA_signal_5903), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3629_s_current_state_reg ( .D(
        new_AGEMA_signal_5906), .CK(clk), .Q(new_AGEMA_signal_5907), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3633_s_current_state_reg ( .D(
        new_AGEMA_signal_5910), .CK(clk), .Q(new_AGEMA_signal_5911), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3637_s_current_state_reg ( .D(
        new_AGEMA_signal_5914), .CK(clk), .Q(new_AGEMA_signal_5915), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3641_s_current_state_reg ( .D(
        new_AGEMA_signal_5918), .CK(clk), .Q(new_AGEMA_signal_5919), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3645_s_current_state_reg ( .D(
        new_AGEMA_signal_5922), .CK(clk), .Q(new_AGEMA_signal_5923), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3649_s_current_state_reg ( .D(
        new_AGEMA_signal_5926), .CK(clk), .Q(new_AGEMA_signal_5927), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3653_s_current_state_reg ( .D(
        new_AGEMA_signal_5930), .CK(clk), .Q(new_AGEMA_signal_5931), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3657_s_current_state_reg ( .D(
        new_AGEMA_signal_5934), .CK(clk), .Q(new_AGEMA_signal_5935), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3661_s_current_state_reg ( .D(
        new_AGEMA_signal_5938), .CK(clk), .Q(new_AGEMA_signal_5939), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3665_s_current_state_reg ( .D(
        new_AGEMA_signal_5942), .CK(clk), .Q(new_AGEMA_signal_5943), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3669_s_current_state_reg ( .D(
        new_AGEMA_signal_5946), .CK(clk), .Q(new_AGEMA_signal_5947), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3673_s_current_state_reg ( .D(
        new_AGEMA_signal_5950), .CK(clk), .Q(new_AGEMA_signal_5951), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3677_s_current_state_reg ( .D(
        new_AGEMA_signal_5954), .CK(clk), .Q(new_AGEMA_signal_5955), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3681_s_current_state_reg ( .D(
        new_AGEMA_signal_5958), .CK(clk), .Q(new_AGEMA_signal_5959), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3685_s_current_state_reg ( .D(
        new_AGEMA_signal_5962), .CK(clk), .Q(new_AGEMA_signal_5963), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3689_s_current_state_reg ( .D(
        new_AGEMA_signal_5966), .CK(clk), .Q(new_AGEMA_signal_5967), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3693_s_current_state_reg ( .D(
        new_AGEMA_signal_5970), .CK(clk), .Q(new_AGEMA_signal_5971), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3697_s_current_state_reg ( .D(
        new_AGEMA_signal_5974), .CK(clk), .Q(new_AGEMA_signal_5975), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3701_s_current_state_reg ( .D(
        new_AGEMA_signal_5978), .CK(clk), .Q(new_AGEMA_signal_5979), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3705_s_current_state_reg ( .D(
        new_AGEMA_signal_5982), .CK(clk), .Q(new_AGEMA_signal_5983), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3709_s_current_state_reg ( .D(
        new_AGEMA_signal_5986), .CK(clk), .Q(new_AGEMA_signal_5987), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3713_s_current_state_reg ( .D(
        new_AGEMA_signal_5990), .CK(clk), .Q(new_AGEMA_signal_5991), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3717_s_current_state_reg ( .D(
        new_AGEMA_signal_5994), .CK(clk), .Q(new_AGEMA_signal_5995), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3721_s_current_state_reg ( .D(
        new_AGEMA_signal_5998), .CK(clk), .Q(new_AGEMA_signal_5999), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3725_s_current_state_reg ( .D(
        new_AGEMA_signal_6002), .CK(clk), .Q(new_AGEMA_signal_6003), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3729_s_current_state_reg ( .D(
        new_AGEMA_signal_6006), .CK(clk), .Q(new_AGEMA_signal_6007), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3733_s_current_state_reg ( .D(
        new_AGEMA_signal_6010), .CK(clk), .Q(new_AGEMA_signal_6011), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3737_s_current_state_reg ( .D(
        new_AGEMA_signal_6014), .CK(clk), .Q(new_AGEMA_signal_6015), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3741_s_current_state_reg ( .D(
        new_AGEMA_signal_6018), .CK(clk), .Q(new_AGEMA_signal_6019), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3745_s_current_state_reg ( .D(
        new_AGEMA_signal_6022), .CK(clk), .Q(new_AGEMA_signal_6023), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3749_s_current_state_reg ( .D(
        new_AGEMA_signal_6026), .CK(clk), .Q(new_AGEMA_signal_6027), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3753_s_current_state_reg ( .D(
        new_AGEMA_signal_6030), .CK(clk), .Q(new_AGEMA_signal_6031), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3757_s_current_state_reg ( .D(
        new_AGEMA_signal_6034), .CK(clk), .Q(new_AGEMA_signal_6035), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3761_s_current_state_reg ( .D(
        new_AGEMA_signal_6038), .CK(clk), .Q(new_AGEMA_signal_6039), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3765_s_current_state_reg ( .D(
        new_AGEMA_signal_6042), .CK(clk), .Q(new_AGEMA_signal_6043), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3769_s_current_state_reg ( .D(
        new_AGEMA_signal_6046), .CK(clk), .Q(new_AGEMA_signal_6047), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3773_s_current_state_reg ( .D(
        new_AGEMA_signal_6050), .CK(clk), .Q(new_AGEMA_signal_6051), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3777_s_current_state_reg ( .D(
        new_AGEMA_signal_6054), .CK(clk), .Q(new_AGEMA_signal_6055), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3781_s_current_state_reg ( .D(
        new_AGEMA_signal_6058), .CK(clk), .Q(new_AGEMA_signal_6059), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3785_s_current_state_reg ( .D(
        new_AGEMA_signal_6062), .CK(clk), .Q(new_AGEMA_signal_6063), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3789_s_current_state_reg ( .D(
        new_AGEMA_signal_6066), .CK(clk), .Q(new_AGEMA_signal_6067), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3793_s_current_state_reg ( .D(
        new_AGEMA_signal_6070), .CK(clk), .Q(new_AGEMA_signal_6071), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3797_s_current_state_reg ( .D(
        new_AGEMA_signal_6074), .CK(clk), .Q(new_AGEMA_signal_6075), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3801_s_current_state_reg ( .D(
        new_AGEMA_signal_6078), .CK(clk), .Q(new_AGEMA_signal_6079), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3805_s_current_state_reg ( .D(
        new_AGEMA_signal_6082), .CK(clk), .Q(new_AGEMA_signal_6083), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3809_s_current_state_reg ( .D(
        new_AGEMA_signal_6086), .CK(clk), .Q(new_AGEMA_signal_6087), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3813_s_current_state_reg ( .D(
        new_AGEMA_signal_6090), .CK(clk), .Q(new_AGEMA_signal_6091), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3817_s_current_state_reg ( .D(
        new_AGEMA_signal_6094), .CK(clk), .Q(new_AGEMA_signal_6095), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3821_s_current_state_reg ( .D(
        new_AGEMA_signal_6098), .CK(clk), .Q(new_AGEMA_signal_6099), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3825_s_current_state_reg ( .D(
        new_AGEMA_signal_6102), .CK(clk), .Q(new_AGEMA_signal_6103), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3829_s_current_state_reg ( .D(
        new_AGEMA_signal_6106), .CK(clk), .Q(new_AGEMA_signal_6107), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1678_s_current_state_reg ( .D(n45), .CK(clk), 
        .Q(new_AGEMA_signal_3956), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1682_s_current_state_reg ( .D(
        new_AGEMA_signal_3959), .CK(clk), .Q(new_AGEMA_signal_3960), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1686_s_current_state_reg ( .D(
        new_AGEMA_signal_3963), .CK(clk), .Q(new_AGEMA_signal_3964), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1690_s_current_state_reg ( .D(
        new_AGEMA_signal_3967), .CK(clk), .Q(new_AGEMA_signal_3968), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1694_s_current_state_reg ( .D(
        new_AGEMA_signal_3971), .CK(clk), .Q(new_AGEMA_signal_3972), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1698_s_current_state_reg ( .D(
        new_AGEMA_signal_3975), .CK(clk), .Q(new_AGEMA_signal_3976), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1702_s_current_state_reg ( .D(
        new_AGEMA_signal_3979), .CK(clk), .Q(new_AGEMA_signal_3980), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1706_s_current_state_reg ( .D(
        new_AGEMA_signal_3983), .CK(clk), .Q(new_AGEMA_signal_3984), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1710_s_current_state_reg ( .D(
        new_AGEMA_signal_3987), .CK(clk), .Q(new_AGEMA_signal_3988), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1714_s_current_state_reg ( .D(
        new_AGEMA_signal_3991), .CK(clk), .Q(new_AGEMA_signal_3992), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1718_s_current_state_reg ( .D(
        new_AGEMA_signal_3995), .CK(clk), .Q(new_AGEMA_signal_3996), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1722_s_current_state_reg ( .D(
        new_AGEMA_signal_3999), .CK(clk), .Q(new_AGEMA_signal_4000), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1726_s_current_state_reg ( .D(
        new_AGEMA_signal_4003), .CK(clk), .Q(new_AGEMA_signal_4004), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1730_s_current_state_reg ( .D(
        new_AGEMA_signal_4007), .CK(clk), .Q(new_AGEMA_signal_4008), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1734_s_current_state_reg ( .D(
        new_AGEMA_signal_4011), .CK(clk), .Q(new_AGEMA_signal_4012), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1738_s_current_state_reg ( .D(
        new_AGEMA_signal_4015), .CK(clk), .Q(new_AGEMA_signal_4016), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1742_s_current_state_reg ( .D(
        new_AGEMA_signal_4019), .CK(clk), .Q(new_AGEMA_signal_4020), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1746_s_current_state_reg ( .D(
        new_AGEMA_signal_4023), .CK(clk), .Q(new_AGEMA_signal_4024), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1750_s_current_state_reg ( .D(
        new_AGEMA_signal_4027), .CK(clk), .Q(new_AGEMA_signal_4028), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1754_s_current_state_reg ( .D(
        new_AGEMA_signal_4031), .CK(clk), .Q(new_AGEMA_signal_4032), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1758_s_current_state_reg ( .D(
        new_AGEMA_signal_4035), .CK(clk), .Q(new_AGEMA_signal_4036), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1762_s_current_state_reg ( .D(
        new_AGEMA_signal_4039), .CK(clk), .Q(new_AGEMA_signal_4040), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1766_s_current_state_reg ( .D(
        new_AGEMA_signal_4043), .CK(clk), .Q(new_AGEMA_signal_4044), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1770_s_current_state_reg ( .D(
        new_AGEMA_signal_4047), .CK(clk), .Q(new_AGEMA_signal_4048), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1774_s_current_state_reg ( .D(
        new_AGEMA_signal_4051), .CK(clk), .Q(new_AGEMA_signal_4052), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1778_s_current_state_reg ( .D(
        new_AGEMA_signal_4055), .CK(clk), .Q(new_AGEMA_signal_4056), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1782_s_current_state_reg ( .D(
        new_AGEMA_signal_4059), .CK(clk), .Q(new_AGEMA_signal_4060), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1786_s_current_state_reg ( .D(
        new_AGEMA_signal_4063), .CK(clk), .Q(new_AGEMA_signal_4064), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1790_s_current_state_reg ( .D(
        new_AGEMA_signal_4067), .CK(clk), .Q(new_AGEMA_signal_4068), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1794_s_current_state_reg ( .D(
        new_AGEMA_signal_4071), .CK(clk), .Q(new_AGEMA_signal_4072), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1798_s_current_state_reg ( .D(
        new_AGEMA_signal_4075), .CK(clk), .Q(new_AGEMA_signal_4076), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1802_s_current_state_reg ( .D(
        new_AGEMA_signal_4079), .CK(clk), .Q(new_AGEMA_signal_4080), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1806_s_current_state_reg ( .D(
        new_AGEMA_signal_4083), .CK(clk), .Q(new_AGEMA_signal_4084), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1810_s_current_state_reg ( .D(
        new_AGEMA_signal_4087), .CK(clk), .Q(new_AGEMA_signal_4088), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1814_s_current_state_reg ( .D(
        new_AGEMA_signal_4091), .CK(clk), .Q(new_AGEMA_signal_4092), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1818_s_current_state_reg ( .D(
        new_AGEMA_signal_4095), .CK(clk), .Q(new_AGEMA_signal_4096), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1822_s_current_state_reg ( .D(
        new_AGEMA_signal_4099), .CK(clk), .Q(new_AGEMA_signal_4100), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1826_s_current_state_reg ( .D(
        new_AGEMA_signal_4103), .CK(clk), .Q(new_AGEMA_signal_4104), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1830_s_current_state_reg ( .D(
        new_AGEMA_signal_4107), .CK(clk), .Q(new_AGEMA_signal_4108), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1834_s_current_state_reg ( .D(
        new_AGEMA_signal_4111), .CK(clk), .Q(new_AGEMA_signal_4112), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1838_s_current_state_reg ( .D(
        new_AGEMA_signal_4115), .CK(clk), .Q(new_AGEMA_signal_4116), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1842_s_current_state_reg ( .D(
        new_AGEMA_signal_4119), .CK(clk), .Q(new_AGEMA_signal_4120), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1846_s_current_state_reg ( .D(
        new_AGEMA_signal_4123), .CK(clk), .Q(new_AGEMA_signal_4124), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1850_s_current_state_reg ( .D(
        new_AGEMA_signal_4127), .CK(clk), .Q(new_AGEMA_signal_4128), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1854_s_current_state_reg ( .D(
        new_AGEMA_signal_4131), .CK(clk), .Q(new_AGEMA_signal_4132), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1858_s_current_state_reg ( .D(
        new_AGEMA_signal_4135), .CK(clk), .Q(new_AGEMA_signal_4136), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1862_s_current_state_reg ( .D(
        new_AGEMA_signal_4139), .CK(clk), .Q(new_AGEMA_signal_4140), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1866_s_current_state_reg ( .D(
        new_AGEMA_signal_4143), .CK(clk), .Q(new_AGEMA_signal_4144), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1870_s_current_state_reg ( .D(
        new_AGEMA_signal_4147), .CK(clk), .Q(new_AGEMA_signal_4148), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1874_s_current_state_reg ( .D(
        new_AGEMA_signal_4151), .CK(clk), .Q(new_AGEMA_signal_4152), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1878_s_current_state_reg ( .D(
        new_AGEMA_signal_4155), .CK(clk), .Q(new_AGEMA_signal_4156), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1882_s_current_state_reg ( .D(
        new_AGEMA_signal_4159), .CK(clk), .Q(new_AGEMA_signal_4160), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1886_s_current_state_reg ( .D(
        new_AGEMA_signal_4163), .CK(clk), .Q(new_AGEMA_signal_4164), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1890_s_current_state_reg ( .D(
        new_AGEMA_signal_4167), .CK(clk), .Q(new_AGEMA_signal_4168), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1894_s_current_state_reg ( .D(
        new_AGEMA_signal_4171), .CK(clk), .Q(new_AGEMA_signal_4172), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1898_s_current_state_reg ( .D(
        new_AGEMA_signal_4175), .CK(clk), .Q(new_AGEMA_signal_4176), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1902_s_current_state_reg ( .D(
        new_AGEMA_signal_4179), .CK(clk), .Q(new_AGEMA_signal_4180), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1906_s_current_state_reg ( .D(
        new_AGEMA_signal_4183), .CK(clk), .Q(new_AGEMA_signal_4184), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1910_s_current_state_reg ( .D(
        new_AGEMA_signal_4187), .CK(clk), .Q(new_AGEMA_signal_4188), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1914_s_current_state_reg ( .D(
        new_AGEMA_signal_4191), .CK(clk), .Q(new_AGEMA_signal_4192), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1918_s_current_state_reg ( .D(
        new_AGEMA_signal_4195), .CK(clk), .Q(new_AGEMA_signal_4196), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1922_s_current_state_reg ( .D(
        new_AGEMA_signal_4199), .CK(clk), .Q(new_AGEMA_signal_4200), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1926_s_current_state_reg ( .D(
        new_AGEMA_signal_4203), .CK(clk), .Q(new_AGEMA_signal_4204), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1930_s_current_state_reg ( .D(
        new_AGEMA_signal_4207), .CK(clk), .Q(new_AGEMA_signal_4208), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1934_s_current_state_reg ( .D(
        new_AGEMA_signal_4211), .CK(clk), .Q(new_AGEMA_signal_4212), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1938_s_current_state_reg ( .D(
        new_AGEMA_signal_4215), .CK(clk), .Q(new_AGEMA_signal_4216), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1942_s_current_state_reg ( .D(
        new_AGEMA_signal_4219), .CK(clk), .Q(new_AGEMA_signal_4220), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1946_s_current_state_reg ( .D(
        new_AGEMA_signal_4223), .CK(clk), .Q(new_AGEMA_signal_4224), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1950_s_current_state_reg ( .D(
        new_AGEMA_signal_4227), .CK(clk), .Q(new_AGEMA_signal_4228), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1954_s_current_state_reg ( .D(
        new_AGEMA_signal_4231), .CK(clk), .Q(new_AGEMA_signal_4232), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1958_s_current_state_reg ( .D(
        new_AGEMA_signal_4235), .CK(clk), .Q(new_AGEMA_signal_4236), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1962_s_current_state_reg ( .D(
        new_AGEMA_signal_4239), .CK(clk), .Q(new_AGEMA_signal_4240), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1966_s_current_state_reg ( .D(
        new_AGEMA_signal_4243), .CK(clk), .Q(new_AGEMA_signal_4244), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1970_s_current_state_reg ( .D(
        new_AGEMA_signal_4247), .CK(clk), .Q(new_AGEMA_signal_4248), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1974_s_current_state_reg ( .D(
        new_AGEMA_signal_4251), .CK(clk), .Q(new_AGEMA_signal_4252), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1978_s_current_state_reg ( .D(
        new_AGEMA_signal_4255), .CK(clk), .Q(new_AGEMA_signal_4256), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1982_s_current_state_reg ( .D(
        new_AGEMA_signal_4259), .CK(clk), .Q(new_AGEMA_signal_4260), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1986_s_current_state_reg ( .D(
        new_AGEMA_signal_4263), .CK(clk), .Q(new_AGEMA_signal_4264), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1990_s_current_state_reg ( .D(
        new_AGEMA_signal_4267), .CK(clk), .Q(new_AGEMA_signal_4268), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1994_s_current_state_reg ( .D(
        new_AGEMA_signal_4271), .CK(clk), .Q(new_AGEMA_signal_4272), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1998_s_current_state_reg ( .D(
        new_AGEMA_signal_4275), .CK(clk), .Q(new_AGEMA_signal_4276), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2002_s_current_state_reg ( .D(
        new_AGEMA_signal_4279), .CK(clk), .Q(new_AGEMA_signal_4280), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2006_s_current_state_reg ( .D(
        new_AGEMA_signal_4283), .CK(clk), .Q(new_AGEMA_signal_4284), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2010_s_current_state_reg ( .D(
        new_AGEMA_signal_4287), .CK(clk), .Q(new_AGEMA_signal_4288), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2014_s_current_state_reg ( .D(
        new_AGEMA_signal_4291), .CK(clk), .Q(new_AGEMA_signal_4292), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2018_s_current_state_reg ( .D(
        new_AGEMA_signal_4295), .CK(clk), .Q(new_AGEMA_signal_4296), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2022_s_current_state_reg ( .D(
        new_AGEMA_signal_4299), .CK(clk), .Q(new_AGEMA_signal_4300), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2026_s_current_state_reg ( .D(
        new_AGEMA_signal_4303), .CK(clk), .Q(new_AGEMA_signal_4304), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2030_s_current_state_reg ( .D(
        new_AGEMA_signal_4307), .CK(clk), .Q(new_AGEMA_signal_4308), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2034_s_current_state_reg ( .D(
        new_AGEMA_signal_4311), .CK(clk), .Q(new_AGEMA_signal_4312), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2038_s_current_state_reg ( .D(
        new_AGEMA_signal_4315), .CK(clk), .Q(new_AGEMA_signal_4316), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2042_s_current_state_reg ( .D(
        new_AGEMA_signal_4319), .CK(clk), .Q(new_AGEMA_signal_4320), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2046_s_current_state_reg ( .D(
        new_AGEMA_signal_4323), .CK(clk), .Q(new_AGEMA_signal_4324), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2050_s_current_state_reg ( .D(
        new_AGEMA_signal_4327), .CK(clk), .Q(new_AGEMA_signal_4328), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2054_s_current_state_reg ( .D(
        new_AGEMA_signal_4331), .CK(clk), .Q(new_AGEMA_signal_4332), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2058_s_current_state_reg ( .D(
        new_AGEMA_signal_4335), .CK(clk), .Q(new_AGEMA_signal_4336), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2062_s_current_state_reg ( .D(
        new_AGEMA_signal_4339), .CK(clk), .Q(new_AGEMA_signal_4340), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2070_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_T2), .CK(clk), .Q(new_AGEMA_signal_4348), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2072_s_current_state_reg ( .D(
        new_AGEMA_signal_1934), .CK(clk), .Q(new_AGEMA_signal_4350), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2074_s_current_state_reg ( .D(
        new_AGEMA_signal_1935), .CK(clk), .Q(new_AGEMA_signal_4352), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2084_s_current_state_reg ( .D(
        new_AGEMA_signal_4361), .CK(clk), .Q(new_AGEMA_signal_4362), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2088_s_current_state_reg ( .D(
        new_AGEMA_signal_4365), .CK(clk), .Q(new_AGEMA_signal_4366), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2092_s_current_state_reg ( .D(
        new_AGEMA_signal_4369), .CK(clk), .Q(new_AGEMA_signal_4370), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2094_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_YY_1_), .CK(clk), .Q(new_AGEMA_signal_4372), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2096_s_current_state_reg ( .D(
        new_AGEMA_signal_2284), .CK(clk), .Q(new_AGEMA_signal_4374), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2098_s_current_state_reg ( .D(
        new_AGEMA_signal_2285), .CK(clk), .Q(new_AGEMA_signal_4376), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2106_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_T2), .CK(clk), .Q(new_AGEMA_signal_4384), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2108_s_current_state_reg ( .D(
        new_AGEMA_signal_1940), .CK(clk), .Q(new_AGEMA_signal_4386), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2110_s_current_state_reg ( .D(
        new_AGEMA_signal_1941), .CK(clk), .Q(new_AGEMA_signal_4388), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2120_s_current_state_reg ( .D(
        new_AGEMA_signal_4397), .CK(clk), .Q(new_AGEMA_signal_4398), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2124_s_current_state_reg ( .D(
        new_AGEMA_signal_4401), .CK(clk), .Q(new_AGEMA_signal_4402), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2128_s_current_state_reg ( .D(
        new_AGEMA_signal_4405), .CK(clk), .Q(new_AGEMA_signal_4406), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2130_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_YY_1_), .CK(clk), .Q(new_AGEMA_signal_4408), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2132_s_current_state_reg ( .D(
        new_AGEMA_signal_2288), .CK(clk), .Q(new_AGEMA_signal_4410), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2134_s_current_state_reg ( .D(
        new_AGEMA_signal_2289), .CK(clk), .Q(new_AGEMA_signal_4412), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2142_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_T2), .CK(clk), .Q(new_AGEMA_signal_4420), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2144_s_current_state_reg ( .D(
        new_AGEMA_signal_1946), .CK(clk), .Q(new_AGEMA_signal_4422), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2146_s_current_state_reg ( .D(
        new_AGEMA_signal_1947), .CK(clk), .Q(new_AGEMA_signal_4424), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2156_s_current_state_reg ( .D(
        new_AGEMA_signal_4433), .CK(clk), .Q(new_AGEMA_signal_4434), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2160_s_current_state_reg ( .D(
        new_AGEMA_signal_4437), .CK(clk), .Q(new_AGEMA_signal_4438), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2164_s_current_state_reg ( .D(
        new_AGEMA_signal_4441), .CK(clk), .Q(new_AGEMA_signal_4442), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2166_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_YY_1_), .CK(clk), .Q(new_AGEMA_signal_4444), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2168_s_current_state_reg ( .D(
        new_AGEMA_signal_2292), .CK(clk), .Q(new_AGEMA_signal_4446), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2170_s_current_state_reg ( .D(
        new_AGEMA_signal_2293), .CK(clk), .Q(new_AGEMA_signal_4448), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2178_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_T2), .CK(clk), .Q(new_AGEMA_signal_4456), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2180_s_current_state_reg ( .D(
        new_AGEMA_signal_1952), .CK(clk), .Q(new_AGEMA_signal_4458), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2182_s_current_state_reg ( .D(
        new_AGEMA_signal_1953), .CK(clk), .Q(new_AGEMA_signal_4460), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2192_s_current_state_reg ( .D(
        new_AGEMA_signal_4469), .CK(clk), .Q(new_AGEMA_signal_4470), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2196_s_current_state_reg ( .D(
        new_AGEMA_signal_4473), .CK(clk), .Q(new_AGEMA_signal_4474), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2200_s_current_state_reg ( .D(
        new_AGEMA_signal_4477), .CK(clk), .Q(new_AGEMA_signal_4478), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2202_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_YY_1_), .CK(clk), .Q(new_AGEMA_signal_4480), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2204_s_current_state_reg ( .D(
        new_AGEMA_signal_2296), .CK(clk), .Q(new_AGEMA_signal_4482), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2206_s_current_state_reg ( .D(
        new_AGEMA_signal_2297), .CK(clk), .Q(new_AGEMA_signal_4484), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2214_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_T2), .CK(clk), .Q(new_AGEMA_signal_4492), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2216_s_current_state_reg ( .D(
        new_AGEMA_signal_1958), .CK(clk), .Q(new_AGEMA_signal_4494), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2218_s_current_state_reg ( .D(
        new_AGEMA_signal_1959), .CK(clk), .Q(new_AGEMA_signal_4496), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2228_s_current_state_reg ( .D(
        new_AGEMA_signal_4505), .CK(clk), .Q(new_AGEMA_signal_4506), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2232_s_current_state_reg ( .D(
        new_AGEMA_signal_4509), .CK(clk), .Q(new_AGEMA_signal_4510), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2236_s_current_state_reg ( .D(
        new_AGEMA_signal_4513), .CK(clk), .Q(new_AGEMA_signal_4514), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2238_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_YY_1_), .CK(clk), .Q(new_AGEMA_signal_4516), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2240_s_current_state_reg ( .D(
        new_AGEMA_signal_2300), .CK(clk), .Q(new_AGEMA_signal_4518), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2242_s_current_state_reg ( .D(
        new_AGEMA_signal_2301), .CK(clk), .Q(new_AGEMA_signal_4520), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2250_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_T2), .CK(clk), .Q(new_AGEMA_signal_4528), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2252_s_current_state_reg ( .D(
        new_AGEMA_signal_1964), .CK(clk), .Q(new_AGEMA_signal_4530), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2254_s_current_state_reg ( .D(
        new_AGEMA_signal_1965), .CK(clk), .Q(new_AGEMA_signal_4532), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2264_s_current_state_reg ( .D(
        new_AGEMA_signal_4541), .CK(clk), .Q(new_AGEMA_signal_4542), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2268_s_current_state_reg ( .D(
        new_AGEMA_signal_4545), .CK(clk), .Q(new_AGEMA_signal_4546), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2272_s_current_state_reg ( .D(
        new_AGEMA_signal_4549), .CK(clk), .Q(new_AGEMA_signal_4550), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2274_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_YY_1_), .CK(clk), .Q(new_AGEMA_signal_4552), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2276_s_current_state_reg ( .D(
        new_AGEMA_signal_2304), .CK(clk), .Q(new_AGEMA_signal_4554), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2278_s_current_state_reg ( .D(
        new_AGEMA_signal_2305), .CK(clk), .Q(new_AGEMA_signal_4556), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2286_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_T2), .CK(clk), .Q(new_AGEMA_signal_4564), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2288_s_current_state_reg ( .D(
        new_AGEMA_signal_1970), .CK(clk), .Q(new_AGEMA_signal_4566), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2290_s_current_state_reg ( .D(
        new_AGEMA_signal_1971), .CK(clk), .Q(new_AGEMA_signal_4568), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2300_s_current_state_reg ( .D(
        new_AGEMA_signal_4577), .CK(clk), .Q(new_AGEMA_signal_4578), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2304_s_current_state_reg ( .D(
        new_AGEMA_signal_4581), .CK(clk), .Q(new_AGEMA_signal_4582), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2308_s_current_state_reg ( .D(
        new_AGEMA_signal_4585), .CK(clk), .Q(new_AGEMA_signal_4586), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2310_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_YY_1_), .CK(clk), .Q(new_AGEMA_signal_4588), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2312_s_current_state_reg ( .D(
        new_AGEMA_signal_2308), .CK(clk), .Q(new_AGEMA_signal_4590), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2314_s_current_state_reg ( .D(
        new_AGEMA_signal_2309), .CK(clk), .Q(new_AGEMA_signal_4592), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2322_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_T2), .CK(clk), .Q(new_AGEMA_signal_4600), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2324_s_current_state_reg ( .D(
        new_AGEMA_signal_1976), .CK(clk), .Q(new_AGEMA_signal_4602), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2326_s_current_state_reg ( .D(
        new_AGEMA_signal_1977), .CK(clk), .Q(new_AGEMA_signal_4604), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2336_s_current_state_reg ( .D(
        new_AGEMA_signal_4613), .CK(clk), .Q(new_AGEMA_signal_4614), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2340_s_current_state_reg ( .D(
        new_AGEMA_signal_4617), .CK(clk), .Q(new_AGEMA_signal_4618), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2344_s_current_state_reg ( .D(
        new_AGEMA_signal_4621), .CK(clk), .Q(new_AGEMA_signal_4622), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2346_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_YY_1_), .CK(clk), .Q(new_AGEMA_signal_4624), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2348_s_current_state_reg ( .D(
        new_AGEMA_signal_2312), .CK(clk), .Q(new_AGEMA_signal_4626), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2350_s_current_state_reg ( .D(
        new_AGEMA_signal_2313), .CK(clk), .Q(new_AGEMA_signal_4628), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2358_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_T2), .CK(clk), .Q(new_AGEMA_signal_4636), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2360_s_current_state_reg ( .D(
        new_AGEMA_signal_1982), .CK(clk), .Q(new_AGEMA_signal_4638), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2362_s_current_state_reg ( .D(
        new_AGEMA_signal_1983), .CK(clk), .Q(new_AGEMA_signal_4640), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2372_s_current_state_reg ( .D(
        new_AGEMA_signal_4649), .CK(clk), .Q(new_AGEMA_signal_4650), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2376_s_current_state_reg ( .D(
        new_AGEMA_signal_4653), .CK(clk), .Q(new_AGEMA_signal_4654), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2380_s_current_state_reg ( .D(
        new_AGEMA_signal_4657), .CK(clk), .Q(new_AGEMA_signal_4658), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2382_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_YY_1_), .CK(clk), .Q(new_AGEMA_signal_4660), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2384_s_current_state_reg ( .D(
        new_AGEMA_signal_2316), .CK(clk), .Q(new_AGEMA_signal_4662), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2386_s_current_state_reg ( .D(
        new_AGEMA_signal_2317), .CK(clk), .Q(new_AGEMA_signal_4664), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2394_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_T2), .CK(clk), .Q(new_AGEMA_signal_4672), .QN()
         );
  DFF_X1 new_AGEMA_reg_buffer_2396_s_current_state_reg ( .D(
        new_AGEMA_signal_1988), .CK(clk), .Q(new_AGEMA_signal_4674), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2398_s_current_state_reg ( .D(
        new_AGEMA_signal_1989), .CK(clk), .Q(new_AGEMA_signal_4676), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2408_s_current_state_reg ( .D(
        new_AGEMA_signal_4685), .CK(clk), .Q(new_AGEMA_signal_4686), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2412_s_current_state_reg ( .D(
        new_AGEMA_signal_4689), .CK(clk), .Q(new_AGEMA_signal_4690), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2416_s_current_state_reg ( .D(
        new_AGEMA_signal_4693), .CK(clk), .Q(new_AGEMA_signal_4694), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2418_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_YY_1_), .CK(clk), .Q(new_AGEMA_signal_4696), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2420_s_current_state_reg ( .D(
        new_AGEMA_signal_2320), .CK(clk), .Q(new_AGEMA_signal_4698), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2422_s_current_state_reg ( .D(
        new_AGEMA_signal_2321), .CK(clk), .Q(new_AGEMA_signal_4700), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2430_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_T2), .CK(clk), .Q(new_AGEMA_signal_4708), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2432_s_current_state_reg ( .D(
        new_AGEMA_signal_1994), .CK(clk), .Q(new_AGEMA_signal_4710), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2434_s_current_state_reg ( .D(
        new_AGEMA_signal_1995), .CK(clk), .Q(new_AGEMA_signal_4712), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2444_s_current_state_reg ( .D(
        new_AGEMA_signal_4721), .CK(clk), .Q(new_AGEMA_signal_4722), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2448_s_current_state_reg ( .D(
        new_AGEMA_signal_4725), .CK(clk), .Q(new_AGEMA_signal_4726), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2452_s_current_state_reg ( .D(
        new_AGEMA_signal_4729), .CK(clk), .Q(new_AGEMA_signal_4730), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2454_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_YY_1_), .CK(clk), .Q(new_AGEMA_signal_4732), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2456_s_current_state_reg ( .D(
        new_AGEMA_signal_2324), .CK(clk), .Q(new_AGEMA_signal_4734), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2458_s_current_state_reg ( .D(
        new_AGEMA_signal_2325), .CK(clk), .Q(new_AGEMA_signal_4736), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2466_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_T2), .CK(clk), .Q(new_AGEMA_signal_4744), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2468_s_current_state_reg ( .D(
        new_AGEMA_signal_2000), .CK(clk), .Q(new_AGEMA_signal_4746), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2470_s_current_state_reg ( .D(
        new_AGEMA_signal_2001), .CK(clk), .Q(new_AGEMA_signal_4748), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2480_s_current_state_reg ( .D(
        new_AGEMA_signal_4757), .CK(clk), .Q(new_AGEMA_signal_4758), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2484_s_current_state_reg ( .D(
        new_AGEMA_signal_4761), .CK(clk), .Q(new_AGEMA_signal_4762), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2488_s_current_state_reg ( .D(
        new_AGEMA_signal_4765), .CK(clk), .Q(new_AGEMA_signal_4766), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2490_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_YY_1_), .CK(clk), .Q(new_AGEMA_signal_4768), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2492_s_current_state_reg ( .D(
        new_AGEMA_signal_2328), .CK(clk), .Q(new_AGEMA_signal_4770), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2494_s_current_state_reg ( .D(
        new_AGEMA_signal_2329), .CK(clk), .Q(new_AGEMA_signal_4772), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2502_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_T2), .CK(clk), .Q(new_AGEMA_signal_4780), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2504_s_current_state_reg ( .D(
        new_AGEMA_signal_2006), .CK(clk), .Q(new_AGEMA_signal_4782), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2506_s_current_state_reg ( .D(
        new_AGEMA_signal_2007), .CK(clk), .Q(new_AGEMA_signal_4784), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2516_s_current_state_reg ( .D(
        new_AGEMA_signal_4793), .CK(clk), .Q(new_AGEMA_signal_4794), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2520_s_current_state_reg ( .D(
        new_AGEMA_signal_4797), .CK(clk), .Q(new_AGEMA_signal_4798), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2524_s_current_state_reg ( .D(
        new_AGEMA_signal_4801), .CK(clk), .Q(new_AGEMA_signal_4802), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2526_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_YY_1_), .CK(clk), .Q(new_AGEMA_signal_4804), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2528_s_current_state_reg ( .D(
        new_AGEMA_signal_2332), .CK(clk), .Q(new_AGEMA_signal_4806), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2530_s_current_state_reg ( .D(
        new_AGEMA_signal_2333), .CK(clk), .Q(new_AGEMA_signal_4808), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2538_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_T2), .CK(clk), .Q(new_AGEMA_signal_4816), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2540_s_current_state_reg ( .D(
        new_AGEMA_signal_2012), .CK(clk), .Q(new_AGEMA_signal_4818), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2542_s_current_state_reg ( .D(
        new_AGEMA_signal_2013), .CK(clk), .Q(new_AGEMA_signal_4820), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2552_s_current_state_reg ( .D(
        new_AGEMA_signal_4829), .CK(clk), .Q(new_AGEMA_signal_4830), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2556_s_current_state_reg ( .D(
        new_AGEMA_signal_4833), .CK(clk), .Q(new_AGEMA_signal_4834), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2560_s_current_state_reg ( .D(
        new_AGEMA_signal_4837), .CK(clk), .Q(new_AGEMA_signal_4838), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2562_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_YY_1_), .CK(clk), .Q(new_AGEMA_signal_4840), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2564_s_current_state_reg ( .D(
        new_AGEMA_signal_2336), .CK(clk), .Q(new_AGEMA_signal_4842), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2566_s_current_state_reg ( .D(
        new_AGEMA_signal_2337), .CK(clk), .Q(new_AGEMA_signal_4844), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2574_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_T2), .CK(clk), .Q(new_AGEMA_signal_4852), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2576_s_current_state_reg ( .D(
        new_AGEMA_signal_2018), .CK(clk), .Q(new_AGEMA_signal_4854), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2578_s_current_state_reg ( .D(
        new_AGEMA_signal_2019), .CK(clk), .Q(new_AGEMA_signal_4856), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2588_s_current_state_reg ( .D(
        new_AGEMA_signal_4865), .CK(clk), .Q(new_AGEMA_signal_4866), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2592_s_current_state_reg ( .D(
        new_AGEMA_signal_4869), .CK(clk), .Q(new_AGEMA_signal_4870), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2596_s_current_state_reg ( .D(
        new_AGEMA_signal_4873), .CK(clk), .Q(new_AGEMA_signal_4874), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2598_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_YY_1_), .CK(clk), .Q(new_AGEMA_signal_4876), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2600_s_current_state_reg ( .D(
        new_AGEMA_signal_2340), .CK(clk), .Q(new_AGEMA_signal_4878), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2602_s_current_state_reg ( .D(
        new_AGEMA_signal_2341), .CK(clk), .Q(new_AGEMA_signal_4880), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2610_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_T2), .CK(clk), .Q(new_AGEMA_signal_4888), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2612_s_current_state_reg ( .D(
        new_AGEMA_signal_2024), .CK(clk), .Q(new_AGEMA_signal_4890), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2614_s_current_state_reg ( .D(
        new_AGEMA_signal_2025), .CK(clk), .Q(new_AGEMA_signal_4892), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2624_s_current_state_reg ( .D(
        new_AGEMA_signal_4901), .CK(clk), .Q(new_AGEMA_signal_4902), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2628_s_current_state_reg ( .D(
        new_AGEMA_signal_4905), .CK(clk), .Q(new_AGEMA_signal_4906), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2632_s_current_state_reg ( .D(
        new_AGEMA_signal_4909), .CK(clk), .Q(new_AGEMA_signal_4910), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2634_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_YY_1_), .CK(clk), .Q(new_AGEMA_signal_4912), 
        .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2636_s_current_state_reg ( .D(
        new_AGEMA_signal_2344), .CK(clk), .Q(new_AGEMA_signal_4914), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2638_s_current_state_reg ( .D(
        new_AGEMA_signal_2345), .CK(clk), .Q(new_AGEMA_signal_4916), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2642_s_current_state_reg ( .D(
        new_AGEMA_signal_4919), .CK(clk), .Q(new_AGEMA_signal_4920), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2646_s_current_state_reg ( .D(
        new_AGEMA_signal_4923), .CK(clk), .Q(new_AGEMA_signal_4924), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2650_s_current_state_reg ( .D(
        new_AGEMA_signal_4927), .CK(clk), .Q(new_AGEMA_signal_4928), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2654_s_current_state_reg ( .D(
        new_AGEMA_signal_4931), .CK(clk), .Q(new_AGEMA_signal_4932), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2658_s_current_state_reg ( .D(
        new_AGEMA_signal_4935), .CK(clk), .Q(new_AGEMA_signal_4936), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2662_s_current_state_reg ( .D(
        new_AGEMA_signal_4939), .CK(clk), .Q(new_AGEMA_signal_4940), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2666_s_current_state_reg ( .D(
        new_AGEMA_signal_4943), .CK(clk), .Q(new_AGEMA_signal_4944), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2670_s_current_state_reg ( .D(
        new_AGEMA_signal_4947), .CK(clk), .Q(new_AGEMA_signal_4948), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2674_s_current_state_reg ( .D(
        new_AGEMA_signal_4951), .CK(clk), .Q(new_AGEMA_signal_4952), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2678_s_current_state_reg ( .D(
        new_AGEMA_signal_4955), .CK(clk), .Q(new_AGEMA_signal_4956), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2682_s_current_state_reg ( .D(
        new_AGEMA_signal_4959), .CK(clk), .Q(new_AGEMA_signal_4960), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2686_s_current_state_reg ( .D(
        new_AGEMA_signal_4963), .CK(clk), .Q(new_AGEMA_signal_4964), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2690_s_current_state_reg ( .D(
        new_AGEMA_signal_4967), .CK(clk), .Q(new_AGEMA_signal_4968), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2694_s_current_state_reg ( .D(
        new_AGEMA_signal_4971), .CK(clk), .Q(new_AGEMA_signal_4972), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2698_s_current_state_reg ( .D(
        new_AGEMA_signal_4975), .CK(clk), .Q(new_AGEMA_signal_4976), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2702_s_current_state_reg ( .D(
        new_AGEMA_signal_4979), .CK(clk), .Q(new_AGEMA_signal_4980), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2706_s_current_state_reg ( .D(
        new_AGEMA_signal_4983), .CK(clk), .Q(new_AGEMA_signal_4984), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2710_s_current_state_reg ( .D(
        new_AGEMA_signal_4987), .CK(clk), .Q(new_AGEMA_signal_4988), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2714_s_current_state_reg ( .D(
        new_AGEMA_signal_4991), .CK(clk), .Q(new_AGEMA_signal_4992), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2718_s_current_state_reg ( .D(
        new_AGEMA_signal_4995), .CK(clk), .Q(new_AGEMA_signal_4996), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2722_s_current_state_reg ( .D(
        new_AGEMA_signal_4999), .CK(clk), .Q(new_AGEMA_signal_5000), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2726_s_current_state_reg ( .D(
        new_AGEMA_signal_5003), .CK(clk), .Q(new_AGEMA_signal_5004), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2730_s_current_state_reg ( .D(
        new_AGEMA_signal_5007), .CK(clk), .Q(new_AGEMA_signal_5008), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2734_s_current_state_reg ( .D(
        new_AGEMA_signal_5011), .CK(clk), .Q(new_AGEMA_signal_5012), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2738_s_current_state_reg ( .D(
        new_AGEMA_signal_5015), .CK(clk), .Q(new_AGEMA_signal_5016), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2742_s_current_state_reg ( .D(
        new_AGEMA_signal_5019), .CK(clk), .Q(new_AGEMA_signal_5020), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2746_s_current_state_reg ( .D(
        new_AGEMA_signal_5023), .CK(clk), .Q(new_AGEMA_signal_5024), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2750_s_current_state_reg ( .D(
        new_AGEMA_signal_5027), .CK(clk), .Q(new_AGEMA_signal_5028), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2754_s_current_state_reg ( .D(
        new_AGEMA_signal_5031), .CK(clk), .Q(new_AGEMA_signal_5032), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2758_s_current_state_reg ( .D(
        new_AGEMA_signal_5035), .CK(clk), .Q(new_AGEMA_signal_5036), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2762_s_current_state_reg ( .D(
        new_AGEMA_signal_5039), .CK(clk), .Q(new_AGEMA_signal_5040), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2766_s_current_state_reg ( .D(
        new_AGEMA_signal_5043), .CK(clk), .Q(new_AGEMA_signal_5044), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2770_s_current_state_reg ( .D(
        new_AGEMA_signal_5047), .CK(clk), .Q(new_AGEMA_signal_5048), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2774_s_current_state_reg ( .D(
        new_AGEMA_signal_5051), .CK(clk), .Q(new_AGEMA_signal_5052), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2778_s_current_state_reg ( .D(
        new_AGEMA_signal_5055), .CK(clk), .Q(new_AGEMA_signal_5056), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2782_s_current_state_reg ( .D(
        new_AGEMA_signal_5059), .CK(clk), .Q(new_AGEMA_signal_5060), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2786_s_current_state_reg ( .D(
        new_AGEMA_signal_5063), .CK(clk), .Q(new_AGEMA_signal_5064), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2790_s_current_state_reg ( .D(
        new_AGEMA_signal_5067), .CK(clk), .Q(new_AGEMA_signal_5068), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2794_s_current_state_reg ( .D(
        new_AGEMA_signal_5071), .CK(clk), .Q(new_AGEMA_signal_5072), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2798_s_current_state_reg ( .D(
        new_AGEMA_signal_5075), .CK(clk), .Q(new_AGEMA_signal_5076), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2802_s_current_state_reg ( .D(
        new_AGEMA_signal_5079), .CK(clk), .Q(new_AGEMA_signal_5080), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2806_s_current_state_reg ( .D(
        new_AGEMA_signal_5083), .CK(clk), .Q(new_AGEMA_signal_5084), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2810_s_current_state_reg ( .D(
        new_AGEMA_signal_5087), .CK(clk), .Q(new_AGEMA_signal_5088), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2814_s_current_state_reg ( .D(
        new_AGEMA_signal_5091), .CK(clk), .Q(new_AGEMA_signal_5092), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2818_s_current_state_reg ( .D(
        new_AGEMA_signal_5095), .CK(clk), .Q(new_AGEMA_signal_5096), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2822_s_current_state_reg ( .D(
        new_AGEMA_signal_5099), .CK(clk), .Q(new_AGEMA_signal_5100), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2826_s_current_state_reg ( .D(
        new_AGEMA_signal_5103), .CK(clk), .Q(new_AGEMA_signal_5104), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2830_s_current_state_reg ( .D(
        new_AGEMA_signal_5107), .CK(clk), .Q(new_AGEMA_signal_5108), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2834_s_current_state_reg ( .D(
        new_AGEMA_signal_5111), .CK(clk), .Q(new_AGEMA_signal_5112), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2838_s_current_state_reg ( .D(
        new_AGEMA_signal_5115), .CK(clk), .Q(new_AGEMA_signal_5116), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2842_s_current_state_reg ( .D(
        new_AGEMA_signal_5119), .CK(clk), .Q(new_AGEMA_signal_5120), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2846_s_current_state_reg ( .D(
        new_AGEMA_signal_5123), .CK(clk), .Q(new_AGEMA_signal_5124), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2848_s_current_state_reg ( .D(StateRegInput[63]), 
        .CK(clk), .Q(new_AGEMA_signal_5126), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2850_s_current_state_reg ( .D(
        new_AGEMA_signal_3042), .CK(clk), .Q(new_AGEMA_signal_5128), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2852_s_current_state_reg ( .D(
        new_AGEMA_signal_3043), .CK(clk), .Q(new_AGEMA_signal_5130), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2854_s_current_state_reg ( .D(StateRegInput[62]), 
        .CK(clk), .Q(new_AGEMA_signal_5132), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2856_s_current_state_reg ( .D(
        new_AGEMA_signal_2956), .CK(clk), .Q(new_AGEMA_signal_5134), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2858_s_current_state_reg ( .D(
        new_AGEMA_signal_2957), .CK(clk), .Q(new_AGEMA_signal_5136), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2860_s_current_state_reg ( .D(StateRegInput[59]), 
        .CK(clk), .Q(new_AGEMA_signal_5138), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2862_s_current_state_reg ( .D(
        new_AGEMA_signal_2848), .CK(clk), .Q(new_AGEMA_signal_5140), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2864_s_current_state_reg ( .D(
        new_AGEMA_signal_2849), .CK(clk), .Q(new_AGEMA_signal_5142), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2866_s_current_state_reg ( .D(StateRegInput[58]), 
        .CK(clk), .Q(new_AGEMA_signal_5144), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2868_s_current_state_reg ( .D(
        new_AGEMA_signal_2728), .CK(clk), .Q(new_AGEMA_signal_5146), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2870_s_current_state_reg ( .D(
        new_AGEMA_signal_2729), .CK(clk), .Q(new_AGEMA_signal_5148), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2872_s_current_state_reg ( .D(StateRegInput[55]), 
        .CK(clk), .Q(new_AGEMA_signal_5150), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2874_s_current_state_reg ( .D(
        new_AGEMA_signal_2844), .CK(clk), .Q(new_AGEMA_signal_5152), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2876_s_current_state_reg ( .D(
        new_AGEMA_signal_2845), .CK(clk), .Q(new_AGEMA_signal_5154), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2878_s_current_state_reg ( .D(StateRegInput[54]), 
        .CK(clk), .Q(new_AGEMA_signal_5156), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2880_s_current_state_reg ( .D(
        new_AGEMA_signal_2724), .CK(clk), .Q(new_AGEMA_signal_5158), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2882_s_current_state_reg ( .D(
        new_AGEMA_signal_2725), .CK(clk), .Q(new_AGEMA_signal_5160), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2884_s_current_state_reg ( .D(StateRegInput[51]), 
        .CK(clk), .Q(new_AGEMA_signal_5162), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2886_s_current_state_reg ( .D(
        new_AGEMA_signal_2840), .CK(clk), .Q(new_AGEMA_signal_5164), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2888_s_current_state_reg ( .D(
        new_AGEMA_signal_2841), .CK(clk), .Q(new_AGEMA_signal_5166), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2890_s_current_state_reg ( .D(StateRegInput[50]), 
        .CK(clk), .Q(new_AGEMA_signal_5168), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2892_s_current_state_reg ( .D(
        new_AGEMA_signal_2720), .CK(clk), .Q(new_AGEMA_signal_5170), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2894_s_current_state_reg ( .D(
        new_AGEMA_signal_2721), .CK(clk), .Q(new_AGEMA_signal_5172), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2896_s_current_state_reg ( .D(StateRegInput[47]), 
        .CK(clk), .Q(new_AGEMA_signal_5174), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2898_s_current_state_reg ( .D(
        new_AGEMA_signal_2836), .CK(clk), .Q(new_AGEMA_signal_5176), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2900_s_current_state_reg ( .D(
        new_AGEMA_signal_2837), .CK(clk), .Q(new_AGEMA_signal_5178), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2902_s_current_state_reg ( .D(StateRegInput[46]), 
        .CK(clk), .Q(new_AGEMA_signal_5180), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2904_s_current_state_reg ( .D(
        new_AGEMA_signal_2716), .CK(clk), .Q(new_AGEMA_signal_5182), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2906_s_current_state_reg ( .D(
        new_AGEMA_signal_2717), .CK(clk), .Q(new_AGEMA_signal_5184), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2908_s_current_state_reg ( .D(StateRegInput[43]), 
        .CK(clk), .Q(new_AGEMA_signal_5186), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2910_s_current_state_reg ( .D(
        new_AGEMA_signal_2592), .CK(clk), .Q(new_AGEMA_signal_5188), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2912_s_current_state_reg ( .D(
        new_AGEMA_signal_2593), .CK(clk), .Q(new_AGEMA_signal_5190), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2914_s_current_state_reg ( .D(StateRegInput[42]), 
        .CK(clk), .Q(new_AGEMA_signal_5192), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2916_s_current_state_reg ( .D(
        new_AGEMA_signal_2486), .CK(clk), .Q(new_AGEMA_signal_5194), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2918_s_current_state_reg ( .D(
        new_AGEMA_signal_2487), .CK(clk), .Q(new_AGEMA_signal_5196), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2920_s_current_state_reg ( .D(StateRegInput[39]), 
        .CK(clk), .Q(new_AGEMA_signal_5198), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2922_s_current_state_reg ( .D(
        new_AGEMA_signal_2588), .CK(clk), .Q(new_AGEMA_signal_5200), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2924_s_current_state_reg ( .D(
        new_AGEMA_signal_2589), .CK(clk), .Q(new_AGEMA_signal_5202), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2926_s_current_state_reg ( .D(StateRegInput[38]), 
        .CK(clk), .Q(new_AGEMA_signal_5204), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2928_s_current_state_reg ( .D(
        new_AGEMA_signal_2482), .CK(clk), .Q(new_AGEMA_signal_5206), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2930_s_current_state_reg ( .D(
        new_AGEMA_signal_2483), .CK(clk), .Q(new_AGEMA_signal_5208), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2932_s_current_state_reg ( .D(StateRegInput[35]), 
        .CK(clk), .Q(new_AGEMA_signal_5210), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2934_s_current_state_reg ( .D(
        new_AGEMA_signal_2584), .CK(clk), .Q(new_AGEMA_signal_5212), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2936_s_current_state_reg ( .D(
        new_AGEMA_signal_2585), .CK(clk), .Q(new_AGEMA_signal_5214), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2938_s_current_state_reg ( .D(StateRegInput[34]), 
        .CK(clk), .Q(new_AGEMA_signal_5216), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2940_s_current_state_reg ( .D(
        new_AGEMA_signal_2478), .CK(clk), .Q(new_AGEMA_signal_5218), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2942_s_current_state_reg ( .D(
        new_AGEMA_signal_2479), .CK(clk), .Q(new_AGEMA_signal_5220), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2944_s_current_state_reg ( .D(StateRegInput[31]), 
        .CK(clk), .Q(new_AGEMA_signal_5222), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2946_s_current_state_reg ( .D(
        new_AGEMA_signal_2820), .CK(clk), .Q(new_AGEMA_signal_5224), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2948_s_current_state_reg ( .D(
        new_AGEMA_signal_2821), .CK(clk), .Q(new_AGEMA_signal_5226), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2950_s_current_state_reg ( .D(StateRegInput[30]), 
        .CK(clk), .Q(new_AGEMA_signal_5228), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2952_s_current_state_reg ( .D(
        new_AGEMA_signal_2700), .CK(clk), .Q(new_AGEMA_signal_5230), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2954_s_current_state_reg ( .D(
        new_AGEMA_signal_2701), .CK(clk), .Q(new_AGEMA_signal_5232), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2956_s_current_state_reg ( .D(StateRegInput[27]), 
        .CK(clk), .Q(new_AGEMA_signal_5234), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2958_s_current_state_reg ( .D(
        new_AGEMA_signal_3018), .CK(clk), .Q(new_AGEMA_signal_5236), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2960_s_current_state_reg ( .D(
        new_AGEMA_signal_3019), .CK(clk), .Q(new_AGEMA_signal_5238), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2962_s_current_state_reg ( .D(StateRegInput[26]), 
        .CK(clk), .Q(new_AGEMA_signal_5240), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2964_s_current_state_reg ( .D(
        new_AGEMA_signal_2932), .CK(clk), .Q(new_AGEMA_signal_5242), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2966_s_current_state_reg ( .D(
        new_AGEMA_signal_2933), .CK(clk), .Q(new_AGEMA_signal_5244), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2968_s_current_state_reg ( .D(StateRegInput[23]), 
        .CK(clk), .Q(new_AGEMA_signal_5246), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2970_s_current_state_reg ( .D(
        new_AGEMA_signal_2816), .CK(clk), .Q(new_AGEMA_signal_5248), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2972_s_current_state_reg ( .D(
        new_AGEMA_signal_2817), .CK(clk), .Q(new_AGEMA_signal_5250), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2974_s_current_state_reg ( .D(StateRegInput[22]), 
        .CK(clk), .Q(new_AGEMA_signal_5252), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2976_s_current_state_reg ( .D(
        new_AGEMA_signal_2696), .CK(clk), .Q(new_AGEMA_signal_5254), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2978_s_current_state_reg ( .D(
        new_AGEMA_signal_2697), .CK(clk), .Q(new_AGEMA_signal_5256), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2980_s_current_state_reg ( .D(StateRegInput[19]), 
        .CK(clk), .Q(new_AGEMA_signal_5258), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2982_s_current_state_reg ( .D(
        new_AGEMA_signal_2812), .CK(clk), .Q(new_AGEMA_signal_5260), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2984_s_current_state_reg ( .D(
        new_AGEMA_signal_2813), .CK(clk), .Q(new_AGEMA_signal_5262), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2986_s_current_state_reg ( .D(StateRegInput[18]), 
        .CK(clk), .Q(new_AGEMA_signal_5264), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2988_s_current_state_reg ( .D(
        new_AGEMA_signal_2692), .CK(clk), .Q(new_AGEMA_signal_5266), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2990_s_current_state_reg ( .D(
        new_AGEMA_signal_2693), .CK(clk), .Q(new_AGEMA_signal_5268), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2992_s_current_state_reg ( .D(StateRegInput[15]), 
        .CK(clk), .Q(new_AGEMA_signal_5270), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2994_s_current_state_reg ( .D(
        new_AGEMA_signal_3006), .CK(clk), .Q(new_AGEMA_signal_5272), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2996_s_current_state_reg ( .D(
        new_AGEMA_signal_3007), .CK(clk), .Q(new_AGEMA_signal_5274), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2998_s_current_state_reg ( .D(StateRegInput[14]), 
        .CK(clk), .Q(new_AGEMA_signal_5276), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3000_s_current_state_reg ( .D(
        new_AGEMA_signal_2920), .CK(clk), .Q(new_AGEMA_signal_5278), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3002_s_current_state_reg ( .D(
        new_AGEMA_signal_2921), .CK(clk), .Q(new_AGEMA_signal_5280), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3004_s_current_state_reg ( .D(StateRegInput[11]), 
        .CK(clk), .Q(new_AGEMA_signal_5282), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3006_s_current_state_reg ( .D(
        new_AGEMA_signal_2808), .CK(clk), .Q(new_AGEMA_signal_5284), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3008_s_current_state_reg ( .D(
        new_AGEMA_signal_2809), .CK(clk), .Q(new_AGEMA_signal_5286), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3010_s_current_state_reg ( .D(StateRegInput[10]), 
        .CK(clk), .Q(new_AGEMA_signal_5288), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3012_s_current_state_reg ( .D(
        new_AGEMA_signal_2688), .CK(clk), .Q(new_AGEMA_signal_5290), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3014_s_current_state_reg ( .D(
        new_AGEMA_signal_2689), .CK(clk), .Q(new_AGEMA_signal_5292), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3016_s_current_state_reg ( .D(StateRegInput[7]), 
        .CK(clk), .Q(new_AGEMA_signal_5294), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3018_s_current_state_reg ( .D(
        new_AGEMA_signal_2804), .CK(clk), .Q(new_AGEMA_signal_5296), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3020_s_current_state_reg ( .D(
        new_AGEMA_signal_2805), .CK(clk), .Q(new_AGEMA_signal_5298), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3022_s_current_state_reg ( .D(StateRegInput[6]), 
        .CK(clk), .Q(new_AGEMA_signal_5300), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3024_s_current_state_reg ( .D(
        new_AGEMA_signal_2684), .CK(clk), .Q(new_AGEMA_signal_5302), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3026_s_current_state_reg ( .D(
        new_AGEMA_signal_2685), .CK(clk), .Q(new_AGEMA_signal_5304), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3028_s_current_state_reg ( .D(StateRegInput[3]), 
        .CK(clk), .Q(new_AGEMA_signal_5306), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3030_s_current_state_reg ( .D(
        new_AGEMA_signal_2800), .CK(clk), .Q(new_AGEMA_signal_5308), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3032_s_current_state_reg ( .D(
        new_AGEMA_signal_2801), .CK(clk), .Q(new_AGEMA_signal_5310), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3034_s_current_state_reg ( .D(StateRegInput[2]), 
        .CK(clk), .Q(new_AGEMA_signal_5312), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3036_s_current_state_reg ( .D(
        new_AGEMA_signal_2680), .CK(clk), .Q(new_AGEMA_signal_5314), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3038_s_current_state_reg ( .D(
        new_AGEMA_signal_2681), .CK(clk), .Q(new_AGEMA_signal_5316), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3042_s_current_state_reg ( .D(
        new_AGEMA_signal_5319), .CK(clk), .Q(new_AGEMA_signal_5320), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3046_s_current_state_reg ( .D(
        new_AGEMA_signal_5323), .CK(clk), .Q(new_AGEMA_signal_5324), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3050_s_current_state_reg ( .D(
        new_AGEMA_signal_5327), .CK(clk), .Q(new_AGEMA_signal_5328), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3054_s_current_state_reg ( .D(
        new_AGEMA_signal_5331), .CK(clk), .Q(new_AGEMA_signal_5332), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3058_s_current_state_reg ( .D(
        new_AGEMA_signal_5335), .CK(clk), .Q(new_AGEMA_signal_5336), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3062_s_current_state_reg ( .D(
        new_AGEMA_signal_5339), .CK(clk), .Q(new_AGEMA_signal_5340), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3066_s_current_state_reg ( .D(
        new_AGEMA_signal_5343), .CK(clk), .Q(new_AGEMA_signal_5344), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3070_s_current_state_reg ( .D(
        new_AGEMA_signal_5347), .CK(clk), .Q(new_AGEMA_signal_5348), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3074_s_current_state_reg ( .D(
        new_AGEMA_signal_5351), .CK(clk), .Q(new_AGEMA_signal_5352), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3078_s_current_state_reg ( .D(
        new_AGEMA_signal_5355), .CK(clk), .Q(new_AGEMA_signal_5356), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3082_s_current_state_reg ( .D(
        new_AGEMA_signal_5359), .CK(clk), .Q(new_AGEMA_signal_5360), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3086_s_current_state_reg ( .D(
        new_AGEMA_signal_5363), .CK(clk), .Q(new_AGEMA_signal_5364), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3090_s_current_state_reg ( .D(
        new_AGEMA_signal_5367), .CK(clk), .Q(new_AGEMA_signal_5368), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3094_s_current_state_reg ( .D(
        new_AGEMA_signal_5371), .CK(clk), .Q(new_AGEMA_signal_5372), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3098_s_current_state_reg ( .D(
        new_AGEMA_signal_5375), .CK(clk), .Q(new_AGEMA_signal_5376), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3102_s_current_state_reg ( .D(
        new_AGEMA_signal_5379), .CK(clk), .Q(new_AGEMA_signal_5380), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3106_s_current_state_reg ( .D(
        new_AGEMA_signal_5383), .CK(clk), .Q(new_AGEMA_signal_5384), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3110_s_current_state_reg ( .D(
        new_AGEMA_signal_5387), .CK(clk), .Q(new_AGEMA_signal_5388), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3114_s_current_state_reg ( .D(
        new_AGEMA_signal_5391), .CK(clk), .Q(new_AGEMA_signal_5392), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3118_s_current_state_reg ( .D(
        new_AGEMA_signal_5395), .CK(clk), .Q(new_AGEMA_signal_5396), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3122_s_current_state_reg ( .D(
        new_AGEMA_signal_5399), .CK(clk), .Q(new_AGEMA_signal_5400), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3126_s_current_state_reg ( .D(
        new_AGEMA_signal_5403), .CK(clk), .Q(new_AGEMA_signal_5404), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3130_s_current_state_reg ( .D(
        new_AGEMA_signal_5407), .CK(clk), .Q(new_AGEMA_signal_5408), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3134_s_current_state_reg ( .D(
        new_AGEMA_signal_5411), .CK(clk), .Q(new_AGEMA_signal_5412), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3138_s_current_state_reg ( .D(
        new_AGEMA_signal_5415), .CK(clk), .Q(new_AGEMA_signal_5416), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3142_s_current_state_reg ( .D(
        new_AGEMA_signal_5419), .CK(clk), .Q(new_AGEMA_signal_5420), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3146_s_current_state_reg ( .D(
        new_AGEMA_signal_5423), .CK(clk), .Q(new_AGEMA_signal_5424), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3150_s_current_state_reg ( .D(
        new_AGEMA_signal_5427), .CK(clk), .Q(new_AGEMA_signal_5428), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3154_s_current_state_reg ( .D(
        new_AGEMA_signal_5431), .CK(clk), .Q(new_AGEMA_signal_5432), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3158_s_current_state_reg ( .D(
        new_AGEMA_signal_5435), .CK(clk), .Q(new_AGEMA_signal_5436), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3162_s_current_state_reg ( .D(
        new_AGEMA_signal_5439), .CK(clk), .Q(new_AGEMA_signal_5440), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3166_s_current_state_reg ( .D(
        new_AGEMA_signal_5443), .CK(clk), .Q(new_AGEMA_signal_5444), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3170_s_current_state_reg ( .D(
        new_AGEMA_signal_5447), .CK(clk), .Q(new_AGEMA_signal_5448), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3174_s_current_state_reg ( .D(
        new_AGEMA_signal_5451), .CK(clk), .Q(new_AGEMA_signal_5452), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3178_s_current_state_reg ( .D(
        new_AGEMA_signal_5455), .CK(clk), .Q(new_AGEMA_signal_5456), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3182_s_current_state_reg ( .D(
        new_AGEMA_signal_5459), .CK(clk), .Q(new_AGEMA_signal_5460), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3186_s_current_state_reg ( .D(
        new_AGEMA_signal_5463), .CK(clk), .Q(new_AGEMA_signal_5464), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3190_s_current_state_reg ( .D(
        new_AGEMA_signal_5467), .CK(clk), .Q(new_AGEMA_signal_5468), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3194_s_current_state_reg ( .D(
        new_AGEMA_signal_5471), .CK(clk), .Q(new_AGEMA_signal_5472), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3198_s_current_state_reg ( .D(
        new_AGEMA_signal_5475), .CK(clk), .Q(new_AGEMA_signal_5476), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3202_s_current_state_reg ( .D(
        new_AGEMA_signal_5479), .CK(clk), .Q(new_AGEMA_signal_5480), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3206_s_current_state_reg ( .D(
        new_AGEMA_signal_5483), .CK(clk), .Q(new_AGEMA_signal_5484), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3210_s_current_state_reg ( .D(
        new_AGEMA_signal_5487), .CK(clk), .Q(new_AGEMA_signal_5488), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3214_s_current_state_reg ( .D(
        new_AGEMA_signal_5491), .CK(clk), .Q(new_AGEMA_signal_5492), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3218_s_current_state_reg ( .D(
        new_AGEMA_signal_5495), .CK(clk), .Q(new_AGEMA_signal_5496), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3222_s_current_state_reg ( .D(
        new_AGEMA_signal_5499), .CK(clk), .Q(new_AGEMA_signal_5500), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3226_s_current_state_reg ( .D(
        new_AGEMA_signal_5503), .CK(clk), .Q(new_AGEMA_signal_5504), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3230_s_current_state_reg ( .D(
        new_AGEMA_signal_5507), .CK(clk), .Q(new_AGEMA_signal_5508), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3234_s_current_state_reg ( .D(
        new_AGEMA_signal_5511), .CK(clk), .Q(new_AGEMA_signal_5512), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3238_s_current_state_reg ( .D(
        new_AGEMA_signal_5515), .CK(clk), .Q(new_AGEMA_signal_5516), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3242_s_current_state_reg ( .D(
        new_AGEMA_signal_5519), .CK(clk), .Q(new_AGEMA_signal_5520), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3246_s_current_state_reg ( .D(
        new_AGEMA_signal_5523), .CK(clk), .Q(new_AGEMA_signal_5524), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3250_s_current_state_reg ( .D(
        new_AGEMA_signal_5527), .CK(clk), .Q(new_AGEMA_signal_5528), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3254_s_current_state_reg ( .D(
        new_AGEMA_signal_5531), .CK(clk), .Q(new_AGEMA_signal_5532), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3258_s_current_state_reg ( .D(
        new_AGEMA_signal_5535), .CK(clk), .Q(new_AGEMA_signal_5536), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3262_s_current_state_reg ( .D(
        new_AGEMA_signal_5539), .CK(clk), .Q(new_AGEMA_signal_5540), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3266_s_current_state_reg ( .D(
        new_AGEMA_signal_5543), .CK(clk), .Q(new_AGEMA_signal_5544), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3270_s_current_state_reg ( .D(
        new_AGEMA_signal_5547), .CK(clk), .Q(new_AGEMA_signal_5548), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3274_s_current_state_reg ( .D(
        new_AGEMA_signal_5551), .CK(clk), .Q(new_AGEMA_signal_5552), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3278_s_current_state_reg ( .D(
        new_AGEMA_signal_5555), .CK(clk), .Q(new_AGEMA_signal_5556), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3282_s_current_state_reg ( .D(
        new_AGEMA_signal_5559), .CK(clk), .Q(new_AGEMA_signal_5560), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3286_s_current_state_reg ( .D(
        new_AGEMA_signal_5563), .CK(clk), .Q(new_AGEMA_signal_5564), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3290_s_current_state_reg ( .D(
        new_AGEMA_signal_5567), .CK(clk), .Q(new_AGEMA_signal_5568), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3294_s_current_state_reg ( .D(
        new_AGEMA_signal_5571), .CK(clk), .Q(new_AGEMA_signal_5572), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3298_s_current_state_reg ( .D(
        new_AGEMA_signal_5575), .CK(clk), .Q(new_AGEMA_signal_5576), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3302_s_current_state_reg ( .D(
        new_AGEMA_signal_5579), .CK(clk), .Q(new_AGEMA_signal_5580), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3306_s_current_state_reg ( .D(
        new_AGEMA_signal_5583), .CK(clk), .Q(new_AGEMA_signal_5584), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3310_s_current_state_reg ( .D(
        new_AGEMA_signal_5587), .CK(clk), .Q(new_AGEMA_signal_5588), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3314_s_current_state_reg ( .D(
        new_AGEMA_signal_5591), .CK(clk), .Q(new_AGEMA_signal_5592), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3318_s_current_state_reg ( .D(
        new_AGEMA_signal_5595), .CK(clk), .Q(new_AGEMA_signal_5596), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3322_s_current_state_reg ( .D(
        new_AGEMA_signal_5599), .CK(clk), .Q(new_AGEMA_signal_5600), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3326_s_current_state_reg ( .D(
        new_AGEMA_signal_5603), .CK(clk), .Q(new_AGEMA_signal_5604), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3330_s_current_state_reg ( .D(
        new_AGEMA_signal_5607), .CK(clk), .Q(new_AGEMA_signal_5608), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3334_s_current_state_reg ( .D(
        new_AGEMA_signal_5611), .CK(clk), .Q(new_AGEMA_signal_5612), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3338_s_current_state_reg ( .D(
        new_AGEMA_signal_5615), .CK(clk), .Q(new_AGEMA_signal_5616), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3342_s_current_state_reg ( .D(
        new_AGEMA_signal_5619), .CK(clk), .Q(new_AGEMA_signal_5620), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3346_s_current_state_reg ( .D(
        new_AGEMA_signal_5623), .CK(clk), .Q(new_AGEMA_signal_5624), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3350_s_current_state_reg ( .D(
        new_AGEMA_signal_5627), .CK(clk), .Q(new_AGEMA_signal_5628), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3354_s_current_state_reg ( .D(
        new_AGEMA_signal_5631), .CK(clk), .Q(new_AGEMA_signal_5632), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3358_s_current_state_reg ( .D(
        new_AGEMA_signal_5635), .CK(clk), .Q(new_AGEMA_signal_5636), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3362_s_current_state_reg ( .D(
        new_AGEMA_signal_5639), .CK(clk), .Q(new_AGEMA_signal_5640), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3366_s_current_state_reg ( .D(
        new_AGEMA_signal_5643), .CK(clk), .Q(new_AGEMA_signal_5644), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3370_s_current_state_reg ( .D(
        new_AGEMA_signal_5647), .CK(clk), .Q(new_AGEMA_signal_5648), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3374_s_current_state_reg ( .D(
        new_AGEMA_signal_5651), .CK(clk), .Q(new_AGEMA_signal_5652), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3378_s_current_state_reg ( .D(
        new_AGEMA_signal_5655), .CK(clk), .Q(new_AGEMA_signal_5656), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3382_s_current_state_reg ( .D(
        new_AGEMA_signal_5659), .CK(clk), .Q(new_AGEMA_signal_5660), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3386_s_current_state_reg ( .D(
        new_AGEMA_signal_5663), .CK(clk), .Q(new_AGEMA_signal_5664), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3390_s_current_state_reg ( .D(
        new_AGEMA_signal_5667), .CK(clk), .Q(new_AGEMA_signal_5668), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3394_s_current_state_reg ( .D(
        new_AGEMA_signal_5671), .CK(clk), .Q(new_AGEMA_signal_5672), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3398_s_current_state_reg ( .D(
        new_AGEMA_signal_5675), .CK(clk), .Q(new_AGEMA_signal_5676), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3402_s_current_state_reg ( .D(
        new_AGEMA_signal_5679), .CK(clk), .Q(new_AGEMA_signal_5680), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3406_s_current_state_reg ( .D(
        new_AGEMA_signal_5683), .CK(clk), .Q(new_AGEMA_signal_5684), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3410_s_current_state_reg ( .D(
        new_AGEMA_signal_5687), .CK(clk), .Q(new_AGEMA_signal_5688), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3414_s_current_state_reg ( .D(
        new_AGEMA_signal_5691), .CK(clk), .Q(new_AGEMA_signal_5692), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3418_s_current_state_reg ( .D(
        new_AGEMA_signal_5695), .CK(clk), .Q(new_AGEMA_signal_5696), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3422_s_current_state_reg ( .D(
        new_AGEMA_signal_5699), .CK(clk), .Q(new_AGEMA_signal_5700), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3426_s_current_state_reg ( .D(
        new_AGEMA_signal_5703), .CK(clk), .Q(new_AGEMA_signal_5704), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3430_s_current_state_reg ( .D(
        new_AGEMA_signal_5707), .CK(clk), .Q(new_AGEMA_signal_5708), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3434_s_current_state_reg ( .D(
        new_AGEMA_signal_5711), .CK(clk), .Q(new_AGEMA_signal_5712), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3438_s_current_state_reg ( .D(
        new_AGEMA_signal_5715), .CK(clk), .Q(new_AGEMA_signal_5716), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3442_s_current_state_reg ( .D(
        new_AGEMA_signal_5719), .CK(clk), .Q(new_AGEMA_signal_5720), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3446_s_current_state_reg ( .D(
        new_AGEMA_signal_5723), .CK(clk), .Q(new_AGEMA_signal_5724), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3450_s_current_state_reg ( .D(
        new_AGEMA_signal_5727), .CK(clk), .Q(new_AGEMA_signal_5728), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3454_s_current_state_reg ( .D(
        new_AGEMA_signal_5731), .CK(clk), .Q(new_AGEMA_signal_5732), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3458_s_current_state_reg ( .D(
        new_AGEMA_signal_5735), .CK(clk), .Q(new_AGEMA_signal_5736), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3462_s_current_state_reg ( .D(
        new_AGEMA_signal_5739), .CK(clk), .Q(new_AGEMA_signal_5740), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3466_s_current_state_reg ( .D(
        new_AGEMA_signal_5743), .CK(clk), .Q(new_AGEMA_signal_5744), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3470_s_current_state_reg ( .D(
        new_AGEMA_signal_5747), .CK(clk), .Q(new_AGEMA_signal_5748), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3474_s_current_state_reg ( .D(
        new_AGEMA_signal_5751), .CK(clk), .Q(new_AGEMA_signal_5752), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3478_s_current_state_reg ( .D(
        new_AGEMA_signal_5755), .CK(clk), .Q(new_AGEMA_signal_5756), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3482_s_current_state_reg ( .D(
        new_AGEMA_signal_5759), .CK(clk), .Q(new_AGEMA_signal_5760), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3486_s_current_state_reg ( .D(
        new_AGEMA_signal_5763), .CK(clk), .Q(new_AGEMA_signal_5764), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3490_s_current_state_reg ( .D(
        new_AGEMA_signal_5767), .CK(clk), .Q(new_AGEMA_signal_5768), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3494_s_current_state_reg ( .D(
        new_AGEMA_signal_5771), .CK(clk), .Q(new_AGEMA_signal_5772), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3498_s_current_state_reg ( .D(
        new_AGEMA_signal_5775), .CK(clk), .Q(new_AGEMA_signal_5776), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3502_s_current_state_reg ( .D(
        new_AGEMA_signal_5779), .CK(clk), .Q(new_AGEMA_signal_5780), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3506_s_current_state_reg ( .D(
        new_AGEMA_signal_5783), .CK(clk), .Q(new_AGEMA_signal_5784), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3510_s_current_state_reg ( .D(
        new_AGEMA_signal_5787), .CK(clk), .Q(new_AGEMA_signal_5788), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3514_s_current_state_reg ( .D(
        new_AGEMA_signal_5791), .CK(clk), .Q(new_AGEMA_signal_5792), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3518_s_current_state_reg ( .D(
        new_AGEMA_signal_5795), .CK(clk), .Q(new_AGEMA_signal_5796), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3522_s_current_state_reg ( .D(
        new_AGEMA_signal_5799), .CK(clk), .Q(new_AGEMA_signal_5800), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3526_s_current_state_reg ( .D(
        new_AGEMA_signal_5803), .CK(clk), .Q(new_AGEMA_signal_5804), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3530_s_current_state_reg ( .D(
        new_AGEMA_signal_5807), .CK(clk), .Q(new_AGEMA_signal_5808), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3534_s_current_state_reg ( .D(
        new_AGEMA_signal_5811), .CK(clk), .Q(new_AGEMA_signal_5812), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3538_s_current_state_reg ( .D(
        new_AGEMA_signal_5815), .CK(clk), .Q(new_AGEMA_signal_5816), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3542_s_current_state_reg ( .D(
        new_AGEMA_signal_5819), .CK(clk), .Q(new_AGEMA_signal_5820), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3546_s_current_state_reg ( .D(
        new_AGEMA_signal_5823), .CK(clk), .Q(new_AGEMA_signal_5824), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3550_s_current_state_reg ( .D(
        new_AGEMA_signal_5827), .CK(clk), .Q(new_AGEMA_signal_5828), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3554_s_current_state_reg ( .D(
        new_AGEMA_signal_5831), .CK(clk), .Q(new_AGEMA_signal_5832), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3558_s_current_state_reg ( .D(
        new_AGEMA_signal_5835), .CK(clk), .Q(new_AGEMA_signal_5836), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3562_s_current_state_reg ( .D(
        new_AGEMA_signal_5839), .CK(clk), .Q(new_AGEMA_signal_5840), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3566_s_current_state_reg ( .D(
        new_AGEMA_signal_5843), .CK(clk), .Q(new_AGEMA_signal_5844), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3570_s_current_state_reg ( .D(
        new_AGEMA_signal_5847), .CK(clk), .Q(new_AGEMA_signal_5848), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3574_s_current_state_reg ( .D(
        new_AGEMA_signal_5851), .CK(clk), .Q(new_AGEMA_signal_5852), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3578_s_current_state_reg ( .D(
        new_AGEMA_signal_5855), .CK(clk), .Q(new_AGEMA_signal_5856), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3582_s_current_state_reg ( .D(
        new_AGEMA_signal_5859), .CK(clk), .Q(new_AGEMA_signal_5860), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3586_s_current_state_reg ( .D(
        new_AGEMA_signal_5863), .CK(clk), .Q(new_AGEMA_signal_5864), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3590_s_current_state_reg ( .D(
        new_AGEMA_signal_5867), .CK(clk), .Q(new_AGEMA_signal_5868), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3594_s_current_state_reg ( .D(
        new_AGEMA_signal_5871), .CK(clk), .Q(new_AGEMA_signal_5872), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3598_s_current_state_reg ( .D(
        new_AGEMA_signal_5875), .CK(clk), .Q(new_AGEMA_signal_5876), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3602_s_current_state_reg ( .D(
        new_AGEMA_signal_5879), .CK(clk), .Q(new_AGEMA_signal_5880), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3606_s_current_state_reg ( .D(
        new_AGEMA_signal_5883), .CK(clk), .Q(new_AGEMA_signal_5884), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3610_s_current_state_reg ( .D(
        new_AGEMA_signal_5887), .CK(clk), .Q(new_AGEMA_signal_5888), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3614_s_current_state_reg ( .D(
        new_AGEMA_signal_5891), .CK(clk), .Q(new_AGEMA_signal_5892), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3618_s_current_state_reg ( .D(
        new_AGEMA_signal_5895), .CK(clk), .Q(new_AGEMA_signal_5896), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3622_s_current_state_reg ( .D(
        new_AGEMA_signal_5899), .CK(clk), .Q(new_AGEMA_signal_5900), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3626_s_current_state_reg ( .D(
        new_AGEMA_signal_5903), .CK(clk), .Q(new_AGEMA_signal_5904), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3630_s_current_state_reg ( .D(
        new_AGEMA_signal_5907), .CK(clk), .Q(new_AGEMA_signal_5908), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3634_s_current_state_reg ( .D(
        new_AGEMA_signal_5911), .CK(clk), .Q(new_AGEMA_signal_5912), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3638_s_current_state_reg ( .D(
        new_AGEMA_signal_5915), .CK(clk), .Q(new_AGEMA_signal_5916), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3642_s_current_state_reg ( .D(
        new_AGEMA_signal_5919), .CK(clk), .Q(new_AGEMA_signal_5920), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3646_s_current_state_reg ( .D(
        new_AGEMA_signal_5923), .CK(clk), .Q(new_AGEMA_signal_5924), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3650_s_current_state_reg ( .D(
        new_AGEMA_signal_5927), .CK(clk), .Q(new_AGEMA_signal_5928), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3654_s_current_state_reg ( .D(
        new_AGEMA_signal_5931), .CK(clk), .Q(new_AGEMA_signal_5932), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3658_s_current_state_reg ( .D(
        new_AGEMA_signal_5935), .CK(clk), .Q(new_AGEMA_signal_5936), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3662_s_current_state_reg ( .D(
        new_AGEMA_signal_5939), .CK(clk), .Q(new_AGEMA_signal_5940), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3666_s_current_state_reg ( .D(
        new_AGEMA_signal_5943), .CK(clk), .Q(new_AGEMA_signal_5944), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3670_s_current_state_reg ( .D(
        new_AGEMA_signal_5947), .CK(clk), .Q(new_AGEMA_signal_5948), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3674_s_current_state_reg ( .D(
        new_AGEMA_signal_5951), .CK(clk), .Q(new_AGEMA_signal_5952), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3678_s_current_state_reg ( .D(
        new_AGEMA_signal_5955), .CK(clk), .Q(new_AGEMA_signal_5956), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3682_s_current_state_reg ( .D(
        new_AGEMA_signal_5959), .CK(clk), .Q(new_AGEMA_signal_5960), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3686_s_current_state_reg ( .D(
        new_AGEMA_signal_5963), .CK(clk), .Q(new_AGEMA_signal_5964), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3690_s_current_state_reg ( .D(
        new_AGEMA_signal_5967), .CK(clk), .Q(new_AGEMA_signal_5968), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3694_s_current_state_reg ( .D(
        new_AGEMA_signal_5971), .CK(clk), .Q(new_AGEMA_signal_5972), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3698_s_current_state_reg ( .D(
        new_AGEMA_signal_5975), .CK(clk), .Q(new_AGEMA_signal_5976), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3702_s_current_state_reg ( .D(
        new_AGEMA_signal_5979), .CK(clk), .Q(new_AGEMA_signal_5980), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3706_s_current_state_reg ( .D(
        new_AGEMA_signal_5983), .CK(clk), .Q(new_AGEMA_signal_5984), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3710_s_current_state_reg ( .D(
        new_AGEMA_signal_5987), .CK(clk), .Q(new_AGEMA_signal_5988), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3714_s_current_state_reg ( .D(
        new_AGEMA_signal_5991), .CK(clk), .Q(new_AGEMA_signal_5992), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3718_s_current_state_reg ( .D(
        new_AGEMA_signal_5995), .CK(clk), .Q(new_AGEMA_signal_5996), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3722_s_current_state_reg ( .D(
        new_AGEMA_signal_5999), .CK(clk), .Q(new_AGEMA_signal_6000), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3726_s_current_state_reg ( .D(
        new_AGEMA_signal_6003), .CK(clk), .Q(new_AGEMA_signal_6004), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3730_s_current_state_reg ( .D(
        new_AGEMA_signal_6007), .CK(clk), .Q(new_AGEMA_signal_6008), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3734_s_current_state_reg ( .D(
        new_AGEMA_signal_6011), .CK(clk), .Q(new_AGEMA_signal_6012), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3738_s_current_state_reg ( .D(
        new_AGEMA_signal_6015), .CK(clk), .Q(new_AGEMA_signal_6016), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3742_s_current_state_reg ( .D(
        new_AGEMA_signal_6019), .CK(clk), .Q(new_AGEMA_signal_6020), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3746_s_current_state_reg ( .D(
        new_AGEMA_signal_6023), .CK(clk), .Q(new_AGEMA_signal_6024), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3750_s_current_state_reg ( .D(
        new_AGEMA_signal_6027), .CK(clk), .Q(new_AGEMA_signal_6028), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3754_s_current_state_reg ( .D(
        new_AGEMA_signal_6031), .CK(clk), .Q(new_AGEMA_signal_6032), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3758_s_current_state_reg ( .D(
        new_AGEMA_signal_6035), .CK(clk), .Q(new_AGEMA_signal_6036), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3762_s_current_state_reg ( .D(
        new_AGEMA_signal_6039), .CK(clk), .Q(new_AGEMA_signal_6040), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3766_s_current_state_reg ( .D(
        new_AGEMA_signal_6043), .CK(clk), .Q(new_AGEMA_signal_6044), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3770_s_current_state_reg ( .D(
        new_AGEMA_signal_6047), .CK(clk), .Q(new_AGEMA_signal_6048), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3774_s_current_state_reg ( .D(
        new_AGEMA_signal_6051), .CK(clk), .Q(new_AGEMA_signal_6052), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3778_s_current_state_reg ( .D(
        new_AGEMA_signal_6055), .CK(clk), .Q(new_AGEMA_signal_6056), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3782_s_current_state_reg ( .D(
        new_AGEMA_signal_6059), .CK(clk), .Q(new_AGEMA_signal_6060), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3786_s_current_state_reg ( .D(
        new_AGEMA_signal_6063), .CK(clk), .Q(new_AGEMA_signal_6064), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3790_s_current_state_reg ( .D(
        new_AGEMA_signal_6067), .CK(clk), .Q(new_AGEMA_signal_6068), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3794_s_current_state_reg ( .D(
        new_AGEMA_signal_6071), .CK(clk), .Q(new_AGEMA_signal_6072), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3798_s_current_state_reg ( .D(
        new_AGEMA_signal_6075), .CK(clk), .Q(new_AGEMA_signal_6076), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3802_s_current_state_reg ( .D(
        new_AGEMA_signal_6079), .CK(clk), .Q(new_AGEMA_signal_6080), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3806_s_current_state_reg ( .D(
        new_AGEMA_signal_6083), .CK(clk), .Q(new_AGEMA_signal_6084), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3810_s_current_state_reg ( .D(
        new_AGEMA_signal_6087), .CK(clk), .Q(new_AGEMA_signal_6088), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3814_s_current_state_reg ( .D(
        new_AGEMA_signal_6091), .CK(clk), .Q(new_AGEMA_signal_6092), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3818_s_current_state_reg ( .D(
        new_AGEMA_signal_6095), .CK(clk), .Q(new_AGEMA_signal_6096), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3822_s_current_state_reg ( .D(
        new_AGEMA_signal_6099), .CK(clk), .Q(new_AGEMA_signal_6100), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3826_s_current_state_reg ( .D(
        new_AGEMA_signal_6103), .CK(clk), .Q(new_AGEMA_signal_6104), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3830_s_current_state_reg ( .D(
        new_AGEMA_signal_6107), .CK(clk), .Q(new_AGEMA_signal_6108), .QN() );
  MUX2_X1 PlaintextMUX_MUXInst_0_U1_Ins_0_U1 ( .A(MCOutput[0]), .B(
        new_AGEMA_signal_3961), .S(n43), .Z(StateRegInput[0]) );
  MUX2_X1 PlaintextMUX_MUXInst_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2890), .B(
        new_AGEMA_signal_3965), .S(n43), .Z(new_AGEMA_signal_2908) );
  MUX2_X1 PlaintextMUX_MUXInst_0_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2891), .B(
        new_AGEMA_signal_3969), .S(n43), .Z(new_AGEMA_signal_2909) );
  MUX2_X1 PlaintextMUX_MUXInst_1_U1_Ins_0_U1 ( .A(MCOutput[1]), .B(
        new_AGEMA_signal_3973), .S(n44), .Z(StateRegInput[1]) );
  MUX2_X1 PlaintextMUX_MUXInst_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2982), .B(
        new_AGEMA_signal_3977), .S(n44), .Z(new_AGEMA_signal_2994) );
  MUX2_X1 PlaintextMUX_MUXInst_1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2983), .B(
        new_AGEMA_signal_3981), .S(n44), .Z(new_AGEMA_signal_2995) );
  MUX2_X1 PlaintextMUX_MUXInst_4_U1_Ins_0_U1 ( .A(MCOutput[4]), .B(
        new_AGEMA_signal_3985), .S(new_AGEMA_signal_3957), .Z(StateRegInput[4]) );
  MUX2_X1 PlaintextMUX_MUXInst_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2894), .B(
        new_AGEMA_signal_3989), .S(new_AGEMA_signal_3957), .Z(
        new_AGEMA_signal_2912) );
  MUX2_X1 PlaintextMUX_MUXInst_4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2895), .B(
        new_AGEMA_signal_3993), .S(new_AGEMA_signal_3957), .Z(
        new_AGEMA_signal_2913) );
  MUX2_X1 PlaintextMUX_MUXInst_5_U1_Ins_0_U1 ( .A(MCOutput[5]), .B(
        new_AGEMA_signal_3997), .S(new_AGEMA_signal_3957), .Z(StateRegInput[5]) );
  MUX2_X1 PlaintextMUX_MUXInst_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2984), .B(
        new_AGEMA_signal_4001), .S(new_AGEMA_signal_3957), .Z(
        new_AGEMA_signal_2998) );
  MUX2_X1 PlaintextMUX_MUXInst_5_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2985), .B(
        new_AGEMA_signal_4005), .S(new_AGEMA_signal_3957), .Z(
        new_AGEMA_signal_2999) );
  MUX2_X1 PlaintextMUX_MUXInst_8_U1_Ins_0_U1 ( .A(MCOutput[8]), .B(
        new_AGEMA_signal_4009), .S(new_AGEMA_signal_3957), .Z(StateRegInput[8]) );
  MUX2_X1 PlaintextMUX_MUXInst_8_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2898), .B(
        new_AGEMA_signal_4013), .S(new_AGEMA_signal_3957), .Z(
        new_AGEMA_signal_2916) );
  MUX2_X1 PlaintextMUX_MUXInst_8_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2899), .B(
        new_AGEMA_signal_4017), .S(new_AGEMA_signal_3957), .Z(
        new_AGEMA_signal_2917) );
  MUX2_X1 PlaintextMUX_MUXInst_9_U1_Ins_0_U1 ( .A(MCOutput[9]), .B(
        new_AGEMA_signal_4021), .S(n40), .Z(StateRegInput[9]) );
  MUX2_X1 PlaintextMUX_MUXInst_9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2986), .B(
        new_AGEMA_signal_4025), .S(n40), .Z(new_AGEMA_signal_3002) );
  MUX2_X1 PlaintextMUX_MUXInst_9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2987), .B(
        new_AGEMA_signal_4029), .S(n40), .Z(new_AGEMA_signal_3003) );
  MUX2_X1 PlaintextMUX_MUXInst_12_U1_Ins_0_U1 ( .A(MCOutput[12]), .B(
        new_AGEMA_signal_4033), .S(n40), .Z(StateRegInput[12]) );
  MUX2_X1 PlaintextMUX_MUXInst_12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3052), .B(
        new_AGEMA_signal_4037), .S(n40), .Z(new_AGEMA_signal_3058) );
  MUX2_X1 PlaintextMUX_MUXInst_12_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3053), .B(
        new_AGEMA_signal_4041), .S(n40), .Z(new_AGEMA_signal_3059) );
  MUX2_X1 PlaintextMUX_MUXInst_13_U1_Ins_0_U1 ( .A(MCOutput[13]), .B(
        new_AGEMA_signal_4045), .S(n40), .Z(StateRegInput[13]) );
  MUX2_X1 PlaintextMUX_MUXInst_13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3072), .B(
        new_AGEMA_signal_4049), .S(n40), .Z(new_AGEMA_signal_3076) );
  MUX2_X1 PlaintextMUX_MUXInst_13_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3073), .B(
        new_AGEMA_signal_4053), .S(n40), .Z(new_AGEMA_signal_3077) );
  MUX2_X1 PlaintextMUX_MUXInst_16_U1_Ins_0_U1 ( .A(MCOutput[16]), .B(
        new_AGEMA_signal_4057), .S(n40), .Z(StateRegInput[16]) );
  MUX2_X1 PlaintextMUX_MUXInst_16_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2874), .B(
        new_AGEMA_signal_4061), .S(n40), .Z(new_AGEMA_signal_2924) );
  MUX2_X1 PlaintextMUX_MUXInst_16_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2875), .B(
        new_AGEMA_signal_4065), .S(n40), .Z(new_AGEMA_signal_2925) );
  MUX2_X1 PlaintextMUX_MUXInst_17_U1_Ins_0_U1 ( .A(MCOutput[17]), .B(
        new_AGEMA_signal_4069), .S(n40), .Z(StateRegInput[17]) );
  MUX2_X1 PlaintextMUX_MUXInst_17_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2972), .B(
        new_AGEMA_signal_4073), .S(n40), .Z(new_AGEMA_signal_3010) );
  MUX2_X1 PlaintextMUX_MUXInst_17_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2973), .B(
        new_AGEMA_signal_4077), .S(n40), .Z(new_AGEMA_signal_3011) );
  MUX2_X1 PlaintextMUX_MUXInst_20_U1_Ins_0_U1 ( .A(MCOutput[20]), .B(
        new_AGEMA_signal_4081), .S(n41), .Z(StateRegInput[20]) );
  MUX2_X1 PlaintextMUX_MUXInst_20_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2878), .B(
        new_AGEMA_signal_4085), .S(n41), .Z(new_AGEMA_signal_2928) );
  MUX2_X1 PlaintextMUX_MUXInst_20_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2879), .B(
        new_AGEMA_signal_4089), .S(n41), .Z(new_AGEMA_signal_2929) );
  MUX2_X1 PlaintextMUX_MUXInst_21_U1_Ins_0_U1 ( .A(MCOutput[21]), .B(
        new_AGEMA_signal_4093), .S(n41), .Z(StateRegInput[21]) );
  MUX2_X1 PlaintextMUX_MUXInst_21_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2974), .B(
        new_AGEMA_signal_4097), .S(n41), .Z(new_AGEMA_signal_3014) );
  MUX2_X1 PlaintextMUX_MUXInst_21_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2975), .B(
        new_AGEMA_signal_4101), .S(n41), .Z(new_AGEMA_signal_3015) );
  MUX2_X1 PlaintextMUX_MUXInst_24_U1_Ins_0_U1 ( .A(MCOutput[24]), .B(
        new_AGEMA_signal_4105), .S(n41), .Z(StateRegInput[24]) );
  MUX2_X1 PlaintextMUX_MUXInst_24_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3048), .B(
        new_AGEMA_signal_4109), .S(n41), .Z(new_AGEMA_signal_3062) );
  MUX2_X1 PlaintextMUX_MUXInst_24_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3049), .B(
        new_AGEMA_signal_4113), .S(n41), .Z(new_AGEMA_signal_3063) );
  MUX2_X1 PlaintextMUX_MUXInst_25_U1_Ins_0_U1 ( .A(MCOutput[25]), .B(
        new_AGEMA_signal_4117), .S(n41), .Z(StateRegInput[25]) );
  MUX2_X1 PlaintextMUX_MUXInst_25_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3070), .B(
        new_AGEMA_signal_4121), .S(n41), .Z(new_AGEMA_signal_3080) );
  MUX2_X1 PlaintextMUX_MUXInst_25_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3071), .B(
        new_AGEMA_signal_4125), .S(n41), .Z(new_AGEMA_signal_3081) );
  MUX2_X1 PlaintextMUX_MUXInst_28_U1_Ins_0_U1 ( .A(MCOutput[28]), .B(
        new_AGEMA_signal_4129), .S(n41), .Z(StateRegInput[28]) );
  MUX2_X1 PlaintextMUX_MUXInst_28_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2886), .B(
        new_AGEMA_signal_4133), .S(n41), .Z(new_AGEMA_signal_2936) );
  MUX2_X1 PlaintextMUX_MUXInst_28_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2887), .B(
        new_AGEMA_signal_4137), .S(n41), .Z(new_AGEMA_signal_2937) );
  MUX2_X1 PlaintextMUX_MUXInst_29_U1_Ins_0_U1 ( .A(MCOutput[29]), .B(
        new_AGEMA_signal_4141), .S(n42), .Z(StateRegInput[29]) );
  MUX2_X1 PlaintextMUX_MUXInst_29_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2980), .B(
        new_AGEMA_signal_4145), .S(n42), .Z(new_AGEMA_signal_3022) );
  MUX2_X1 PlaintextMUX_MUXInst_29_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2981), .B(
        new_AGEMA_signal_4149), .S(n42), .Z(new_AGEMA_signal_3023) );
  MUX2_X1 PlaintextMUX_MUXInst_32_U1_Ins_0_U1 ( .A(MCOutput[32]), .B(
        new_AGEMA_signal_4153), .S(n42), .Z(StateRegInput[32]) );
  MUX2_X1 PlaintextMUX_MUXInst_32_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2620), .B(
        new_AGEMA_signal_4157), .S(n42), .Z(new_AGEMA_signal_2704) );
  MUX2_X1 PlaintextMUX_MUXInst_32_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2621), .B(
        new_AGEMA_signal_4161), .S(n42), .Z(new_AGEMA_signal_2705) );
  MUX2_X1 PlaintextMUX_MUXInst_33_U1_Ins_0_U1 ( .A(MCOutput[33]), .B(
        new_AGEMA_signal_4165), .S(n42), .Z(StateRegInput[33]) );
  MUX2_X1 PlaintextMUX_MUXInst_33_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2744), .B(
        new_AGEMA_signal_4169), .S(n42), .Z(new_AGEMA_signal_2824) );
  MUX2_X1 PlaintextMUX_MUXInst_33_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2745), .B(
        new_AGEMA_signal_4173), .S(n42), .Z(new_AGEMA_signal_2825) );
  MUX2_X1 PlaintextMUX_MUXInst_36_U1_Ins_0_U1 ( .A(MCOutput[36]), .B(
        new_AGEMA_signal_4177), .S(n42), .Z(StateRegInput[36]) );
  MUX2_X1 PlaintextMUX_MUXInst_36_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2624), .B(
        new_AGEMA_signal_4181), .S(n42), .Z(new_AGEMA_signal_2708) );
  MUX2_X1 PlaintextMUX_MUXInst_36_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2625), .B(
        new_AGEMA_signal_4185), .S(n42), .Z(new_AGEMA_signal_2709) );
  MUX2_X1 PlaintextMUX_MUXInst_37_U1_Ins_0_U1 ( .A(MCOutput[37]), .B(
        new_AGEMA_signal_4189), .S(n42), .Z(StateRegInput[37]) );
  MUX2_X1 PlaintextMUX_MUXInst_37_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2746), .B(
        new_AGEMA_signal_4193), .S(n42), .Z(new_AGEMA_signal_2828) );
  MUX2_X1 PlaintextMUX_MUXInst_37_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2747), .B(
        new_AGEMA_signal_4197), .S(n42), .Z(new_AGEMA_signal_2829) );
  MUX2_X1 PlaintextMUX_MUXInst_40_U1_Ins_0_U1 ( .A(MCOutput[40]), .B(
        new_AGEMA_signal_4201), .S(n43), .Z(StateRegInput[40]) );
  MUX2_X1 PlaintextMUX_MUXInst_40_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2628), .B(
        new_AGEMA_signal_4205), .S(n43), .Z(new_AGEMA_signal_2712) );
  MUX2_X1 PlaintextMUX_MUXInst_40_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2629), .B(
        new_AGEMA_signal_4209), .S(n43), .Z(new_AGEMA_signal_2713) );
  MUX2_X1 PlaintextMUX_MUXInst_41_U1_Ins_0_U1 ( .A(MCOutput[41]), .B(
        new_AGEMA_signal_4213), .S(n43), .Z(StateRegInput[41]) );
  MUX2_X1 PlaintextMUX_MUXInst_41_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2748), .B(
        new_AGEMA_signal_4217), .S(n43), .Z(new_AGEMA_signal_2832) );
  MUX2_X1 PlaintextMUX_MUXInst_41_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2749), .B(
        new_AGEMA_signal_4221), .S(n43), .Z(new_AGEMA_signal_2833) );
  MUX2_X1 PlaintextMUX_MUXInst_44_U1_Ins_0_U1 ( .A(MCOutput[44]), .B(
        new_AGEMA_signal_4225), .S(n43), .Z(StateRegInput[44]) );
  MUX2_X1 PlaintextMUX_MUXInst_44_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2854), .B(
        new_AGEMA_signal_4229), .S(n43), .Z(new_AGEMA_signal_2940) );
  MUX2_X1 PlaintextMUX_MUXInst_44_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2855), .B(
        new_AGEMA_signal_4233), .S(n43), .Z(new_AGEMA_signal_2941) );
  MUX2_X1 PlaintextMUX_MUXInst_45_U1_Ins_0_U1 ( .A(MCOutput[45]), .B(
        new_AGEMA_signal_4237), .S(n43), .Z(StateRegInput[45]) );
  MUX2_X1 PlaintextMUX_MUXInst_45_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2960), .B(
        new_AGEMA_signal_4241), .S(n43), .Z(new_AGEMA_signal_3026) );
  MUX2_X1 PlaintextMUX_MUXInst_45_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2961), .B(
        new_AGEMA_signal_4245), .S(n43), .Z(new_AGEMA_signal_3027) );
  MUX2_X1 PlaintextMUX_MUXInst_48_U1_Ins_0_U1 ( .A(MCOutput[48]), .B(
        new_AGEMA_signal_4249), .S(n43), .Z(StateRegInput[48]) );
  MUX2_X1 PlaintextMUX_MUXInst_48_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2858), .B(
        new_AGEMA_signal_4253), .S(n43), .Z(new_AGEMA_signal_2944) );
  MUX2_X1 PlaintextMUX_MUXInst_48_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2859), .B(
        new_AGEMA_signal_4257), .S(n43), .Z(new_AGEMA_signal_2945) );
  MUX2_X1 PlaintextMUX_MUXInst_49_U1_Ins_0_U1 ( .A(MCOutput[49]), .B(
        new_AGEMA_signal_4261), .S(n44), .Z(StateRegInput[49]) );
  MUX2_X1 PlaintextMUX_MUXInst_49_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2962), .B(
        new_AGEMA_signal_4265), .S(n44), .Z(new_AGEMA_signal_3030) );
  MUX2_X1 PlaintextMUX_MUXInst_49_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2963), .B(
        new_AGEMA_signal_4269), .S(n44), .Z(new_AGEMA_signal_3031) );
  MUX2_X1 PlaintextMUX_MUXInst_52_U1_Ins_0_U1 ( .A(MCOutput[52]), .B(
        new_AGEMA_signal_4273), .S(n44), .Z(StateRegInput[52]) );
  MUX2_X1 PlaintextMUX_MUXInst_52_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2862), .B(
        new_AGEMA_signal_4277), .S(n44), .Z(new_AGEMA_signal_2948) );
  MUX2_X1 PlaintextMUX_MUXInst_52_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2863), .B(
        new_AGEMA_signal_4281), .S(n44), .Z(new_AGEMA_signal_2949) );
  MUX2_X1 PlaintextMUX_MUXInst_53_U1_Ins_0_U1 ( .A(MCOutput[53]), .B(
        new_AGEMA_signal_4285), .S(n44), .Z(StateRegInput[53]) );
  MUX2_X1 PlaintextMUX_MUXInst_53_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2964), .B(
        new_AGEMA_signal_4289), .S(n44), .Z(new_AGEMA_signal_3034) );
  MUX2_X1 PlaintextMUX_MUXInst_53_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2965), .B(
        new_AGEMA_signal_4293), .S(n44), .Z(new_AGEMA_signal_3035) );
  MUX2_X1 PlaintextMUX_MUXInst_56_U1_Ins_0_U1 ( .A(MCOutput[56]), .B(
        new_AGEMA_signal_4297), .S(n44), .Z(StateRegInput[56]) );
  MUX2_X1 PlaintextMUX_MUXInst_56_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2866), .B(
        new_AGEMA_signal_4301), .S(n44), .Z(new_AGEMA_signal_2952) );
  MUX2_X1 PlaintextMUX_MUXInst_56_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2867), .B(
        new_AGEMA_signal_4305), .S(n44), .Z(new_AGEMA_signal_2953) );
  MUX2_X1 PlaintextMUX_MUXInst_57_U1_Ins_0_U1 ( .A(MCOutput[57]), .B(
        new_AGEMA_signal_4309), .S(n44), .Z(StateRegInput[57]) );
  MUX2_X1 PlaintextMUX_MUXInst_57_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2966), .B(
        new_AGEMA_signal_4313), .S(n44), .Z(new_AGEMA_signal_3038) );
  MUX2_X1 PlaintextMUX_MUXInst_57_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2967), .B(
        new_AGEMA_signal_4317), .S(n44), .Z(new_AGEMA_signal_3039) );
  MUX2_X1 PlaintextMUX_MUXInst_60_U1_Ins_0_U1 ( .A(MCOutput[60]), .B(
        new_AGEMA_signal_4321), .S(new_AGEMA_signal_3957), .Z(
        StateRegInput[60]) );
  MUX2_X1 PlaintextMUX_MUXInst_60_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3044), .B(
        new_AGEMA_signal_4325), .S(new_AGEMA_signal_3957), .Z(
        new_AGEMA_signal_3066) );
  MUX2_X1 PlaintextMUX_MUXInst_60_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3045), .B(
        new_AGEMA_signal_4329), .S(new_AGEMA_signal_3957), .Z(
        new_AGEMA_signal_3067) );
  MUX2_X1 PlaintextMUX_MUXInst_61_U1_Ins_0_U1 ( .A(MCOutput[61]), .B(
        new_AGEMA_signal_4333), .S(new_AGEMA_signal_3957), .Z(
        StateRegInput[61]) );
  MUX2_X1 PlaintextMUX_MUXInst_61_U1_Ins_1_U1 ( .A(new_AGEMA_signal_3068), .B(
        new_AGEMA_signal_4337), .S(new_AGEMA_signal_3957), .Z(
        new_AGEMA_signal_3084) );
  MUX2_X1 PlaintextMUX_MUXInst_61_U1_Ins_2_U1 ( .A(new_AGEMA_signal_3069), .B(
        new_AGEMA_signal_4341), .S(new_AGEMA_signal_3957), .Z(
        new_AGEMA_signal_3085) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U37 ( .A(new_AGEMA_signal_2028), .B(
        Fresh[98]), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U36 ( .A(Fresh[97]), .B(
        SubCellInst_SboxInst_0_Q2), .Z(
        SubCellInst_SboxInst_0_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U35 ( .A(new_AGEMA_signal_2029), .B(
        Fresh[98]), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U34 ( .A(Fresh[96]), .B(
        SubCellInst_SboxInst_0_Q2), .Z(
        SubCellInst_SboxInst_0_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U33 ( .A(Fresh[97]), .B(
        new_AGEMA_signal_2029), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U32 ( .A(new_AGEMA_signal_2028), .B(
        Fresh[96]), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U25 ( .A1(new_AGEMA_signal_4347), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U24 ( .A1(new_AGEMA_signal_4347), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U23 ( .A1(new_AGEMA_signal_4345), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND2_U1_U22 ( .A(Fresh[98]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U21 ( .A1(new_AGEMA_signal_4345), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U20 ( .A1(new_AGEMA_signal_4343), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND2_U1_U19 ( .A(Fresh[97]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U18 ( .A1(new_AGEMA_signal_4343), 
        .A2(SubCellInst_SboxInst_0_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND2_U1_U17 ( .A(Fresh[96]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U16 ( .A1(new_AGEMA_signal_2029), 
        .A2(new_AGEMA_signal_4347), .ZN(SubCellInst_SboxInst_0_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U15 ( .A1(new_AGEMA_signal_2028), 
        .A2(new_AGEMA_signal_4345), .ZN(SubCellInst_SboxInst_0_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_0_Q2), 
        .A2(new_AGEMA_signal_4343), .ZN(SubCellInst_SboxInst_0_AND2_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND2_U1_n33), .Z(new_AGEMA_signal_2159) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n32), .B(
        SubCellInst_SboxInst_0_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_0_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND2_U1_n30), .Z(new_AGEMA_signal_2158) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n29), .B(
        SubCellInst_SboxInst_0_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_0_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND2_U1_n27), .Z(SubCellInst_SboxInst_0_T1) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n26), .B(
        SubCellInst_SboxInst_0_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_0_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4343), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4345), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4347), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_T1), .B(new_AGEMA_signal_4349), .Z(
        SubCellInst_SboxInst_0_L0) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2158), 
        .B(new_AGEMA_signal_4351), .Z(new_AGEMA_signal_2286) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2159), 
        .B(new_AGEMA_signal_4353), .Z(new_AGEMA_signal_2287) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U37 ( .A(new_AGEMA_signal_2030), .B(
        Fresh[101]), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U36 ( .A(Fresh[100]), .B(
        SubCellInst_SboxInst_0_Q7), .Z(
        SubCellInst_SboxInst_0_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U35 ( .A(new_AGEMA_signal_2031), .B(
        Fresh[101]), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U34 ( .A(Fresh[99]), .B(
        SubCellInst_SboxInst_0_Q7), .Z(
        SubCellInst_SboxInst_0_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U33 ( .A(Fresh[100]), .B(
        new_AGEMA_signal_2031), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U32 ( .A(new_AGEMA_signal_2030), .B(
        Fresh[99]), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U25 ( .A1(new_AGEMA_signal_4359), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U24 ( .A1(new_AGEMA_signal_4359), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U23 ( .A1(new_AGEMA_signal_4357), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND4_U1_U22 ( .A(Fresh[101]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U21 ( .A1(new_AGEMA_signal_4357), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U20 ( .A1(new_AGEMA_signal_4355), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_0_AND4_U1_U19 ( .A(Fresh[100]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U18 ( .A1(new_AGEMA_signal_4355), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND4_U1_U17 ( .A(Fresh[99]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U16 ( .A1(new_AGEMA_signal_2031), 
        .A2(new_AGEMA_signal_4359), .ZN(SubCellInst_SboxInst_0_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U15 ( .A1(new_AGEMA_signal_2030), 
        .A2(new_AGEMA_signal_4357), .ZN(SubCellInst_SboxInst_0_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_0_Q7), 
        .A2(new_AGEMA_signal_4355), .ZN(SubCellInst_SboxInst_0_AND4_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND4_U1_n33), .Z(new_AGEMA_signal_2161) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n32), .B(
        SubCellInst_SboxInst_0_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_0_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_0_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND4_U1_n30), .Z(new_AGEMA_signal_2160) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n29), .B(
        SubCellInst_SboxInst_0_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_0_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND4_U1_n27), .Z(SubCellInst_SboxInst_0_T3) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n26), .B(
        SubCellInst_SboxInst_0_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_0_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4355), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4357), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4359), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L0), .B(new_AGEMA_signal_4363), .Z(
        SubCellInst_SboxInst_0_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2286), 
        .B(new_AGEMA_signal_4367), .Z(new_AGEMA_signal_2372) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2287), 
        .B(new_AGEMA_signal_4371), .Z(new_AGEMA_signal_2373) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L0), .B(SubCellInst_SboxInst_0_T3), .Z(
        ShiftRowsOutput[4]) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2286), 
        .B(new_AGEMA_signal_2160), .Z(new_AGEMA_signal_2374) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2287), 
        .B(new_AGEMA_signal_2161), .Z(new_AGEMA_signal_2375) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_4373), .B(SubCellInst_SboxInst_0_YY_3), .ZN(ShiftRowsOutput[5]) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4375), .B(new_AGEMA_signal_2372), .Z(new_AGEMA_signal_2488) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4377), .B(new_AGEMA_signal_2373), .Z(new_AGEMA_signal_2489) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U37 ( .A(new_AGEMA_signal_2036), .B(
        Fresh[104]), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U36 ( .A(Fresh[103]), .B(
        SubCellInst_SboxInst_1_Q2), .Z(
        SubCellInst_SboxInst_1_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U35 ( .A(new_AGEMA_signal_2037), .B(
        Fresh[104]), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U34 ( .A(Fresh[102]), .B(
        SubCellInst_SboxInst_1_Q2), .Z(
        SubCellInst_SboxInst_1_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U33 ( .A(Fresh[103]), .B(
        new_AGEMA_signal_2037), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U32 ( .A(new_AGEMA_signal_2036), .B(
        Fresh[102]), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U25 ( .A1(new_AGEMA_signal_4383), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U24 ( .A1(new_AGEMA_signal_4383), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U23 ( .A1(new_AGEMA_signal_4381), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND2_U1_U22 ( .A(Fresh[104]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U21 ( .A1(new_AGEMA_signal_4381), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U20 ( .A1(new_AGEMA_signal_4379), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND2_U1_U19 ( .A(Fresh[103]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U18 ( .A1(new_AGEMA_signal_4379), 
        .A2(SubCellInst_SboxInst_1_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND2_U1_U17 ( .A(Fresh[102]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U16 ( .A1(new_AGEMA_signal_2037), 
        .A2(new_AGEMA_signal_4383), .ZN(SubCellInst_SboxInst_1_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U15 ( .A1(new_AGEMA_signal_2036), 
        .A2(new_AGEMA_signal_4381), .ZN(SubCellInst_SboxInst_1_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_1_Q2), 
        .A2(new_AGEMA_signal_4379), .ZN(SubCellInst_SboxInst_1_AND2_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND2_U1_n33), .Z(new_AGEMA_signal_2167) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n32), .B(
        SubCellInst_SboxInst_1_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_1_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND2_U1_n30), .Z(new_AGEMA_signal_2166) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n29), .B(
        SubCellInst_SboxInst_1_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_1_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND2_U1_n27), .Z(SubCellInst_SboxInst_1_T1) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n26), .B(
        SubCellInst_SboxInst_1_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_1_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4379), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4381), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4383), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_T1), .B(new_AGEMA_signal_4385), .Z(
        SubCellInst_SboxInst_1_L0) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2166), 
        .B(new_AGEMA_signal_4387), .Z(new_AGEMA_signal_2290) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2167), 
        .B(new_AGEMA_signal_4389), .Z(new_AGEMA_signal_2291) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U37 ( .A(new_AGEMA_signal_2038), .B(
        Fresh[107]), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U36 ( .A(Fresh[106]), .B(
        SubCellInst_SboxInst_1_Q7), .Z(
        SubCellInst_SboxInst_1_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U35 ( .A(new_AGEMA_signal_2039), .B(
        Fresh[107]), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U34 ( .A(Fresh[105]), .B(
        SubCellInst_SboxInst_1_Q7), .Z(
        SubCellInst_SboxInst_1_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U33 ( .A(Fresh[106]), .B(
        new_AGEMA_signal_2039), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U32 ( .A(new_AGEMA_signal_2038), .B(
        Fresh[105]), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U25 ( .A1(new_AGEMA_signal_4395), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U24 ( .A1(new_AGEMA_signal_4395), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U23 ( .A1(new_AGEMA_signal_4393), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND4_U1_U22 ( .A(Fresh[107]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U21 ( .A1(new_AGEMA_signal_4393), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U20 ( .A1(new_AGEMA_signal_4391), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_1_AND4_U1_U19 ( .A(Fresh[106]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U18 ( .A1(new_AGEMA_signal_4391), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND4_U1_U17 ( .A(Fresh[105]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U16 ( .A1(new_AGEMA_signal_2039), 
        .A2(new_AGEMA_signal_4395), .ZN(SubCellInst_SboxInst_1_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U15 ( .A1(new_AGEMA_signal_2038), 
        .A2(new_AGEMA_signal_4393), .ZN(SubCellInst_SboxInst_1_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_1_Q7), 
        .A2(new_AGEMA_signal_4391), .ZN(SubCellInst_SboxInst_1_AND4_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND4_U1_n33), .Z(new_AGEMA_signal_2169) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n32), .B(
        SubCellInst_SboxInst_1_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_1_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_1_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND4_U1_n30), .Z(new_AGEMA_signal_2168) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n29), .B(
        SubCellInst_SboxInst_1_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_1_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND4_U1_n27), .Z(SubCellInst_SboxInst_1_T3) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n26), .B(
        SubCellInst_SboxInst_1_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_1_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4391), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4393), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4395), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L0), .B(new_AGEMA_signal_4399), .Z(
        SubCellInst_SboxInst_1_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2290), 
        .B(new_AGEMA_signal_4403), .Z(new_AGEMA_signal_2376) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2291), 
        .B(new_AGEMA_signal_4407), .Z(new_AGEMA_signal_2377) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L0), .B(SubCellInst_SboxInst_1_T3), .Z(
        ShiftRowsOutput[8]) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2290), 
        .B(new_AGEMA_signal_2168), .Z(new_AGEMA_signal_2378) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2291), 
        .B(new_AGEMA_signal_2169), .Z(new_AGEMA_signal_2379) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_4409), .B(SubCellInst_SboxInst_1_YY_3), .ZN(ShiftRowsOutput[9]) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4411), .B(new_AGEMA_signal_2376), .Z(new_AGEMA_signal_2490) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4413), .B(new_AGEMA_signal_2377), .Z(new_AGEMA_signal_2491) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U37 ( .A(new_AGEMA_signal_2044), .B(
        Fresh[110]), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U36 ( .A(Fresh[109]), .B(
        SubCellInst_SboxInst_2_Q2), .Z(
        SubCellInst_SboxInst_2_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U35 ( .A(new_AGEMA_signal_2045), .B(
        Fresh[110]), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U34 ( .A(Fresh[108]), .B(
        SubCellInst_SboxInst_2_Q2), .Z(
        SubCellInst_SboxInst_2_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U33 ( .A(Fresh[109]), .B(
        new_AGEMA_signal_2045), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U32 ( .A(new_AGEMA_signal_2044), .B(
        Fresh[108]), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U25 ( .A1(new_AGEMA_signal_4419), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U24 ( .A1(new_AGEMA_signal_4419), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U23 ( .A1(new_AGEMA_signal_4417), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND2_U1_U22 ( .A(Fresh[110]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U21 ( .A1(new_AGEMA_signal_4417), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U20 ( .A1(new_AGEMA_signal_4415), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND2_U1_U19 ( .A(Fresh[109]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U18 ( .A1(new_AGEMA_signal_4415), 
        .A2(SubCellInst_SboxInst_2_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND2_U1_U17 ( .A(Fresh[108]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U16 ( .A1(new_AGEMA_signal_2045), 
        .A2(new_AGEMA_signal_4419), .ZN(SubCellInst_SboxInst_2_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U15 ( .A1(new_AGEMA_signal_2044), 
        .A2(new_AGEMA_signal_4417), .ZN(SubCellInst_SboxInst_2_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_2_Q2), 
        .A2(new_AGEMA_signal_4415), .ZN(SubCellInst_SboxInst_2_AND2_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND2_U1_n33), .Z(new_AGEMA_signal_2175) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n32), .B(
        SubCellInst_SboxInst_2_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_2_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND2_U1_n30), .Z(new_AGEMA_signal_2174) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n29), .B(
        SubCellInst_SboxInst_2_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_2_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND2_U1_n27), .Z(SubCellInst_SboxInst_2_T1) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n26), .B(
        SubCellInst_SboxInst_2_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_2_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4415), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4417), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4419), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_T1), .B(new_AGEMA_signal_4421), .Z(
        SubCellInst_SboxInst_2_L0) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2174), 
        .B(new_AGEMA_signal_4423), .Z(new_AGEMA_signal_2294) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2175), 
        .B(new_AGEMA_signal_4425), .Z(new_AGEMA_signal_2295) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U37 ( .A(new_AGEMA_signal_2046), .B(
        Fresh[113]), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U36 ( .A(Fresh[112]), .B(
        SubCellInst_SboxInst_2_Q7), .Z(
        SubCellInst_SboxInst_2_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U35 ( .A(new_AGEMA_signal_2047), .B(
        Fresh[113]), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U34 ( .A(Fresh[111]), .B(
        SubCellInst_SboxInst_2_Q7), .Z(
        SubCellInst_SboxInst_2_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U33 ( .A(Fresh[112]), .B(
        new_AGEMA_signal_2047), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U32 ( .A(new_AGEMA_signal_2046), .B(
        Fresh[111]), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U25 ( .A1(new_AGEMA_signal_4431), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U24 ( .A1(new_AGEMA_signal_4431), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U23 ( .A1(new_AGEMA_signal_4429), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND4_U1_U22 ( .A(Fresh[113]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U21 ( .A1(new_AGEMA_signal_4429), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U20 ( .A1(new_AGEMA_signal_4427), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_2_AND4_U1_U19 ( .A(Fresh[112]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U18 ( .A1(new_AGEMA_signal_4427), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND4_U1_U17 ( .A(Fresh[111]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U16 ( .A1(new_AGEMA_signal_2047), 
        .A2(new_AGEMA_signal_4431), .ZN(SubCellInst_SboxInst_2_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U15 ( .A1(new_AGEMA_signal_2046), 
        .A2(new_AGEMA_signal_4429), .ZN(SubCellInst_SboxInst_2_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_2_Q7), 
        .A2(new_AGEMA_signal_4427), .ZN(SubCellInst_SboxInst_2_AND4_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND4_U1_n33), .Z(new_AGEMA_signal_2177) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n32), .B(
        SubCellInst_SboxInst_2_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_2_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_2_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND4_U1_n30), .Z(new_AGEMA_signal_2176) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n29), .B(
        SubCellInst_SboxInst_2_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_2_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND4_U1_n27), .Z(SubCellInst_SboxInst_2_T3) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n26), .B(
        SubCellInst_SboxInst_2_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_2_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4427), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4429), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4431), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L0), .B(new_AGEMA_signal_4435), .Z(
        SubCellInst_SboxInst_2_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2294), 
        .B(new_AGEMA_signal_4439), .Z(new_AGEMA_signal_2380) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2295), 
        .B(new_AGEMA_signal_4443), .Z(new_AGEMA_signal_2381) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L0), .B(SubCellInst_SboxInst_2_T3), .Z(
        ShiftRowsOutput[12]) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2294), 
        .B(new_AGEMA_signal_2176), .Z(new_AGEMA_signal_2382) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2295), 
        .B(new_AGEMA_signal_2177), .Z(new_AGEMA_signal_2383) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_4445), .B(SubCellInst_SboxInst_2_YY_3), .ZN(ShiftRowsOutput[13]) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4447), .B(new_AGEMA_signal_2380), .Z(new_AGEMA_signal_2492) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4449), .B(new_AGEMA_signal_2381), .Z(new_AGEMA_signal_2493) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U37 ( .A(new_AGEMA_signal_2052), .B(
        Fresh[116]), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U36 ( .A(Fresh[115]), .B(
        SubCellInst_SboxInst_3_Q2), .Z(
        SubCellInst_SboxInst_3_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U35 ( .A(new_AGEMA_signal_2053), .B(
        Fresh[116]), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U34 ( .A(Fresh[114]), .B(
        SubCellInst_SboxInst_3_Q2), .Z(
        SubCellInst_SboxInst_3_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U33 ( .A(Fresh[115]), .B(
        new_AGEMA_signal_2053), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U32 ( .A(new_AGEMA_signal_2052), .B(
        Fresh[114]), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U25 ( .A1(new_AGEMA_signal_4455), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U24 ( .A1(new_AGEMA_signal_4455), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U23 ( .A1(new_AGEMA_signal_4453), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND2_U1_U22 ( .A(Fresh[116]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U21 ( .A1(new_AGEMA_signal_4453), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U20 ( .A1(new_AGEMA_signal_4451), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND2_U1_U19 ( .A(Fresh[115]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U18 ( .A1(new_AGEMA_signal_4451), 
        .A2(SubCellInst_SboxInst_3_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND2_U1_U17 ( .A(Fresh[114]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U16 ( .A1(new_AGEMA_signal_2053), 
        .A2(new_AGEMA_signal_4455), .ZN(SubCellInst_SboxInst_3_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U15 ( .A1(new_AGEMA_signal_2052), 
        .A2(new_AGEMA_signal_4453), .ZN(SubCellInst_SboxInst_3_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_3_Q2), 
        .A2(new_AGEMA_signal_4451), .ZN(SubCellInst_SboxInst_3_AND2_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND2_U1_n33), .Z(new_AGEMA_signal_2183) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n32), .B(
        SubCellInst_SboxInst_3_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_3_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND2_U1_n30), .Z(new_AGEMA_signal_2182) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n29), .B(
        SubCellInst_SboxInst_3_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_3_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND2_U1_n27), .Z(SubCellInst_SboxInst_3_T1) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n26), .B(
        SubCellInst_SboxInst_3_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_3_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4451), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4453), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4455), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_T1), .B(new_AGEMA_signal_4457), .Z(
        SubCellInst_SboxInst_3_L0) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2182), 
        .B(new_AGEMA_signal_4459), .Z(new_AGEMA_signal_2298) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2183), 
        .B(new_AGEMA_signal_4461), .Z(new_AGEMA_signal_2299) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U37 ( .A(new_AGEMA_signal_2054), .B(
        Fresh[119]), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U36 ( .A(Fresh[118]), .B(
        SubCellInst_SboxInst_3_Q7), .Z(
        SubCellInst_SboxInst_3_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U35 ( .A(new_AGEMA_signal_2055), .B(
        Fresh[119]), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U34 ( .A(Fresh[117]), .B(
        SubCellInst_SboxInst_3_Q7), .Z(
        SubCellInst_SboxInst_3_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U33 ( .A(Fresh[118]), .B(
        new_AGEMA_signal_2055), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U32 ( .A(new_AGEMA_signal_2054), .B(
        Fresh[117]), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U25 ( .A1(new_AGEMA_signal_4467), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U24 ( .A1(new_AGEMA_signal_4467), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U23 ( .A1(new_AGEMA_signal_4465), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND4_U1_U22 ( .A(Fresh[119]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U21 ( .A1(new_AGEMA_signal_4465), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U20 ( .A1(new_AGEMA_signal_4463), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_3_AND4_U1_U19 ( .A(Fresh[118]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U18 ( .A1(new_AGEMA_signal_4463), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND4_U1_U17 ( .A(Fresh[117]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U16 ( .A1(new_AGEMA_signal_2055), 
        .A2(new_AGEMA_signal_4467), .ZN(SubCellInst_SboxInst_3_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U15 ( .A1(new_AGEMA_signal_2054), 
        .A2(new_AGEMA_signal_4465), .ZN(SubCellInst_SboxInst_3_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_3_Q7), 
        .A2(new_AGEMA_signal_4463), .ZN(SubCellInst_SboxInst_3_AND4_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND4_U1_n33), .Z(new_AGEMA_signal_2185) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n32), .B(
        SubCellInst_SboxInst_3_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_3_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_3_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND4_U1_n30), .Z(new_AGEMA_signal_2184) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n29), .B(
        SubCellInst_SboxInst_3_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_3_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND4_U1_n27), .Z(SubCellInst_SboxInst_3_T3) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n26), .B(
        SubCellInst_SboxInst_3_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_3_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4463), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4465), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4467), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L0), .B(new_AGEMA_signal_4471), .Z(
        SubCellInst_SboxInst_3_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2298), 
        .B(new_AGEMA_signal_4475), .Z(new_AGEMA_signal_2384) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2299), 
        .B(new_AGEMA_signal_4479), .Z(new_AGEMA_signal_2385) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L0), .B(SubCellInst_SboxInst_3_T3), .Z(
        ShiftRowsOutput[0]) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2298), 
        .B(new_AGEMA_signal_2184), .Z(new_AGEMA_signal_2386) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2299), 
        .B(new_AGEMA_signal_2185), .Z(new_AGEMA_signal_2387) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_4481), .B(SubCellInst_SboxInst_3_YY_3), .ZN(ShiftRowsOutput[1]) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4483), .B(new_AGEMA_signal_2384), .Z(new_AGEMA_signal_2494) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4485), .B(new_AGEMA_signal_2385), .Z(new_AGEMA_signal_2495) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U37 ( .A(new_AGEMA_signal_2060), .B(
        Fresh[122]), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U36 ( .A(Fresh[121]), .B(
        SubCellInst_SboxInst_4_Q2), .Z(
        SubCellInst_SboxInst_4_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U35 ( .A(new_AGEMA_signal_2061), .B(
        Fresh[122]), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U34 ( .A(Fresh[120]), .B(
        SubCellInst_SboxInst_4_Q2), .Z(
        SubCellInst_SboxInst_4_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U33 ( .A(Fresh[121]), .B(
        new_AGEMA_signal_2061), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U32 ( .A(new_AGEMA_signal_2060), .B(
        Fresh[120]), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U25 ( .A1(new_AGEMA_signal_4491), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U24 ( .A1(new_AGEMA_signal_4491), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U23 ( .A1(new_AGEMA_signal_4489), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND2_U1_U22 ( .A(Fresh[122]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U21 ( .A1(new_AGEMA_signal_4489), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U20 ( .A1(new_AGEMA_signal_4487), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND2_U1_U19 ( .A(Fresh[121]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U18 ( .A1(new_AGEMA_signal_4487), 
        .A2(SubCellInst_SboxInst_4_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND2_U1_U17 ( .A(Fresh[120]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U16 ( .A1(new_AGEMA_signal_2061), 
        .A2(new_AGEMA_signal_4491), .ZN(SubCellInst_SboxInst_4_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U15 ( .A1(new_AGEMA_signal_2060), 
        .A2(new_AGEMA_signal_4489), .ZN(SubCellInst_SboxInst_4_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_4_Q2), 
        .A2(new_AGEMA_signal_4487), .ZN(SubCellInst_SboxInst_4_AND2_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND2_U1_n33), .Z(new_AGEMA_signal_2191) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n32), .B(
        SubCellInst_SboxInst_4_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_4_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND2_U1_n30), .Z(new_AGEMA_signal_2190) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n29), .B(
        SubCellInst_SboxInst_4_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_4_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND2_U1_n27), .Z(SubCellInst_SboxInst_4_T1) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n26), .B(
        SubCellInst_SboxInst_4_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_4_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4487), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4489), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4491), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_T1), .B(new_AGEMA_signal_4493), .Z(
        SubCellInst_SboxInst_4_L0) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2190), 
        .B(new_AGEMA_signal_4495), .Z(new_AGEMA_signal_2302) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2191), 
        .B(new_AGEMA_signal_4497), .Z(new_AGEMA_signal_2303) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U37 ( .A(new_AGEMA_signal_2062), .B(
        Fresh[125]), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U36 ( .A(Fresh[124]), .B(
        SubCellInst_SboxInst_4_Q7), .Z(
        SubCellInst_SboxInst_4_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U35 ( .A(new_AGEMA_signal_2063), .B(
        Fresh[125]), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U34 ( .A(Fresh[123]), .B(
        SubCellInst_SboxInst_4_Q7), .Z(
        SubCellInst_SboxInst_4_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U33 ( .A(Fresh[124]), .B(
        new_AGEMA_signal_2063), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U32 ( .A(new_AGEMA_signal_2062), .B(
        Fresh[123]), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U25 ( .A1(new_AGEMA_signal_4503), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U24 ( .A1(new_AGEMA_signal_4503), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U23 ( .A1(new_AGEMA_signal_4501), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND4_U1_U22 ( .A(Fresh[125]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U21 ( .A1(new_AGEMA_signal_4501), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U20 ( .A1(new_AGEMA_signal_4499), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_4_AND4_U1_U19 ( .A(Fresh[124]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U18 ( .A1(new_AGEMA_signal_4499), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND4_U1_U17 ( .A(Fresh[123]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U16 ( .A1(new_AGEMA_signal_2063), 
        .A2(new_AGEMA_signal_4503), .ZN(SubCellInst_SboxInst_4_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U15 ( .A1(new_AGEMA_signal_2062), 
        .A2(new_AGEMA_signal_4501), .ZN(SubCellInst_SboxInst_4_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_4_Q7), 
        .A2(new_AGEMA_signal_4499), .ZN(SubCellInst_SboxInst_4_AND4_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND4_U1_n33), .Z(new_AGEMA_signal_2193) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n32), .B(
        SubCellInst_SboxInst_4_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_4_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_4_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND4_U1_n30), .Z(new_AGEMA_signal_2192) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n29), .B(
        SubCellInst_SboxInst_4_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_4_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND4_U1_n27), .Z(SubCellInst_SboxInst_4_T3) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n26), .B(
        SubCellInst_SboxInst_4_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_4_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4499), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4501), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4503), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L0), .B(new_AGEMA_signal_4507), .Z(
        SubCellInst_SboxInst_4_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2302), 
        .B(new_AGEMA_signal_4511), .Z(new_AGEMA_signal_2388) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2303), 
        .B(new_AGEMA_signal_4515), .Z(new_AGEMA_signal_2389) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L0), .B(SubCellInst_SboxInst_4_T3), .Z(
        ShiftRowsOutput[24]) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2302), 
        .B(new_AGEMA_signal_2192), .Z(new_AGEMA_signal_2390) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2303), 
        .B(new_AGEMA_signal_2193), .Z(new_AGEMA_signal_2391) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_4517), .B(SubCellInst_SboxInst_4_YY_3), .ZN(ShiftRowsOutput[25]) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4519), .B(new_AGEMA_signal_2388), .Z(new_AGEMA_signal_2496) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4521), .B(new_AGEMA_signal_2389), .Z(new_AGEMA_signal_2497) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U37 ( .A(new_AGEMA_signal_2068), .B(
        Fresh[128]), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U36 ( .A(Fresh[127]), .B(
        SubCellInst_SboxInst_5_Q2), .Z(
        SubCellInst_SboxInst_5_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U35 ( .A(new_AGEMA_signal_2069), .B(
        Fresh[128]), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U34 ( .A(Fresh[126]), .B(
        SubCellInst_SboxInst_5_Q2), .Z(
        SubCellInst_SboxInst_5_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U33 ( .A(Fresh[127]), .B(
        new_AGEMA_signal_2069), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U32 ( .A(new_AGEMA_signal_2068), .B(
        Fresh[126]), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U25 ( .A1(new_AGEMA_signal_4527), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U24 ( .A1(new_AGEMA_signal_4527), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U23 ( .A1(new_AGEMA_signal_4525), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND2_U1_U22 ( .A(Fresh[128]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U21 ( .A1(new_AGEMA_signal_4525), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U20 ( .A1(new_AGEMA_signal_4523), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND2_U1_U19 ( .A(Fresh[127]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U18 ( .A1(new_AGEMA_signal_4523), 
        .A2(SubCellInst_SboxInst_5_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND2_U1_U17 ( .A(Fresh[126]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U16 ( .A1(new_AGEMA_signal_2069), 
        .A2(new_AGEMA_signal_4527), .ZN(SubCellInst_SboxInst_5_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U15 ( .A1(new_AGEMA_signal_2068), 
        .A2(new_AGEMA_signal_4525), .ZN(SubCellInst_SboxInst_5_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_5_Q2), 
        .A2(new_AGEMA_signal_4523), .ZN(SubCellInst_SboxInst_5_AND2_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND2_U1_n33), .Z(new_AGEMA_signal_2199) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n32), .B(
        SubCellInst_SboxInst_5_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_5_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND2_U1_n30), .Z(new_AGEMA_signal_2198) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n29), .B(
        SubCellInst_SboxInst_5_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_5_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND2_U1_n27), .Z(SubCellInst_SboxInst_5_T1) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n26), .B(
        SubCellInst_SboxInst_5_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_5_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4523), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4525), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4527), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_T1), .B(new_AGEMA_signal_4529), .Z(
        SubCellInst_SboxInst_5_L0) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2198), 
        .B(new_AGEMA_signal_4531), .Z(new_AGEMA_signal_2306) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2199), 
        .B(new_AGEMA_signal_4533), .Z(new_AGEMA_signal_2307) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U37 ( .A(new_AGEMA_signal_2070), .B(
        Fresh[131]), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U36 ( .A(Fresh[130]), .B(
        SubCellInst_SboxInst_5_Q7), .Z(
        SubCellInst_SboxInst_5_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U35 ( .A(new_AGEMA_signal_2071), .B(
        Fresh[131]), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U34 ( .A(Fresh[129]), .B(
        SubCellInst_SboxInst_5_Q7), .Z(
        SubCellInst_SboxInst_5_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U33 ( .A(Fresh[130]), .B(
        new_AGEMA_signal_2071), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U32 ( .A(new_AGEMA_signal_2070), .B(
        Fresh[129]), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U25 ( .A1(new_AGEMA_signal_4539), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U24 ( .A1(new_AGEMA_signal_4539), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U23 ( .A1(new_AGEMA_signal_4537), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND4_U1_U22 ( .A(Fresh[131]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U21 ( .A1(new_AGEMA_signal_4537), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U20 ( .A1(new_AGEMA_signal_4535), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_5_AND4_U1_U19 ( .A(Fresh[130]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U18 ( .A1(new_AGEMA_signal_4535), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND4_U1_U17 ( .A(Fresh[129]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U16 ( .A1(new_AGEMA_signal_2071), 
        .A2(new_AGEMA_signal_4539), .ZN(SubCellInst_SboxInst_5_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U15 ( .A1(new_AGEMA_signal_2070), 
        .A2(new_AGEMA_signal_4537), .ZN(SubCellInst_SboxInst_5_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_5_Q7), 
        .A2(new_AGEMA_signal_4535), .ZN(SubCellInst_SboxInst_5_AND4_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND4_U1_n33), .Z(new_AGEMA_signal_2201) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n32), .B(
        SubCellInst_SboxInst_5_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_5_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_5_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND4_U1_n30), .Z(new_AGEMA_signal_2200) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n29), .B(
        SubCellInst_SboxInst_5_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_5_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND4_U1_n27), .Z(SubCellInst_SboxInst_5_T3) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n26), .B(
        SubCellInst_SboxInst_5_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_5_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4535), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4537), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4539), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L0), .B(new_AGEMA_signal_4543), .Z(
        SubCellInst_SboxInst_5_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2306), 
        .B(new_AGEMA_signal_4547), .Z(new_AGEMA_signal_2392) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2307), 
        .B(new_AGEMA_signal_4551), .Z(new_AGEMA_signal_2393) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L0), .B(SubCellInst_SboxInst_5_T3), .Z(
        ShiftRowsOutput[28]) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2306), 
        .B(new_AGEMA_signal_2200), .Z(new_AGEMA_signal_2394) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2307), 
        .B(new_AGEMA_signal_2201), .Z(new_AGEMA_signal_2395) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_4553), .B(SubCellInst_SboxInst_5_YY_3), .ZN(ShiftRowsOutput[29]) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4555), .B(new_AGEMA_signal_2392), .Z(new_AGEMA_signal_2498) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4557), .B(new_AGEMA_signal_2393), .Z(new_AGEMA_signal_2499) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U37 ( .A(new_AGEMA_signal_2076), .B(
        Fresh[134]), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U36 ( .A(Fresh[133]), .B(
        SubCellInst_SboxInst_6_Q2), .Z(
        SubCellInst_SboxInst_6_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U35 ( .A(new_AGEMA_signal_2077), .B(
        Fresh[134]), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U34 ( .A(Fresh[132]), .B(
        SubCellInst_SboxInst_6_Q2), .Z(
        SubCellInst_SboxInst_6_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U33 ( .A(Fresh[133]), .B(
        new_AGEMA_signal_2077), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U32 ( .A(new_AGEMA_signal_2076), .B(
        Fresh[132]), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U25 ( .A1(new_AGEMA_signal_4563), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U24 ( .A1(new_AGEMA_signal_4563), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U23 ( .A1(new_AGEMA_signal_4561), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND2_U1_U22 ( .A(Fresh[134]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U21 ( .A1(new_AGEMA_signal_4561), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U20 ( .A1(new_AGEMA_signal_4559), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND2_U1_U19 ( .A(Fresh[133]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U18 ( .A1(new_AGEMA_signal_4559), 
        .A2(SubCellInst_SboxInst_6_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND2_U1_U17 ( .A(Fresh[132]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U16 ( .A1(new_AGEMA_signal_2077), 
        .A2(new_AGEMA_signal_4563), .ZN(SubCellInst_SboxInst_6_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U15 ( .A1(new_AGEMA_signal_2076), 
        .A2(new_AGEMA_signal_4561), .ZN(SubCellInst_SboxInst_6_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_6_Q2), 
        .A2(new_AGEMA_signal_4559), .ZN(SubCellInst_SboxInst_6_AND2_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND2_U1_n33), .Z(new_AGEMA_signal_2207) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n32), .B(
        SubCellInst_SboxInst_6_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_6_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND2_U1_n30), .Z(new_AGEMA_signal_2206) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n29), .B(
        SubCellInst_SboxInst_6_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_6_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND2_U1_n27), .Z(SubCellInst_SboxInst_6_T1) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n26), .B(
        SubCellInst_SboxInst_6_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_6_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4559), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4561), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4563), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_T1), .B(new_AGEMA_signal_4565), .Z(
        SubCellInst_SboxInst_6_L0) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2206), 
        .B(new_AGEMA_signal_4567), .Z(new_AGEMA_signal_2310) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2207), 
        .B(new_AGEMA_signal_4569), .Z(new_AGEMA_signal_2311) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U37 ( .A(new_AGEMA_signal_2078), .B(
        Fresh[137]), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U36 ( .A(Fresh[136]), .B(
        SubCellInst_SboxInst_6_Q7), .Z(
        SubCellInst_SboxInst_6_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U35 ( .A(new_AGEMA_signal_2079), .B(
        Fresh[137]), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U34 ( .A(Fresh[135]), .B(
        SubCellInst_SboxInst_6_Q7), .Z(
        SubCellInst_SboxInst_6_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U33 ( .A(Fresh[136]), .B(
        new_AGEMA_signal_2079), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U32 ( .A(new_AGEMA_signal_2078), .B(
        Fresh[135]), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U25 ( .A1(new_AGEMA_signal_4575), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U24 ( .A1(new_AGEMA_signal_4575), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U23 ( .A1(new_AGEMA_signal_4573), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND4_U1_U22 ( .A(Fresh[137]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U21 ( .A1(new_AGEMA_signal_4573), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U20 ( .A1(new_AGEMA_signal_4571), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_6_AND4_U1_U19 ( .A(Fresh[136]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U18 ( .A1(new_AGEMA_signal_4571), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND4_U1_U17 ( .A(Fresh[135]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U16 ( .A1(new_AGEMA_signal_2079), 
        .A2(new_AGEMA_signal_4575), .ZN(SubCellInst_SboxInst_6_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U15 ( .A1(new_AGEMA_signal_2078), 
        .A2(new_AGEMA_signal_4573), .ZN(SubCellInst_SboxInst_6_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_6_Q7), 
        .A2(new_AGEMA_signal_4571), .ZN(SubCellInst_SboxInst_6_AND4_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND4_U1_n33), .Z(new_AGEMA_signal_2209) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n32), .B(
        SubCellInst_SboxInst_6_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_6_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_6_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND4_U1_n30), .Z(new_AGEMA_signal_2208) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n29), .B(
        SubCellInst_SboxInst_6_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_6_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND4_U1_n27), .Z(SubCellInst_SboxInst_6_T3) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n26), .B(
        SubCellInst_SboxInst_6_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_6_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4571), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4573), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4575), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L0), .B(new_AGEMA_signal_4579), .Z(
        SubCellInst_SboxInst_6_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2310), 
        .B(new_AGEMA_signal_4583), .Z(new_AGEMA_signal_2396) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2311), 
        .B(new_AGEMA_signal_4587), .Z(new_AGEMA_signal_2397) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L0), .B(SubCellInst_SboxInst_6_T3), .Z(
        ShiftRowsOutput[16]) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2310), 
        .B(new_AGEMA_signal_2208), .Z(new_AGEMA_signal_2398) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2311), 
        .B(new_AGEMA_signal_2209), .Z(new_AGEMA_signal_2399) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_4589), .B(SubCellInst_SboxInst_6_YY_3), .ZN(ShiftRowsOutput[17]) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4591), .B(new_AGEMA_signal_2396), .Z(new_AGEMA_signal_2500) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4593), .B(new_AGEMA_signal_2397), .Z(new_AGEMA_signal_2501) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U37 ( .A(new_AGEMA_signal_2084), .B(
        Fresh[140]), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U36 ( .A(Fresh[139]), .B(
        SubCellInst_SboxInst_7_Q2), .Z(
        SubCellInst_SboxInst_7_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U35 ( .A(new_AGEMA_signal_2085), .B(
        Fresh[140]), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U34 ( .A(Fresh[138]), .B(
        SubCellInst_SboxInst_7_Q2), .Z(
        SubCellInst_SboxInst_7_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U33 ( .A(Fresh[139]), .B(
        new_AGEMA_signal_2085), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U32 ( .A(new_AGEMA_signal_2084), .B(
        Fresh[138]), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U25 ( .A1(new_AGEMA_signal_4599), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U24 ( .A1(new_AGEMA_signal_4599), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U23 ( .A1(new_AGEMA_signal_4597), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND2_U1_U22 ( .A(Fresh[140]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U21 ( .A1(new_AGEMA_signal_4597), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U20 ( .A1(new_AGEMA_signal_4595), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND2_U1_U19 ( .A(Fresh[139]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U18 ( .A1(new_AGEMA_signal_4595), 
        .A2(SubCellInst_SboxInst_7_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND2_U1_U17 ( .A(Fresh[138]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U16 ( .A1(new_AGEMA_signal_2085), 
        .A2(new_AGEMA_signal_4599), .ZN(SubCellInst_SboxInst_7_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U15 ( .A1(new_AGEMA_signal_2084), 
        .A2(new_AGEMA_signal_4597), .ZN(SubCellInst_SboxInst_7_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_7_Q2), 
        .A2(new_AGEMA_signal_4595), .ZN(SubCellInst_SboxInst_7_AND2_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND2_U1_n33), .Z(new_AGEMA_signal_2215) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n32), .B(
        SubCellInst_SboxInst_7_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_7_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND2_U1_n30), .Z(new_AGEMA_signal_2214) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n29), .B(
        SubCellInst_SboxInst_7_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_7_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND2_U1_n27), .Z(SubCellInst_SboxInst_7_T1) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n26), .B(
        SubCellInst_SboxInst_7_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_7_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4595), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4597), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4599), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_T1), .B(new_AGEMA_signal_4601), .Z(
        SubCellInst_SboxInst_7_L0) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2214), 
        .B(new_AGEMA_signal_4603), .Z(new_AGEMA_signal_2314) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2215), 
        .B(new_AGEMA_signal_4605), .Z(new_AGEMA_signal_2315) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U37 ( .A(new_AGEMA_signal_2086), .B(
        Fresh[143]), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U36 ( .A(Fresh[142]), .B(
        SubCellInst_SboxInst_7_Q7), .Z(
        SubCellInst_SboxInst_7_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U35 ( .A(new_AGEMA_signal_2087), .B(
        Fresh[143]), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U34 ( .A(Fresh[141]), .B(
        SubCellInst_SboxInst_7_Q7), .Z(
        SubCellInst_SboxInst_7_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U33 ( .A(Fresh[142]), .B(
        new_AGEMA_signal_2087), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U32 ( .A(new_AGEMA_signal_2086), .B(
        Fresh[141]), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U25 ( .A1(new_AGEMA_signal_4611), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U24 ( .A1(new_AGEMA_signal_4611), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U23 ( .A1(new_AGEMA_signal_4609), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND4_U1_U22 ( .A(Fresh[143]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U21 ( .A1(new_AGEMA_signal_4609), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U20 ( .A1(new_AGEMA_signal_4607), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_7_AND4_U1_U19 ( .A(Fresh[142]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U18 ( .A1(new_AGEMA_signal_4607), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND4_U1_U17 ( .A(Fresh[141]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U16 ( .A1(new_AGEMA_signal_2087), 
        .A2(new_AGEMA_signal_4611), .ZN(SubCellInst_SboxInst_7_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U15 ( .A1(new_AGEMA_signal_2086), 
        .A2(new_AGEMA_signal_4609), .ZN(SubCellInst_SboxInst_7_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_7_Q7), 
        .A2(new_AGEMA_signal_4607), .ZN(SubCellInst_SboxInst_7_AND4_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND4_U1_n33), .Z(new_AGEMA_signal_2217) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n32), .B(
        SubCellInst_SboxInst_7_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_7_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_7_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND4_U1_n30), .Z(new_AGEMA_signal_2216) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n29), .B(
        SubCellInst_SboxInst_7_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_7_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND4_U1_n27), .Z(SubCellInst_SboxInst_7_T3) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n26), .B(
        SubCellInst_SboxInst_7_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_7_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4607), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4609), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4611), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L0), .B(new_AGEMA_signal_4615), .Z(
        SubCellInst_SboxInst_7_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2314), 
        .B(new_AGEMA_signal_4619), .Z(new_AGEMA_signal_2400) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2315), 
        .B(new_AGEMA_signal_4623), .Z(new_AGEMA_signal_2401) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L0), .B(SubCellInst_SboxInst_7_T3), .Z(
        ShiftRowsOutput[20]) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2314), 
        .B(new_AGEMA_signal_2216), .Z(new_AGEMA_signal_2402) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2315), 
        .B(new_AGEMA_signal_2217), .Z(new_AGEMA_signal_2403) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_4625), .B(SubCellInst_SboxInst_7_YY_3), .ZN(SubCellOutput_29) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4627), .B(new_AGEMA_signal_2400), .Z(new_AGEMA_signal_2594) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4629), .B(new_AGEMA_signal_2401), .Z(new_AGEMA_signal_2595) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U37 ( .A(new_AGEMA_signal_2092), .B(
        Fresh[146]), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U36 ( .A(Fresh[145]), .B(
        SubCellInst_SboxInst_8_Q2), .Z(
        SubCellInst_SboxInst_8_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U35 ( .A(new_AGEMA_signal_2093), .B(
        Fresh[146]), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U34 ( .A(Fresh[144]), .B(
        SubCellInst_SboxInst_8_Q2), .Z(
        SubCellInst_SboxInst_8_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U33 ( .A(Fresh[145]), .B(
        new_AGEMA_signal_2093), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U32 ( .A(new_AGEMA_signal_2092), .B(
        Fresh[144]), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U25 ( .A1(new_AGEMA_signal_4635), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U24 ( .A1(new_AGEMA_signal_4635), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U23 ( .A1(new_AGEMA_signal_4633), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND2_U1_U22 ( .A(Fresh[146]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U21 ( .A1(new_AGEMA_signal_4633), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U20 ( .A1(new_AGEMA_signal_4631), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND2_U1_U19 ( .A(Fresh[145]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U18 ( .A1(new_AGEMA_signal_4631), 
        .A2(SubCellInst_SboxInst_8_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND2_U1_U17 ( .A(Fresh[144]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U16 ( .A1(new_AGEMA_signal_2093), 
        .A2(new_AGEMA_signal_4635), .ZN(SubCellInst_SboxInst_8_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U15 ( .A1(new_AGEMA_signal_2092), 
        .A2(new_AGEMA_signal_4633), .ZN(SubCellInst_SboxInst_8_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_8_Q2), 
        .A2(new_AGEMA_signal_4631), .ZN(SubCellInst_SboxInst_8_AND2_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND2_U1_n33), .Z(new_AGEMA_signal_2223) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n32), .B(
        SubCellInst_SboxInst_8_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_8_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND2_U1_n30), .Z(new_AGEMA_signal_2222) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n29), .B(
        SubCellInst_SboxInst_8_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_8_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND2_U1_n27), .Z(SubCellInst_SboxInst_8_T1) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n26), .B(
        SubCellInst_SboxInst_8_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_8_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4631), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4633), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4635), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_T1), .B(new_AGEMA_signal_4637), .Z(
        SubCellInst_SboxInst_8_L0) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2222), 
        .B(new_AGEMA_signal_4639), .Z(new_AGEMA_signal_2318) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2223), 
        .B(new_AGEMA_signal_4641), .Z(new_AGEMA_signal_2319) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U37 ( .A(new_AGEMA_signal_2094), .B(
        Fresh[149]), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U36 ( .A(Fresh[148]), .B(
        SubCellInst_SboxInst_8_Q7), .Z(
        SubCellInst_SboxInst_8_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U35 ( .A(new_AGEMA_signal_2095), .B(
        Fresh[149]), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U34 ( .A(Fresh[147]), .B(
        SubCellInst_SboxInst_8_Q7), .Z(
        SubCellInst_SboxInst_8_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U33 ( .A(Fresh[148]), .B(
        new_AGEMA_signal_2095), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U32 ( .A(new_AGEMA_signal_2094), .B(
        Fresh[147]), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U25 ( .A1(new_AGEMA_signal_4647), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U24 ( .A1(new_AGEMA_signal_4647), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U23 ( .A1(new_AGEMA_signal_4645), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND4_U1_U22 ( .A(Fresh[149]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U21 ( .A1(new_AGEMA_signal_4645), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U20 ( .A1(new_AGEMA_signal_4643), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_8_AND4_U1_U19 ( .A(Fresh[148]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U18 ( .A1(new_AGEMA_signal_4643), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND4_U1_U17 ( .A(Fresh[147]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U16 ( .A1(new_AGEMA_signal_2095), 
        .A2(new_AGEMA_signal_4647), .ZN(SubCellInst_SboxInst_8_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U15 ( .A1(new_AGEMA_signal_2094), 
        .A2(new_AGEMA_signal_4645), .ZN(SubCellInst_SboxInst_8_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_8_Q7), 
        .A2(new_AGEMA_signal_4643), .ZN(SubCellInst_SboxInst_8_AND4_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND4_U1_n33), .Z(new_AGEMA_signal_2225) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n32), .B(
        SubCellInst_SboxInst_8_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_8_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_8_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND4_U1_n30), .Z(new_AGEMA_signal_2224) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n29), .B(
        SubCellInst_SboxInst_8_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_8_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND4_U1_n27), .Z(SubCellInst_SboxInst_8_T3) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n26), .B(
        SubCellInst_SboxInst_8_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_8_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4643), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4645), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4647), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L0), .B(new_AGEMA_signal_4651), .Z(
        SubCellInst_SboxInst_8_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2318), 
        .B(new_AGEMA_signal_4655), .Z(new_AGEMA_signal_2404) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2319), 
        .B(new_AGEMA_signal_4659), .Z(new_AGEMA_signal_2405) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L0), .B(SubCellInst_SboxInst_8_T3), .Z(
        AddRoundConstantOutput[32]) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2318), 
        .B(new_AGEMA_signal_2224), .Z(new_AGEMA_signal_2406) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2319), 
        .B(new_AGEMA_signal_2225), .Z(new_AGEMA_signal_2407) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_4661), .B(SubCellInst_SboxInst_8_YY_3), .ZN(AddRoundConstantOutput[33]) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4663), .B(new_AGEMA_signal_2404), .Z(new_AGEMA_signal_2504) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4665), .B(new_AGEMA_signal_2405), .Z(new_AGEMA_signal_2505) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U37 ( .A(new_AGEMA_signal_2100), .B(
        Fresh[152]), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U36 ( .A(Fresh[151]), .B(
        SubCellInst_SboxInst_9_Q2), .Z(
        SubCellInst_SboxInst_9_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U35 ( .A(new_AGEMA_signal_2101), .B(
        Fresh[152]), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U34 ( .A(Fresh[150]), .B(
        SubCellInst_SboxInst_9_Q2), .Z(
        SubCellInst_SboxInst_9_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U33 ( .A(Fresh[151]), .B(
        new_AGEMA_signal_2101), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U32 ( .A(new_AGEMA_signal_2100), .B(
        Fresh[150]), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U25 ( .A1(new_AGEMA_signal_4671), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U24 ( .A1(new_AGEMA_signal_4671), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U23 ( .A1(new_AGEMA_signal_4669), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND2_U1_U22 ( .A(Fresh[152]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U21 ( .A1(new_AGEMA_signal_4669), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U20 ( .A1(new_AGEMA_signal_4667), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND2_U1_U19 ( .A(Fresh[151]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U18 ( .A1(new_AGEMA_signal_4667), 
        .A2(SubCellInst_SboxInst_9_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND2_U1_U17 ( .A(Fresh[150]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U16 ( .A1(new_AGEMA_signal_2101), 
        .A2(new_AGEMA_signal_4671), .ZN(SubCellInst_SboxInst_9_AND2_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U15 ( .A1(new_AGEMA_signal_2100), 
        .A2(new_AGEMA_signal_4669), .ZN(SubCellInst_SboxInst_9_AND2_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_9_Q2), 
        .A2(new_AGEMA_signal_4667), .ZN(SubCellInst_SboxInst_9_AND2_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND2_U1_n33), .Z(new_AGEMA_signal_2231) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n32), .B(
        SubCellInst_SboxInst_9_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_9_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND2_U1_n30), .Z(new_AGEMA_signal_2230) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n29), .B(
        SubCellInst_SboxInst_9_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_9_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND2_U1_n27), .Z(SubCellInst_SboxInst_9_T1) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n26), .B(
        SubCellInst_SboxInst_9_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_9_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4667), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4669), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4671), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_T1), .B(new_AGEMA_signal_4673), .Z(
        SubCellInst_SboxInst_9_L0) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2230), 
        .B(new_AGEMA_signal_4675), .Z(new_AGEMA_signal_2322) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2231), 
        .B(new_AGEMA_signal_4677), .Z(new_AGEMA_signal_2323) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U37 ( .A(new_AGEMA_signal_2102), .B(
        Fresh[155]), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U36 ( .A(Fresh[154]), .B(
        SubCellInst_SboxInst_9_Q7), .Z(
        SubCellInst_SboxInst_9_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U35 ( .A(new_AGEMA_signal_2103), .B(
        Fresh[155]), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U34 ( .A(Fresh[153]), .B(
        SubCellInst_SboxInst_9_Q7), .Z(
        SubCellInst_SboxInst_9_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U33 ( .A(Fresh[154]), .B(
        new_AGEMA_signal_2103), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U32 ( .A(new_AGEMA_signal_2102), .B(
        Fresh[153]), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U25 ( .A1(new_AGEMA_signal_4683), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U24 ( .A1(new_AGEMA_signal_4683), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U23 ( .A1(new_AGEMA_signal_4681), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND4_U1_U22 ( .A(Fresh[155]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U21 ( .A1(new_AGEMA_signal_4681), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U20 ( .A1(new_AGEMA_signal_4679), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_9_AND4_U1_U19 ( .A(Fresh[154]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U18 ( .A1(new_AGEMA_signal_4679), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND4_U1_U17 ( .A(Fresh[153]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U16 ( .A1(new_AGEMA_signal_2103), 
        .A2(new_AGEMA_signal_4683), .ZN(SubCellInst_SboxInst_9_AND4_U1_mul[2])
         );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U15 ( .A1(new_AGEMA_signal_2102), 
        .A2(new_AGEMA_signal_4681), .ZN(SubCellInst_SboxInst_9_AND4_U1_mul[1])
         );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_9_Q7), 
        .A2(new_AGEMA_signal_4679), .ZN(SubCellInst_SboxInst_9_AND4_U1_mul[0])
         );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND4_U1_n33), .Z(new_AGEMA_signal_2233) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n32), .B(
        SubCellInst_SboxInst_9_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_9_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_9_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND4_U1_n30), .Z(new_AGEMA_signal_2232) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n29), .B(
        SubCellInst_SboxInst_9_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_9_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND4_U1_n27), .Z(SubCellInst_SboxInst_9_T3) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n26), .B(
        SubCellInst_SboxInst_9_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_9_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4679), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4681), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4683), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L0), .B(new_AGEMA_signal_4687), .Z(
        SubCellInst_SboxInst_9_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2322), 
        .B(new_AGEMA_signal_4691), .Z(new_AGEMA_signal_2408) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2323), 
        .B(new_AGEMA_signal_4695), .Z(new_AGEMA_signal_2409) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L0), .B(SubCellInst_SboxInst_9_T3), .Z(
        AddRoundConstantOutput[36]) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2322), 
        .B(new_AGEMA_signal_2232), .Z(new_AGEMA_signal_2410) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2323), 
        .B(new_AGEMA_signal_2233), .Z(new_AGEMA_signal_2411) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR_o1_U1_Ins0_U1 ( .A(new_AGEMA_signal_4697), .B(SubCellInst_SboxInst_9_YY_3), .ZN(AddRoundConstantOutput[37]) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_4699), .B(new_AGEMA_signal_2408), .Z(new_AGEMA_signal_2506) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_o1_U1_Ins_2_U1 ( .A(new_AGEMA_signal_4701), .B(new_AGEMA_signal_2409), .Z(new_AGEMA_signal_2507) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U37 ( .A(new_AGEMA_signal_2108), .B(
        Fresh[158]), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U36 ( .A(Fresh[157]), .B(
        SubCellInst_SboxInst_10_Q2), .Z(
        SubCellInst_SboxInst_10_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U35 ( .A(new_AGEMA_signal_2109), .B(
        Fresh[158]), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U34 ( .A(Fresh[156]), .B(
        SubCellInst_SboxInst_10_Q2), .Z(
        SubCellInst_SboxInst_10_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U33 ( .A(Fresh[157]), .B(
        new_AGEMA_signal_2109), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U32 ( .A(new_AGEMA_signal_2108), .B(
        Fresh[156]), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U25 ( .A1(new_AGEMA_signal_4707), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U24 ( .A1(new_AGEMA_signal_4707), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U23 ( .A1(new_AGEMA_signal_4705), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND2_U1_U22 ( .A(Fresh[158]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U21 ( .A1(new_AGEMA_signal_4705), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U20 ( .A1(new_AGEMA_signal_4703), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND2_U1_U19 ( .A(Fresh[157]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U18 ( .A1(new_AGEMA_signal_4703), 
        .A2(SubCellInst_SboxInst_10_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND2_U1_U17 ( .A(Fresh[156]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U16 ( .A1(new_AGEMA_signal_2109), 
        .A2(new_AGEMA_signal_4707), .ZN(SubCellInst_SboxInst_10_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U15 ( .A1(new_AGEMA_signal_2108), 
        .A2(new_AGEMA_signal_4705), .ZN(SubCellInst_SboxInst_10_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_10_Q2), .A2(new_AGEMA_signal_4703), .ZN(SubCellInst_SboxInst_10_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND2_U1_n33), .Z(new_AGEMA_signal_2239) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n32), .B(
        SubCellInst_SboxInst_10_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_10_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND2_U1_n30), .Z(new_AGEMA_signal_2238) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n29), .B(
        SubCellInst_SboxInst_10_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_10_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND2_U1_n27), .Z(SubCellInst_SboxInst_10_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n26), .B(
        SubCellInst_SboxInst_10_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_10_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4703), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4705), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4707), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_T1), .B(new_AGEMA_signal_4709), .Z(
        SubCellInst_SboxInst_10_L0) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2238), 
        .B(new_AGEMA_signal_4711), .Z(new_AGEMA_signal_2326) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2239), 
        .B(new_AGEMA_signal_4713), .Z(new_AGEMA_signal_2327) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U37 ( .A(new_AGEMA_signal_2110), .B(
        Fresh[161]), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U36 ( .A(Fresh[160]), .B(
        SubCellInst_SboxInst_10_Q7), .Z(
        SubCellInst_SboxInst_10_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U35 ( .A(new_AGEMA_signal_2111), .B(
        Fresh[161]), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U34 ( .A(Fresh[159]), .B(
        SubCellInst_SboxInst_10_Q7), .Z(
        SubCellInst_SboxInst_10_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U33 ( .A(Fresh[160]), .B(
        new_AGEMA_signal_2111), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U32 ( .A(new_AGEMA_signal_2110), .B(
        Fresh[159]), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U25 ( .A1(new_AGEMA_signal_4719), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U24 ( .A1(new_AGEMA_signal_4719), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U23 ( .A1(new_AGEMA_signal_4717), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND4_U1_U22 ( .A(Fresh[161]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U21 ( .A1(new_AGEMA_signal_4717), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U20 ( .A1(new_AGEMA_signal_4715), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_10_AND4_U1_U19 ( .A(Fresh[160]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U18 ( .A1(new_AGEMA_signal_4715), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND4_U1_U17 ( .A(Fresh[159]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U16 ( .A1(new_AGEMA_signal_2111), 
        .A2(new_AGEMA_signal_4719), .ZN(SubCellInst_SboxInst_10_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U15 ( .A1(new_AGEMA_signal_2110), 
        .A2(new_AGEMA_signal_4717), .ZN(SubCellInst_SboxInst_10_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_10_Q7), .A2(new_AGEMA_signal_4715), .ZN(SubCellInst_SboxInst_10_AND4_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND4_U1_n33), .Z(new_AGEMA_signal_2241) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n32), .B(
        SubCellInst_SboxInst_10_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_10_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_10_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND4_U1_n30), .Z(new_AGEMA_signal_2240) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n29), .B(
        SubCellInst_SboxInst_10_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_10_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND4_U1_n27), .Z(SubCellInst_SboxInst_10_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n26), .B(
        SubCellInst_SboxInst_10_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_10_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4715), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4717), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4719), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L0), .B(new_AGEMA_signal_4723), .Z(
        SubCellInst_SboxInst_10_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2326), 
        .B(new_AGEMA_signal_4727), .Z(new_AGEMA_signal_2412) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2327), 
        .B(new_AGEMA_signal_4731), .Z(new_AGEMA_signal_2413) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L0), .B(SubCellInst_SboxInst_10_T3), .Z(
        AddRoundConstantOutput[40]) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2326), .B(new_AGEMA_signal_2240), .Z(new_AGEMA_signal_2414) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2327), .B(new_AGEMA_signal_2241), .Z(new_AGEMA_signal_2415) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_4733), .B(SubCellInst_SboxInst_10_YY_3), .ZN(
        AddRoundConstantOutput[41]) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_4735), .B(new_AGEMA_signal_2412), .Z(
        new_AGEMA_signal_2508) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_4737), .B(new_AGEMA_signal_2413), .Z(
        new_AGEMA_signal_2509) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U37 ( .A(new_AGEMA_signal_2116), .B(
        Fresh[164]), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U36 ( .A(Fresh[163]), .B(
        SubCellInst_SboxInst_11_Q2), .Z(
        SubCellInst_SboxInst_11_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U35 ( .A(new_AGEMA_signal_2117), .B(
        Fresh[164]), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U34 ( .A(Fresh[162]), .B(
        SubCellInst_SboxInst_11_Q2), .Z(
        SubCellInst_SboxInst_11_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U33 ( .A(Fresh[163]), .B(
        new_AGEMA_signal_2117), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U32 ( .A(new_AGEMA_signal_2116), .B(
        Fresh[162]), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U25 ( .A1(new_AGEMA_signal_4743), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U24 ( .A1(new_AGEMA_signal_4743), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U23 ( .A1(new_AGEMA_signal_4741), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND2_U1_U22 ( .A(Fresh[164]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U21 ( .A1(new_AGEMA_signal_4741), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U20 ( .A1(new_AGEMA_signal_4739), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND2_U1_U19 ( .A(Fresh[163]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U18 ( .A1(new_AGEMA_signal_4739), 
        .A2(SubCellInst_SboxInst_11_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND2_U1_U17 ( .A(Fresh[162]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U16 ( .A1(new_AGEMA_signal_2117), 
        .A2(new_AGEMA_signal_4743), .ZN(SubCellInst_SboxInst_11_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U15 ( .A1(new_AGEMA_signal_2116), 
        .A2(new_AGEMA_signal_4741), .ZN(SubCellInst_SboxInst_11_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_11_Q2), .A2(new_AGEMA_signal_4739), .ZN(SubCellInst_SboxInst_11_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND2_U1_n33), .Z(new_AGEMA_signal_2247) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n32), .B(
        SubCellInst_SboxInst_11_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_11_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND2_U1_n30), .Z(new_AGEMA_signal_2246) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n29), .B(
        SubCellInst_SboxInst_11_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_11_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND2_U1_n27), .Z(SubCellInst_SboxInst_11_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n26), .B(
        SubCellInst_SboxInst_11_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_11_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4739), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4741), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4743), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_T1), .B(new_AGEMA_signal_4745), .Z(
        SubCellInst_SboxInst_11_L0) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2246), 
        .B(new_AGEMA_signal_4747), .Z(new_AGEMA_signal_2330) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2247), 
        .B(new_AGEMA_signal_4749), .Z(new_AGEMA_signal_2331) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U37 ( .A(new_AGEMA_signal_2118), .B(
        Fresh[167]), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U36 ( .A(Fresh[166]), .B(
        SubCellInst_SboxInst_11_Q7), .Z(
        SubCellInst_SboxInst_11_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U35 ( .A(new_AGEMA_signal_2119), .B(
        Fresh[167]), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U34 ( .A(Fresh[165]), .B(
        SubCellInst_SboxInst_11_Q7), .Z(
        SubCellInst_SboxInst_11_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U33 ( .A(Fresh[166]), .B(
        new_AGEMA_signal_2119), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U32 ( .A(new_AGEMA_signal_2118), .B(
        Fresh[165]), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U25 ( .A1(new_AGEMA_signal_4755), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U24 ( .A1(new_AGEMA_signal_4755), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U23 ( .A1(new_AGEMA_signal_4753), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND4_U1_U22 ( .A(Fresh[167]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U21 ( .A1(new_AGEMA_signal_4753), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U20 ( .A1(new_AGEMA_signal_4751), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_11_AND4_U1_U19 ( .A(Fresh[166]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U18 ( .A1(new_AGEMA_signal_4751), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND4_U1_U17 ( .A(Fresh[165]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U16 ( .A1(new_AGEMA_signal_2119), 
        .A2(new_AGEMA_signal_4755), .ZN(SubCellInst_SboxInst_11_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U15 ( .A1(new_AGEMA_signal_2118), 
        .A2(new_AGEMA_signal_4753), .ZN(SubCellInst_SboxInst_11_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_11_Q7), .A2(new_AGEMA_signal_4751), .ZN(SubCellInst_SboxInst_11_AND4_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND4_U1_n33), .Z(new_AGEMA_signal_2249) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n32), .B(
        SubCellInst_SboxInst_11_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_11_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_11_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND4_U1_n30), .Z(new_AGEMA_signal_2248) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n29), .B(
        SubCellInst_SboxInst_11_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_11_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND4_U1_n27), .Z(SubCellInst_SboxInst_11_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n26), .B(
        SubCellInst_SboxInst_11_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_11_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4751), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4753), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4755), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L0), .B(new_AGEMA_signal_4759), .Z(
        SubCellInst_SboxInst_11_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2330), 
        .B(new_AGEMA_signal_4763), .Z(new_AGEMA_signal_2416) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2331), 
        .B(new_AGEMA_signal_4767), .Z(new_AGEMA_signal_2417) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L0), .B(SubCellInst_SboxInst_11_T3), .Z(
        SubCellOutput_44) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2330), .B(new_AGEMA_signal_2248), .Z(new_AGEMA_signal_2418) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2331), .B(new_AGEMA_signal_2249), .Z(new_AGEMA_signal_2419) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_4769), .B(SubCellInst_SboxInst_11_YY_3), .ZN(
        SubCellOutput_45) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_4771), .B(new_AGEMA_signal_2416), .Z(
        new_AGEMA_signal_2510) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_4773), .B(new_AGEMA_signal_2417), .Z(
        new_AGEMA_signal_2511) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U37 ( .A(new_AGEMA_signal_2124), .B(
        Fresh[170]), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U36 ( .A(Fresh[169]), .B(
        SubCellInst_SboxInst_12_Q2), .Z(
        SubCellInst_SboxInst_12_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U35 ( .A(new_AGEMA_signal_2125), .B(
        Fresh[170]), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U34 ( .A(Fresh[168]), .B(
        SubCellInst_SboxInst_12_Q2), .Z(
        SubCellInst_SboxInst_12_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U33 ( .A(Fresh[169]), .B(
        new_AGEMA_signal_2125), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U32 ( .A(new_AGEMA_signal_2124), .B(
        Fresh[168]), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U25 ( .A1(new_AGEMA_signal_4779), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U24 ( .A1(new_AGEMA_signal_4779), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U23 ( .A1(new_AGEMA_signal_4777), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND2_U1_U22 ( .A(Fresh[170]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U21 ( .A1(new_AGEMA_signal_4777), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U20 ( .A1(new_AGEMA_signal_4775), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND2_U1_U19 ( .A(Fresh[169]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U18 ( .A1(new_AGEMA_signal_4775), 
        .A2(SubCellInst_SboxInst_12_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND2_U1_U17 ( .A(Fresh[168]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U16 ( .A1(new_AGEMA_signal_2125), 
        .A2(new_AGEMA_signal_4779), .ZN(SubCellInst_SboxInst_12_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U15 ( .A1(new_AGEMA_signal_2124), 
        .A2(new_AGEMA_signal_4777), .ZN(SubCellInst_SboxInst_12_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_12_Q2), .A2(new_AGEMA_signal_4775), .ZN(SubCellInst_SboxInst_12_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND2_U1_n33), .Z(new_AGEMA_signal_2255) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n32), .B(
        SubCellInst_SboxInst_12_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_12_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND2_U1_n30), .Z(new_AGEMA_signal_2254) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n29), .B(
        SubCellInst_SboxInst_12_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_12_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND2_U1_n27), .Z(SubCellInst_SboxInst_12_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n26), .B(
        SubCellInst_SboxInst_12_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_12_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4775), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4777), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4779), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_T1), .B(new_AGEMA_signal_4781), .Z(
        SubCellInst_SboxInst_12_L0) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2254), 
        .B(new_AGEMA_signal_4783), .Z(new_AGEMA_signal_2334) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2255), 
        .B(new_AGEMA_signal_4785), .Z(new_AGEMA_signal_2335) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U37 ( .A(new_AGEMA_signal_2126), .B(
        Fresh[173]), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U36 ( .A(Fresh[172]), .B(
        SubCellInst_SboxInst_12_Q7), .Z(
        SubCellInst_SboxInst_12_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U35 ( .A(new_AGEMA_signal_2127), .B(
        Fresh[173]), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U34 ( .A(Fresh[171]), .B(
        SubCellInst_SboxInst_12_Q7), .Z(
        SubCellInst_SboxInst_12_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U33 ( .A(Fresh[172]), .B(
        new_AGEMA_signal_2127), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U32 ( .A(new_AGEMA_signal_2126), .B(
        Fresh[171]), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U25 ( .A1(new_AGEMA_signal_4791), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U24 ( .A1(new_AGEMA_signal_4791), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U23 ( .A1(new_AGEMA_signal_4789), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND4_U1_U22 ( .A(Fresh[173]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U21 ( .A1(new_AGEMA_signal_4789), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U20 ( .A1(new_AGEMA_signal_4787), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_12_AND4_U1_U19 ( .A(Fresh[172]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U18 ( .A1(new_AGEMA_signal_4787), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND4_U1_U17 ( .A(Fresh[171]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U16 ( .A1(new_AGEMA_signal_2127), 
        .A2(new_AGEMA_signal_4791), .ZN(SubCellInst_SboxInst_12_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U15 ( .A1(new_AGEMA_signal_2126), 
        .A2(new_AGEMA_signal_4789), .ZN(SubCellInst_SboxInst_12_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_12_Q7), .A2(new_AGEMA_signal_4787), .ZN(SubCellInst_SboxInst_12_AND4_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND4_U1_n33), .Z(new_AGEMA_signal_2257) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n32), .B(
        SubCellInst_SboxInst_12_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_12_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_12_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND4_U1_n30), .Z(new_AGEMA_signal_2256) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n29), .B(
        SubCellInst_SboxInst_12_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_12_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND4_U1_n27), .Z(SubCellInst_SboxInst_12_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n26), .B(
        SubCellInst_SboxInst_12_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_12_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4787), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4789), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4791), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L0), .B(new_AGEMA_signal_4795), .Z(
        SubCellInst_SboxInst_12_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2334), 
        .B(new_AGEMA_signal_4799), .Z(new_AGEMA_signal_2420) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2335), 
        .B(new_AGEMA_signal_4803), .Z(new_AGEMA_signal_2421) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L0), .B(SubCellInst_SboxInst_12_T3), .Z(
        AddRoundConstantOutput[48]) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2334), .B(new_AGEMA_signal_2256), .Z(new_AGEMA_signal_2422) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2335), .B(new_AGEMA_signal_2257), .Z(new_AGEMA_signal_2423) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_4805), .B(SubCellInst_SboxInst_12_YY_3), .ZN(
        AddRoundConstantOutput[49]) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_4807), .B(new_AGEMA_signal_2420), .Z(
        new_AGEMA_signal_2512) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_4809), .B(new_AGEMA_signal_2421), .Z(
        new_AGEMA_signal_2513) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U37 ( .A(new_AGEMA_signal_2132), .B(
        Fresh[176]), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U36 ( .A(Fresh[175]), .B(
        SubCellInst_SboxInst_13_Q2), .Z(
        SubCellInst_SboxInst_13_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U35 ( .A(new_AGEMA_signal_2133), .B(
        Fresh[176]), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U34 ( .A(Fresh[174]), .B(
        SubCellInst_SboxInst_13_Q2), .Z(
        SubCellInst_SboxInst_13_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U33 ( .A(Fresh[175]), .B(
        new_AGEMA_signal_2133), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U32 ( .A(new_AGEMA_signal_2132), .B(
        Fresh[174]), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U25 ( .A1(new_AGEMA_signal_4815), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U24 ( .A1(new_AGEMA_signal_4815), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U23 ( .A1(new_AGEMA_signal_4813), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND2_U1_U22 ( .A(Fresh[176]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U21 ( .A1(new_AGEMA_signal_4813), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U20 ( .A1(new_AGEMA_signal_4811), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND2_U1_U19 ( .A(Fresh[175]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U18 ( .A1(new_AGEMA_signal_4811), 
        .A2(SubCellInst_SboxInst_13_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND2_U1_U17 ( .A(Fresh[174]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U16 ( .A1(new_AGEMA_signal_2133), 
        .A2(new_AGEMA_signal_4815), .ZN(SubCellInst_SboxInst_13_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U15 ( .A1(new_AGEMA_signal_2132), 
        .A2(new_AGEMA_signal_4813), .ZN(SubCellInst_SboxInst_13_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_13_Q2), .A2(new_AGEMA_signal_4811), .ZN(SubCellInst_SboxInst_13_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND2_U1_n33), .Z(new_AGEMA_signal_2263) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n32), .B(
        SubCellInst_SboxInst_13_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_13_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND2_U1_n30), .Z(new_AGEMA_signal_2262) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n29), .B(
        SubCellInst_SboxInst_13_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_13_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND2_U1_n27), .Z(SubCellInst_SboxInst_13_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n26), .B(
        SubCellInst_SboxInst_13_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_13_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4811), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4813), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4815), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_T1), .B(new_AGEMA_signal_4817), .Z(
        SubCellInst_SboxInst_13_L0) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2262), 
        .B(new_AGEMA_signal_4819), .Z(new_AGEMA_signal_2338) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2263), 
        .B(new_AGEMA_signal_4821), .Z(new_AGEMA_signal_2339) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U37 ( .A(new_AGEMA_signal_2134), .B(
        Fresh[179]), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U36 ( .A(Fresh[178]), .B(
        SubCellInst_SboxInst_13_Q7), .Z(
        SubCellInst_SboxInst_13_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U35 ( .A(new_AGEMA_signal_2135), .B(
        Fresh[179]), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U34 ( .A(Fresh[177]), .B(
        SubCellInst_SboxInst_13_Q7), .Z(
        SubCellInst_SboxInst_13_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U33 ( .A(Fresh[178]), .B(
        new_AGEMA_signal_2135), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U32 ( .A(new_AGEMA_signal_2134), .B(
        Fresh[177]), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U25 ( .A1(new_AGEMA_signal_4827), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U24 ( .A1(new_AGEMA_signal_4827), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U23 ( .A1(new_AGEMA_signal_4825), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND4_U1_U22 ( .A(Fresh[179]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U21 ( .A1(new_AGEMA_signal_4825), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U20 ( .A1(new_AGEMA_signal_4823), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_13_AND4_U1_U19 ( .A(Fresh[178]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U18 ( .A1(new_AGEMA_signal_4823), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND4_U1_U17 ( .A(Fresh[177]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U16 ( .A1(new_AGEMA_signal_2135), 
        .A2(new_AGEMA_signal_4827), .ZN(SubCellInst_SboxInst_13_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U15 ( .A1(new_AGEMA_signal_2134), 
        .A2(new_AGEMA_signal_4825), .ZN(SubCellInst_SboxInst_13_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_13_Q7), .A2(new_AGEMA_signal_4823), .ZN(SubCellInst_SboxInst_13_AND4_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND4_U1_n33), .Z(new_AGEMA_signal_2265) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n32), .B(
        SubCellInst_SboxInst_13_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_13_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_13_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND4_U1_n30), .Z(new_AGEMA_signal_2264) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n29), .B(
        SubCellInst_SboxInst_13_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_13_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND4_U1_n27), .Z(SubCellInst_SboxInst_13_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n26), .B(
        SubCellInst_SboxInst_13_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_13_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4823), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4825), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4827), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L0), .B(new_AGEMA_signal_4831), .Z(
        SubCellInst_SboxInst_13_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2338), 
        .B(new_AGEMA_signal_4835), .Z(new_AGEMA_signal_2424) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2339), 
        .B(new_AGEMA_signal_4839), .Z(new_AGEMA_signal_2425) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L0), .B(SubCellInst_SboxInst_13_T3), .Z(
        AddRoundConstantOutput[52]) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2338), .B(new_AGEMA_signal_2264), .Z(new_AGEMA_signal_2426) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2339), .B(new_AGEMA_signal_2265), .Z(new_AGEMA_signal_2427) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_4841), .B(SubCellInst_SboxInst_13_YY_3), .ZN(
        AddRoundConstantOutput[53]) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_4843), .B(new_AGEMA_signal_2424), .Z(
        new_AGEMA_signal_2514) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_4845), .B(new_AGEMA_signal_2425), .Z(
        new_AGEMA_signal_2515) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U37 ( .A(new_AGEMA_signal_2140), .B(
        Fresh[182]), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U36 ( .A(Fresh[181]), .B(
        SubCellInst_SboxInst_14_Q2), .Z(
        SubCellInst_SboxInst_14_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U35 ( .A(new_AGEMA_signal_2141), .B(
        Fresh[182]), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U34 ( .A(Fresh[180]), .B(
        SubCellInst_SboxInst_14_Q2), .Z(
        SubCellInst_SboxInst_14_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U33 ( .A(Fresh[181]), .B(
        new_AGEMA_signal_2141), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U32 ( .A(new_AGEMA_signal_2140), .B(
        Fresh[180]), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U25 ( .A1(new_AGEMA_signal_4851), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U24 ( .A1(new_AGEMA_signal_4851), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U23 ( .A1(new_AGEMA_signal_4849), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND2_U1_U22 ( .A(Fresh[182]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U21 ( .A1(new_AGEMA_signal_4849), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U20 ( .A1(new_AGEMA_signal_4847), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND2_U1_U19 ( .A(Fresh[181]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U18 ( .A1(new_AGEMA_signal_4847), 
        .A2(SubCellInst_SboxInst_14_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND2_U1_U17 ( .A(Fresh[180]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U16 ( .A1(new_AGEMA_signal_2141), 
        .A2(new_AGEMA_signal_4851), .ZN(SubCellInst_SboxInst_14_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U15 ( .A1(new_AGEMA_signal_2140), 
        .A2(new_AGEMA_signal_4849), .ZN(SubCellInst_SboxInst_14_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_14_Q2), .A2(new_AGEMA_signal_4847), .ZN(SubCellInst_SboxInst_14_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND2_U1_n33), .Z(new_AGEMA_signal_2271) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n32), .B(
        SubCellInst_SboxInst_14_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_14_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND2_U1_n30), .Z(new_AGEMA_signal_2270) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n29), .B(
        SubCellInst_SboxInst_14_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_14_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND2_U1_n27), .Z(SubCellInst_SboxInst_14_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n26), .B(
        SubCellInst_SboxInst_14_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_14_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4847), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4849), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4851), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_T1), .B(new_AGEMA_signal_4853), .Z(
        SubCellInst_SboxInst_14_L0) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2270), 
        .B(new_AGEMA_signal_4855), .Z(new_AGEMA_signal_2342) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2271), 
        .B(new_AGEMA_signal_4857), .Z(new_AGEMA_signal_2343) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U37 ( .A(new_AGEMA_signal_2142), .B(
        Fresh[185]), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U36 ( .A(Fresh[184]), .B(
        SubCellInst_SboxInst_14_Q7), .Z(
        SubCellInst_SboxInst_14_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U35 ( .A(new_AGEMA_signal_2143), .B(
        Fresh[185]), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U34 ( .A(Fresh[183]), .B(
        SubCellInst_SboxInst_14_Q7), .Z(
        SubCellInst_SboxInst_14_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U33 ( .A(Fresh[184]), .B(
        new_AGEMA_signal_2143), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U32 ( .A(new_AGEMA_signal_2142), .B(
        Fresh[183]), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U25 ( .A1(new_AGEMA_signal_4863), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U24 ( .A1(new_AGEMA_signal_4863), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U23 ( .A1(new_AGEMA_signal_4861), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND4_U1_U22 ( .A(Fresh[185]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U21 ( .A1(new_AGEMA_signal_4861), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U20 ( .A1(new_AGEMA_signal_4859), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_14_AND4_U1_U19 ( .A(Fresh[184]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U18 ( .A1(new_AGEMA_signal_4859), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND4_U1_U17 ( .A(Fresh[183]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U16 ( .A1(new_AGEMA_signal_2143), 
        .A2(new_AGEMA_signal_4863), .ZN(SubCellInst_SboxInst_14_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U15 ( .A1(new_AGEMA_signal_2142), 
        .A2(new_AGEMA_signal_4861), .ZN(SubCellInst_SboxInst_14_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_14_Q7), .A2(new_AGEMA_signal_4859), .ZN(SubCellInst_SboxInst_14_AND4_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND4_U1_n33), .Z(new_AGEMA_signal_2273) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n32), .B(
        SubCellInst_SboxInst_14_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_14_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_14_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND4_U1_n30), .Z(new_AGEMA_signal_2272) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n29), .B(
        SubCellInst_SboxInst_14_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_14_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND4_U1_n27), .Z(SubCellInst_SboxInst_14_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n26), .B(
        SubCellInst_SboxInst_14_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_14_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4859), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4861), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4863), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L0), .B(new_AGEMA_signal_4867), .Z(
        SubCellInst_SboxInst_14_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2342), 
        .B(new_AGEMA_signal_4871), .Z(new_AGEMA_signal_2428) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2343), 
        .B(new_AGEMA_signal_4875), .Z(new_AGEMA_signal_2429) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L0), .B(SubCellInst_SboxInst_14_T3), .Z(
        AddRoundConstantOutput[56]) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2342), .B(new_AGEMA_signal_2272), .Z(new_AGEMA_signal_2430) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2343), .B(new_AGEMA_signal_2273), .Z(new_AGEMA_signal_2431) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_4877), .B(SubCellInst_SboxInst_14_YY_3), .ZN(
        AddRoundConstantOutput[57]) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_4879), .B(new_AGEMA_signal_2428), .Z(
        new_AGEMA_signal_2516) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_4881), .B(new_AGEMA_signal_2429), .Z(
        new_AGEMA_signal_2517) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U37 ( .A(new_AGEMA_signal_2148), .B(
        Fresh[188]), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U36 ( .A(Fresh[187]), .B(
        SubCellInst_SboxInst_15_Q2), .Z(
        SubCellInst_SboxInst_15_AND2_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U35 ( .A(new_AGEMA_signal_2149), .B(
        Fresh[188]), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U34 ( .A(Fresh[186]), .B(
        SubCellInst_SboxInst_15_Q2), .Z(
        SubCellInst_SboxInst_15_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U33 ( .A(Fresh[187]), .B(
        new_AGEMA_signal_2149), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U32 ( .A(new_AGEMA_signal_2148), .B(
        Fresh[186]), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U31 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U30 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U29 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U28 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U27 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U26 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U25 ( .A1(new_AGEMA_signal_4887), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U24 ( .A1(new_AGEMA_signal_4887), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U23 ( .A1(new_AGEMA_signal_4885), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n36), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND2_U1_U22 ( .A(Fresh[188]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U21 ( .A1(new_AGEMA_signal_4885), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U20 ( .A1(new_AGEMA_signal_4883), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n35), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND2_U1_U19 ( .A(Fresh[187]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U18 ( .A1(new_AGEMA_signal_4883), 
        .A2(SubCellInst_SboxInst_15_AND2_U1_n34), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND2_U1_U17 ( .A(Fresh[186]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U16 ( .A1(new_AGEMA_signal_2149), 
        .A2(new_AGEMA_signal_4887), .ZN(SubCellInst_SboxInst_15_AND2_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U15 ( .A1(new_AGEMA_signal_2148), 
        .A2(new_AGEMA_signal_4885), .ZN(SubCellInst_SboxInst_15_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U14 ( .A1(SubCellInst_SboxInst_15_Q2), .A2(new_AGEMA_signal_4883), .ZN(SubCellInst_SboxInst_15_AND2_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U13 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND2_U1_n33), .Z(new_AGEMA_signal_2279) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U12 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n32), .B(
        SubCellInst_SboxInst_15_AND2_U1_n31), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U11 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND2_U1_z[2]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U10 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_15_AND2_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U9 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND2_U1_n30), .Z(new_AGEMA_signal_2278) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U8 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n29), .B(
        SubCellInst_SboxInst_15_AND2_U1_n28), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U7 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND2_U1_z[1]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U6 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_15_AND2_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND2_U1_n27), .Z(SubCellInst_SboxInst_15_T1)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n26), .B(
        SubCellInst_SboxInst_15_AND2_U1_n25), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND2_U1_z[0]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_15_AND2_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4883), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4885), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4887), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_T1), .B(new_AGEMA_signal_4889), .Z(
        SubCellInst_SboxInst_15_L0) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2278), 
        .B(new_AGEMA_signal_4891), .Z(new_AGEMA_signal_2346) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR4_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2279), 
        .B(new_AGEMA_signal_4893), .Z(new_AGEMA_signal_2347) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U37 ( .A(new_AGEMA_signal_2150), .B(
        Fresh[191]), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_2__1_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U36 ( .A(Fresh[190]), .B(
        SubCellInst_SboxInst_15_Q7), .Z(
        SubCellInst_SboxInst_15_AND4_U1_s_in_2__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U35 ( .A(new_AGEMA_signal_2151), .B(
        Fresh[191]), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_1__2_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U34 ( .A(Fresh[189]), .B(
        SubCellInst_SboxInst_15_Q7), .Z(
        SubCellInst_SboxInst_15_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U33 ( .A(Fresh[190]), .B(
        new_AGEMA_signal_2151), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_0__2_)
         );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U32 ( .A(new_AGEMA_signal_2150), .B(
        Fresh[189]), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_0__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U31 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_2__1_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__1_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U30 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_2_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_2__0_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U29 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__2_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U28 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_1_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U27 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__2_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__2_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U26 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_0_), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U25 ( .A1(new_AGEMA_signal_4899), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U24 ( .A1(new_AGEMA_signal_4899), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U23 ( .A1(new_AGEMA_signal_4897), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n36), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND4_U1_U22 ( .A(Fresh[191]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n36) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U21 ( .A1(new_AGEMA_signal_4897), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U20 ( .A1(new_AGEMA_signal_4895), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n35), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__2_) );
  INV_X1 SubCellInst_SboxInst_15_AND4_U1_U19 ( .A(Fresh[190]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n35) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U18 ( .A1(new_AGEMA_signal_4895), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n34), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND4_U1_U17 ( .A(Fresh[189]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n34) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U16 ( .A1(new_AGEMA_signal_2151), 
        .A2(new_AGEMA_signal_4899), .ZN(SubCellInst_SboxInst_15_AND4_U1_mul[2]) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U15 ( .A1(new_AGEMA_signal_2150), 
        .A2(new_AGEMA_signal_4897), .ZN(SubCellInst_SboxInst_15_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U14 ( .A1(SubCellInst_SboxInst_15_Q7), .A2(new_AGEMA_signal_4895), .ZN(SubCellInst_SboxInst_15_AND4_U1_mul[0]) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U13 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND4_U1_n33), .Z(new_AGEMA_signal_2281) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U12 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n32), .B(
        SubCellInst_SboxInst_15_AND4_U1_n31), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n33) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U11 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__0_), .B(
        SubCellInst_SboxInst_15_AND4_U1_z[2]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n31) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U10 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__1_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__1_), .Z(
        SubCellInst_SboxInst_15_AND4_U1_n32) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U9 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND4_U1_n30), .Z(new_AGEMA_signal_2280) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U8 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n29), .B(
        SubCellInst_SboxInst_15_AND4_U1_n28), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n30) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U7 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND4_U1_z[1]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n28) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U6 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__2_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__2_), .Z(
        SubCellInst_SboxInst_15_AND4_U1_n29) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND4_U1_n27), .Z(SubCellInst_SboxInst_15_T3)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n26), .B(
        SubCellInst_SboxInst_15_AND4_U1_n25), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n27) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND4_U1_z[0]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n25) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__2_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__2_), .Z(
        SubCellInst_SboxInst_15_AND4_U1_n26) );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_z[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_a_i_0_s_current_state_reg ( .D(
        new_AGEMA_signal_4895), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_0_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_0_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_z[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_4897), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_1_2_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__2_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s1_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s2_2_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_z[2]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_a_i_2_s_current_state_reg ( .D(
        new_AGEMA_signal_4899), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_a_reg_2_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_2_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_2_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_2__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_2__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_2__1_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L0), .B(new_AGEMA_signal_4903), .Z(
        SubCellInst_SboxInst_15_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2346), 
        .B(new_AGEMA_signal_4907), .Z(new_AGEMA_signal_2432) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR9_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2347), 
        .B(new_AGEMA_signal_4911), .Z(new_AGEMA_signal_2433) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L0), .B(SubCellInst_SboxInst_15_T3), .Z(
        SubCellOutput[60]) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2346), .B(new_AGEMA_signal_2280), .Z(new_AGEMA_signal_2434) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR10_U1_Ins_2_U1 ( .A(new_AGEMA_signal_2347), .B(new_AGEMA_signal_2281), .Z(new_AGEMA_signal_2435) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR_o1_U1_Ins0_U1 ( .A(
        new_AGEMA_signal_4913), .B(SubCellInst_SboxInst_15_YY_3), .ZN(
        SubCellOutput[61]) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_4915), .B(new_AGEMA_signal_2432), .Z(
        new_AGEMA_signal_2518) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_o1_U1_Ins_2_U1 ( .A(
        new_AGEMA_signal_4917), .B(new_AGEMA_signal_2433), .Z(
        new_AGEMA_signal_2519) );
  INV_X1 AddConstXOR_U2_U1 ( .A(SubCellOutput_29), .ZN(ShiftRowsOutput[21]) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_0_n1), .B(new_AGEMA_signal_4921), 
        .ZN(AddRoundConstantOutput[60]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2520), .B(1'b0), .Z(new_AGEMA_signal_2596) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2521), .B(1'b0), .Z(new_AGEMA_signal_2597) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[60]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_0_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2434), .Z(new_AGEMA_signal_2520) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2435), .Z(new_AGEMA_signal_2521) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_1_n1), .B(new_AGEMA_signal_4925), 
        .ZN(AddRoundConstantOutput[61]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2598), .B(1'b0), .Z(new_AGEMA_signal_2730) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2599), .B(1'b0), .Z(new_AGEMA_signal_2731) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[61]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_1_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2518), .Z(new_AGEMA_signal_2598) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2519), .Z(new_AGEMA_signal_2599) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_0_n1), .B(new_AGEMA_signal_4929), 
        .ZN(AddRoundConstantOutput[44]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2524), .B(1'b0), .Z(new_AGEMA_signal_2600) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2525), .B(1'b0), .Z(new_AGEMA_signal_2601) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_44), .ZN(AddConstXOR_AddConstXOR_XORInst_1_0_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2418), .Z(new_AGEMA_signal_2524) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2419), .Z(new_AGEMA_signal_2525) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_1_n1), .B(new_AGEMA_signal_4933), 
        .ZN(AddRoundConstantOutput[45]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2602), .B(1'b0), .Z(new_AGEMA_signal_2732) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2603), .B(1'b0), .Z(new_AGEMA_signal_2733) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_45), .ZN(AddConstXOR_AddConstXOR_XORInst_1_1_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2510), .Z(new_AGEMA_signal_2602) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2511), .Z(new_AGEMA_signal_2603) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_0_n1), .B(new_AGEMA_signal_4937), .ZN(
        ShiftRowsOutput[44]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2528), .B(new_AGEMA_signal_4941), .Z(
        new_AGEMA_signal_2604) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2529), .B(new_AGEMA_signal_4945), .Z(
        new_AGEMA_signal_2605) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[32]), .ZN(AddRoundTweakeyXOR_XORInst_0_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2406), .Z(new_AGEMA_signal_2528) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2407), .Z(new_AGEMA_signal_2529) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_1_n1), .B(new_AGEMA_signal_4949), .ZN(
        ShiftRowsOutput[45]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2606), .B(new_AGEMA_signal_4953), .Z(
        new_AGEMA_signal_2734) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2607), .B(new_AGEMA_signal_4957), .Z(
        new_AGEMA_signal_2735) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[33]), .ZN(AddRoundTweakeyXOR_XORInst_0_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2504), .Z(new_AGEMA_signal_2606) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2505), .Z(new_AGEMA_signal_2607) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_0_n1), .B(new_AGEMA_signal_4961), .ZN(
        ShiftRowsOutput[32]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2532), .B(new_AGEMA_signal_4965), .Z(
        new_AGEMA_signal_2608) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2533), .B(new_AGEMA_signal_4969), .Z(
        new_AGEMA_signal_2609) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[36]), .ZN(AddRoundTweakeyXOR_XORInst_1_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2410), .Z(new_AGEMA_signal_2532) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2411), .Z(new_AGEMA_signal_2533) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_1_n1), .B(new_AGEMA_signal_4973), .ZN(
        ShiftRowsOutput[33]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2610), .B(new_AGEMA_signal_4977), .Z(
        new_AGEMA_signal_2736) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2611), .B(new_AGEMA_signal_4981), .Z(
        new_AGEMA_signal_2737) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[37]), .ZN(AddRoundTweakeyXOR_XORInst_1_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2506), .Z(new_AGEMA_signal_2610) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2507), .Z(new_AGEMA_signal_2611) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_0_n1), .B(new_AGEMA_signal_4985), .ZN(
        ShiftRowsOutput[36]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2536), .B(new_AGEMA_signal_4989), .Z(
        new_AGEMA_signal_2612) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2537), .B(new_AGEMA_signal_4993), .Z(
        new_AGEMA_signal_2613) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[40]), .ZN(AddRoundTweakeyXOR_XORInst_2_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2414), .Z(new_AGEMA_signal_2536) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2415), .Z(new_AGEMA_signal_2537) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_1_n1), .B(new_AGEMA_signal_4997), .ZN(
        ShiftRowsOutput[37]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2614), .B(new_AGEMA_signal_5001), .Z(
        new_AGEMA_signal_2738) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2615), .B(new_AGEMA_signal_5005), .Z(
        new_AGEMA_signal_2739) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[41]), .ZN(AddRoundTweakeyXOR_XORInst_2_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2508), .Z(new_AGEMA_signal_2614) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2509), .Z(new_AGEMA_signal_2615) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_0_n1), .B(new_AGEMA_signal_5009), .ZN(
        ShiftRowsOutput[40]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2740), .B(new_AGEMA_signal_5013), .Z(
        new_AGEMA_signal_2850) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2741), .B(new_AGEMA_signal_5017), .Z(
        new_AGEMA_signal_2851) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[44]), .ZN(AddRoundTweakeyXOR_XORInst_3_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2600), .Z(new_AGEMA_signal_2740) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2601), .Z(new_AGEMA_signal_2741) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_1_n1), .B(new_AGEMA_signal_5021), .ZN(
        ShiftRowsOutput[41]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2852), .B(new_AGEMA_signal_5025), .Z(
        new_AGEMA_signal_2958) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2853), .B(new_AGEMA_signal_5029), .Z(
        new_AGEMA_signal_2959) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[45]), .ZN(AddRoundTweakeyXOR_XORInst_3_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2732), .Z(new_AGEMA_signal_2852) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2733), .Z(new_AGEMA_signal_2853) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_0_n1), .B(new_AGEMA_signal_5033), .ZN(
        MCOutput[32]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2542), .B(new_AGEMA_signal_5037), .Z(
        new_AGEMA_signal_2620) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2543), .B(new_AGEMA_signal_5041), .Z(
        new_AGEMA_signal_2621) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[48]), .ZN(AddRoundTweakeyXOR_XORInst_4_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2422), .Z(new_AGEMA_signal_2542) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2423), .Z(new_AGEMA_signal_2543) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_1_n1), .B(new_AGEMA_signal_5045), .ZN(
        MCOutput[33]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2622), .B(new_AGEMA_signal_5049), .Z(
        new_AGEMA_signal_2744) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2623), .B(new_AGEMA_signal_5053), .Z(
        new_AGEMA_signal_2745) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[49]), .ZN(AddRoundTweakeyXOR_XORInst_4_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2512), .Z(new_AGEMA_signal_2622) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2513), .Z(new_AGEMA_signal_2623) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_0_n1), .B(new_AGEMA_signal_5057), .ZN(
        MCOutput[36]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2546), .B(new_AGEMA_signal_5061), .Z(
        new_AGEMA_signal_2624) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2547), .B(new_AGEMA_signal_5065), .Z(
        new_AGEMA_signal_2625) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[52]), .ZN(AddRoundTweakeyXOR_XORInst_5_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2426), .Z(new_AGEMA_signal_2546) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2427), .Z(new_AGEMA_signal_2547) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_1_n1), .B(new_AGEMA_signal_5069), .ZN(
        MCOutput[37]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2626), .B(new_AGEMA_signal_5073), .Z(
        new_AGEMA_signal_2746) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2627), .B(new_AGEMA_signal_5077), .Z(
        new_AGEMA_signal_2747) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[53]), .ZN(AddRoundTweakeyXOR_XORInst_5_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2514), .Z(new_AGEMA_signal_2626) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2515), .Z(new_AGEMA_signal_2627) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_0_n1), .B(new_AGEMA_signal_5081), .ZN(
        MCOutput[40]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2550), .B(new_AGEMA_signal_5085), .Z(
        new_AGEMA_signal_2628) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2551), .B(new_AGEMA_signal_5089), .Z(
        new_AGEMA_signal_2629) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[56]), .ZN(AddRoundTweakeyXOR_XORInst_6_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2430), .Z(new_AGEMA_signal_2550) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2431), .Z(new_AGEMA_signal_2551) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_1_n1), .B(new_AGEMA_signal_5093), .ZN(
        MCOutput[41]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2630), .B(new_AGEMA_signal_5097), .Z(
        new_AGEMA_signal_2748) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2631), .B(new_AGEMA_signal_5101), .Z(
        new_AGEMA_signal_2749) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[57]), .ZN(AddRoundTweakeyXOR_XORInst_6_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2516), .Z(new_AGEMA_signal_2630) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2517), .Z(new_AGEMA_signal_2631) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_0_n1), .B(new_AGEMA_signal_5105), .ZN(
        MCOutput[44]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2750), .B(new_AGEMA_signal_5109), .Z(
        new_AGEMA_signal_2854) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2751), .B(new_AGEMA_signal_5113), .Z(
        new_AGEMA_signal_2855) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[60]), .ZN(AddRoundTweakeyXOR_XORInst_7_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2596), .Z(new_AGEMA_signal_2750) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2597), .Z(new_AGEMA_signal_2751) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_1_n1), .B(new_AGEMA_signal_5117), .ZN(
        MCOutput[45]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2856), .B(new_AGEMA_signal_5121), .Z(
        new_AGEMA_signal_2960) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U2_Ins_2_U1 ( .A(
        new_AGEMA_signal_2857), .B(new_AGEMA_signal_5125), .Z(
        new_AGEMA_signal_2961) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[61]), .ZN(AddRoundTweakeyXOR_XORInst_7_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2730), .Z(new_AGEMA_signal_2856) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2731), .Z(new_AGEMA_signal_2857) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_0_n2), 
        .B(MCInst_MCR0_XORInst_0_0_n1), .ZN(MCOutput[48]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2754), .B(
        new_AGEMA_signal_2556), .Z(new_AGEMA_signal_2858) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2755), .B(
        new_AGEMA_signal_2557), .Z(new_AGEMA_signal_2859) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[16]), .B(
        ShiftRowsOutput[0]), .ZN(MCInst_MCR0_XORInst_0_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2398), .B(
        new_AGEMA_signal_2386), .Z(new_AGEMA_signal_2556) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2399), .B(
        new_AGEMA_signal_2387), .Z(new_AGEMA_signal_2557) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[32]), 
        .Z(MCInst_MCR0_XORInst_0_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2620), .Z(new_AGEMA_signal_2754) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2621), .Z(new_AGEMA_signal_2755) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_1_n2), 
        .B(MCInst_MCR0_XORInst_0_1_n1), .ZN(MCOutput[49]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2860), .B(
        new_AGEMA_signal_2636), .Z(new_AGEMA_signal_2962) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2861), .B(
        new_AGEMA_signal_2637), .Z(new_AGEMA_signal_2963) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[17]), .B(
        ShiftRowsOutput[1]), .ZN(MCInst_MCR0_XORInst_0_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2500), .B(
        new_AGEMA_signal_2494), .Z(new_AGEMA_signal_2636) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2501), .B(
        new_AGEMA_signal_2495), .Z(new_AGEMA_signal_2637) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[33]), 
        .Z(MCInst_MCR0_XORInst_0_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2744), .Z(new_AGEMA_signal_2860) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2745), .Z(new_AGEMA_signal_2861) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_0_n2), 
        .B(MCInst_MCR0_XORInst_1_0_n1), .ZN(MCOutput[52]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2758), .B(
        new_AGEMA_signal_2560), .Z(new_AGEMA_signal_2862) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2759), .B(
        new_AGEMA_signal_2561), .Z(new_AGEMA_signal_2863) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[20]), .B(
        ShiftRowsOutput[4]), .ZN(MCInst_MCR0_XORInst_1_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2402), .B(
        new_AGEMA_signal_2374), .Z(new_AGEMA_signal_2560) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2403), .B(
        new_AGEMA_signal_2375), .Z(new_AGEMA_signal_2561) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[36]), 
        .Z(MCInst_MCR0_XORInst_1_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2624), .Z(new_AGEMA_signal_2758) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2625), .Z(new_AGEMA_signal_2759) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_1_n2), 
        .B(MCInst_MCR0_XORInst_1_1_n1), .ZN(MCOutput[53]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2864), .B(
        new_AGEMA_signal_2760), .Z(new_AGEMA_signal_2964) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2865), .B(
        new_AGEMA_signal_2761), .Z(new_AGEMA_signal_2965) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[21]), .B(
        ShiftRowsOutput[5]), .ZN(MCInst_MCR0_XORInst_1_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2594), .B(
        new_AGEMA_signal_2488), .Z(new_AGEMA_signal_2760) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2595), .B(
        new_AGEMA_signal_2489), .Z(new_AGEMA_signal_2761) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[37]), 
        .Z(MCInst_MCR0_XORInst_1_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2746), .Z(new_AGEMA_signal_2864) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2747), .Z(new_AGEMA_signal_2865) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_0_n2), 
        .B(MCInst_MCR0_XORInst_2_0_n1), .ZN(MCOutput[56]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2764), .B(
        new_AGEMA_signal_2564), .Z(new_AGEMA_signal_2866) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2765), .B(
        new_AGEMA_signal_2565), .Z(new_AGEMA_signal_2867) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[24]), .B(
        ShiftRowsOutput[8]), .ZN(MCInst_MCR0_XORInst_2_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2390), .B(
        new_AGEMA_signal_2378), .Z(new_AGEMA_signal_2564) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2391), .B(
        new_AGEMA_signal_2379), .Z(new_AGEMA_signal_2565) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[40]), 
        .Z(MCInst_MCR0_XORInst_2_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2628), .Z(new_AGEMA_signal_2764) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2629), .Z(new_AGEMA_signal_2765) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_1_n2), 
        .B(MCInst_MCR0_XORInst_2_1_n1), .ZN(MCOutput[57]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2868), .B(
        new_AGEMA_signal_2646), .Z(new_AGEMA_signal_2966) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2869), .B(
        new_AGEMA_signal_2647), .Z(new_AGEMA_signal_2967) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[25]), .B(
        ShiftRowsOutput[9]), .ZN(MCInst_MCR0_XORInst_2_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2496), .B(
        new_AGEMA_signal_2490), .Z(new_AGEMA_signal_2646) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2497), .B(
        new_AGEMA_signal_2491), .Z(new_AGEMA_signal_2647) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[41]), 
        .Z(MCInst_MCR0_XORInst_2_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2748), .Z(new_AGEMA_signal_2868) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2749), .Z(new_AGEMA_signal_2869) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_0_n2), 
        .B(MCInst_MCR0_XORInst_3_0_n1), .ZN(MCOutput[60]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2968), .B(
        new_AGEMA_signal_2568), .Z(new_AGEMA_signal_3044) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U3_Ins_2_U1 ( .A(new_AGEMA_signal_2969), .B(
        new_AGEMA_signal_2569), .Z(new_AGEMA_signal_3045) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[28]), .B(
        ShiftRowsOutput[12]), .ZN(MCInst_MCR0_XORInst_3_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2394), .B(
        new_AGEMA_signal_2382), .Z(new_AGEMA_signal_2568) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2395), .B(
        new_AGEMA_signal_2383), .Z(new_AGEMA_signal_2569) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[44]), 
        .Z(MCInst_MCR0_XORInst_3_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2854), .Z(new_AGEMA_signal_2968) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2855), .Z(new_AGEMA_signal_2969) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_1_n2), 
        .B(MCInst_MCR0_XORInst_3_1_n1), .ZN(MCOutput[61]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_3046), .B(
        new_AGEMA_signal_2652), .Z(new_AGEMA_signal_3068) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U3_Ins_2_U1 ( .A(new_AGEMA_signal_3047), .B(
        new_AGEMA_signal_2653), .Z(new_AGEMA_signal_3069) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[29]), .B(
        ShiftRowsOutput[13]), .ZN(MCInst_MCR0_XORInst_3_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2498), .B(
        new_AGEMA_signal_2492), .Z(new_AGEMA_signal_2652) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2499), .B(
        new_AGEMA_signal_2493), .Z(new_AGEMA_signal_2653) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[45]), 
        .Z(MCInst_MCR0_XORInst_3_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2960), .Z(new_AGEMA_signal_3046) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2961), .Z(new_AGEMA_signal_3047) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_0_n1), 
        .B(ShiftRowsOutput[16]), .ZN(MCOutput[16]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2770), .B(
        new_AGEMA_signal_2398), .Z(new_AGEMA_signal_2874) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2771), .B(
        new_AGEMA_signal_2399), .Z(new_AGEMA_signal_2875) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[32]), .ZN(MCInst_MCR2_XORInst_0_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2608), .Z(new_AGEMA_signal_2770) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2609), .Z(new_AGEMA_signal_2771) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_1_n1), 
        .B(ShiftRowsOutput[17]), .ZN(MCOutput[17]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2876), .B(
        new_AGEMA_signal_2500), .Z(new_AGEMA_signal_2972) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2877), .B(
        new_AGEMA_signal_2501), .Z(new_AGEMA_signal_2973) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[33]), .ZN(MCInst_MCR2_XORInst_0_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2736), .Z(new_AGEMA_signal_2876) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2737), .Z(new_AGEMA_signal_2877) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_0_n1), 
        .B(ShiftRowsOutput[20]), .ZN(MCOutput[20]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2774), .B(
        new_AGEMA_signal_2402), .Z(new_AGEMA_signal_2878) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2775), .B(
        new_AGEMA_signal_2403), .Z(new_AGEMA_signal_2879) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[36]), .ZN(MCInst_MCR2_XORInst_1_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2612), .Z(new_AGEMA_signal_2774) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2613), .Z(new_AGEMA_signal_2775) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_1_n1), 
        .B(ShiftRowsOutput[21]), .ZN(MCOutput[21]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2880), .B(
        new_AGEMA_signal_2594), .Z(new_AGEMA_signal_2974) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2881), .B(
        new_AGEMA_signal_2595), .Z(new_AGEMA_signal_2975) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[37]), .ZN(MCInst_MCR2_XORInst_1_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2738), .Z(new_AGEMA_signal_2880) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2739), .Z(new_AGEMA_signal_2881) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_0_n1), 
        .B(ShiftRowsOutput[24]), .ZN(MCOutput[24]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2976), .B(
        new_AGEMA_signal_2390), .Z(new_AGEMA_signal_3048) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2977), .B(
        new_AGEMA_signal_2391), .Z(new_AGEMA_signal_3049) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[40]), .ZN(MCInst_MCR2_XORInst_2_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2850), .Z(new_AGEMA_signal_2976) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2851), .Z(new_AGEMA_signal_2977) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_1_n1), 
        .B(ShiftRowsOutput[25]), .ZN(MCOutput[25]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3050), .B(
        new_AGEMA_signal_2496), .Z(new_AGEMA_signal_3070) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3051), .B(
        new_AGEMA_signal_2497), .Z(new_AGEMA_signal_3071) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[41]), .ZN(MCInst_MCR2_XORInst_2_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2958), .Z(new_AGEMA_signal_3050) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2959), .Z(new_AGEMA_signal_3051) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_0_n1), 
        .B(ShiftRowsOutput[28]), .ZN(MCOutput[28]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2780), .B(
        new_AGEMA_signal_2394), .Z(new_AGEMA_signal_2886) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2781), .B(
        new_AGEMA_signal_2395), .Z(new_AGEMA_signal_2887) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[44]), .ZN(MCInst_MCR2_XORInst_3_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2604), .Z(new_AGEMA_signal_2780) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2605), .Z(new_AGEMA_signal_2781) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_1_n1), 
        .B(ShiftRowsOutput[29]), .ZN(MCOutput[29]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2888), .B(
        new_AGEMA_signal_2498), .Z(new_AGEMA_signal_2980) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2889), .B(
        new_AGEMA_signal_2499), .Z(new_AGEMA_signal_2981) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[45]), .ZN(MCInst_MCR2_XORInst_3_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2734), .Z(new_AGEMA_signal_2888) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2735), .Z(new_AGEMA_signal_2889) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_0_n1), 
        .B(ShiftRowsOutput[16]), .ZN(MCOutput[0]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2784), .B(
        new_AGEMA_signal_2398), .Z(new_AGEMA_signal_2890) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2785), .B(
        new_AGEMA_signal_2399), .Z(new_AGEMA_signal_2891) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[32]), 
        .ZN(MCInst_MCR3_XORInst_0_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2620), .Z(new_AGEMA_signal_2784) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2621), .Z(new_AGEMA_signal_2785) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_1_n1), 
        .B(ShiftRowsOutput[17]), .ZN(MCOutput[1]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2892), .B(
        new_AGEMA_signal_2500), .Z(new_AGEMA_signal_2982) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2893), .B(
        new_AGEMA_signal_2501), .Z(new_AGEMA_signal_2983) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[33]), 
        .ZN(MCInst_MCR3_XORInst_0_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2744), .Z(new_AGEMA_signal_2892) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2745), .Z(new_AGEMA_signal_2893) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_0_n1), 
        .B(ShiftRowsOutput[20]), .ZN(MCOutput[4]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2788), .B(
        new_AGEMA_signal_2402), .Z(new_AGEMA_signal_2894) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2789), .B(
        new_AGEMA_signal_2403), .Z(new_AGEMA_signal_2895) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[36]), 
        .ZN(MCInst_MCR3_XORInst_1_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2624), .Z(new_AGEMA_signal_2788) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2625), .Z(new_AGEMA_signal_2789) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_1_n1), 
        .B(ShiftRowsOutput[21]), .ZN(MCOutput[5]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2896), .B(
        new_AGEMA_signal_2594), .Z(new_AGEMA_signal_2984) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2897), .B(
        new_AGEMA_signal_2595), .Z(new_AGEMA_signal_2985) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[37]), 
        .ZN(MCInst_MCR3_XORInst_1_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2746), .Z(new_AGEMA_signal_2896) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2747), .Z(new_AGEMA_signal_2897) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_0_n1), 
        .B(ShiftRowsOutput[24]), .ZN(MCOutput[8]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2792), .B(
        new_AGEMA_signal_2390), .Z(new_AGEMA_signal_2898) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2793), .B(
        new_AGEMA_signal_2391), .Z(new_AGEMA_signal_2899) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[40]), 
        .ZN(MCInst_MCR3_XORInst_2_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2628), .Z(new_AGEMA_signal_2792) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2629), .Z(new_AGEMA_signal_2793) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_1_n1), 
        .B(ShiftRowsOutput[25]), .ZN(MCOutput[9]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2900), .B(
        new_AGEMA_signal_2496), .Z(new_AGEMA_signal_2986) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2901), .B(
        new_AGEMA_signal_2497), .Z(new_AGEMA_signal_2987) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[41]), 
        .ZN(MCInst_MCR3_XORInst_2_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2748), .Z(new_AGEMA_signal_2900) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2749), .Z(new_AGEMA_signal_2901) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_0_n1), 
        .B(ShiftRowsOutput[28]), .ZN(MCOutput[12]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2988), .B(
        new_AGEMA_signal_2394), .Z(new_AGEMA_signal_3052) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U2_Ins_2_U1 ( .A(new_AGEMA_signal_2989), .B(
        new_AGEMA_signal_2395), .Z(new_AGEMA_signal_3053) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[44]), 
        .ZN(MCInst_MCR3_XORInst_3_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2854), .Z(new_AGEMA_signal_2988) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2855), .Z(new_AGEMA_signal_2989) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_1_n1), 
        .B(ShiftRowsOutput[29]), .ZN(MCOutput[13]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_3054), .B(
        new_AGEMA_signal_2498), .Z(new_AGEMA_signal_3072) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U2_Ins_2_U1 ( .A(new_AGEMA_signal_3055), .B(
        new_AGEMA_signal_2499), .Z(new_AGEMA_signal_3073) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[45]), 
        .ZN(MCInst_MCR3_XORInst_3_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2960), .Z(new_AGEMA_signal_3054) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U1_Ins_2_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2961), .Z(new_AGEMA_signal_3055) );
  DFF_X1 new_AGEMA_reg_buffer_1679_s_current_state_reg ( .D(
        new_AGEMA_signal_3956), .CK(clk), .Q(new_AGEMA_signal_3957), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1683_s_current_state_reg ( .D(
        new_AGEMA_signal_3960), .CK(clk), .Q(new_AGEMA_signal_3961), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1687_s_current_state_reg ( .D(
        new_AGEMA_signal_3964), .CK(clk), .Q(new_AGEMA_signal_3965), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1691_s_current_state_reg ( .D(
        new_AGEMA_signal_3968), .CK(clk), .Q(new_AGEMA_signal_3969), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1695_s_current_state_reg ( .D(
        new_AGEMA_signal_3972), .CK(clk), .Q(new_AGEMA_signal_3973), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1699_s_current_state_reg ( .D(
        new_AGEMA_signal_3976), .CK(clk), .Q(new_AGEMA_signal_3977), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1703_s_current_state_reg ( .D(
        new_AGEMA_signal_3980), .CK(clk), .Q(new_AGEMA_signal_3981), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1707_s_current_state_reg ( .D(
        new_AGEMA_signal_3984), .CK(clk), .Q(new_AGEMA_signal_3985), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1711_s_current_state_reg ( .D(
        new_AGEMA_signal_3988), .CK(clk), .Q(new_AGEMA_signal_3989), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1715_s_current_state_reg ( .D(
        new_AGEMA_signal_3992), .CK(clk), .Q(new_AGEMA_signal_3993), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1719_s_current_state_reg ( .D(
        new_AGEMA_signal_3996), .CK(clk), .Q(new_AGEMA_signal_3997), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1723_s_current_state_reg ( .D(
        new_AGEMA_signal_4000), .CK(clk), .Q(new_AGEMA_signal_4001), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1727_s_current_state_reg ( .D(
        new_AGEMA_signal_4004), .CK(clk), .Q(new_AGEMA_signal_4005), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1731_s_current_state_reg ( .D(
        new_AGEMA_signal_4008), .CK(clk), .Q(new_AGEMA_signal_4009), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1735_s_current_state_reg ( .D(
        new_AGEMA_signal_4012), .CK(clk), .Q(new_AGEMA_signal_4013), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1739_s_current_state_reg ( .D(
        new_AGEMA_signal_4016), .CK(clk), .Q(new_AGEMA_signal_4017), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1743_s_current_state_reg ( .D(
        new_AGEMA_signal_4020), .CK(clk), .Q(new_AGEMA_signal_4021), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1747_s_current_state_reg ( .D(
        new_AGEMA_signal_4024), .CK(clk), .Q(new_AGEMA_signal_4025), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1751_s_current_state_reg ( .D(
        new_AGEMA_signal_4028), .CK(clk), .Q(new_AGEMA_signal_4029), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1755_s_current_state_reg ( .D(
        new_AGEMA_signal_4032), .CK(clk), .Q(new_AGEMA_signal_4033), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1759_s_current_state_reg ( .D(
        new_AGEMA_signal_4036), .CK(clk), .Q(new_AGEMA_signal_4037), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1763_s_current_state_reg ( .D(
        new_AGEMA_signal_4040), .CK(clk), .Q(new_AGEMA_signal_4041), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1767_s_current_state_reg ( .D(
        new_AGEMA_signal_4044), .CK(clk), .Q(new_AGEMA_signal_4045), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1771_s_current_state_reg ( .D(
        new_AGEMA_signal_4048), .CK(clk), .Q(new_AGEMA_signal_4049), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1775_s_current_state_reg ( .D(
        new_AGEMA_signal_4052), .CK(clk), .Q(new_AGEMA_signal_4053), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1779_s_current_state_reg ( .D(
        new_AGEMA_signal_4056), .CK(clk), .Q(new_AGEMA_signal_4057), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1783_s_current_state_reg ( .D(
        new_AGEMA_signal_4060), .CK(clk), .Q(new_AGEMA_signal_4061), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1787_s_current_state_reg ( .D(
        new_AGEMA_signal_4064), .CK(clk), .Q(new_AGEMA_signal_4065), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1791_s_current_state_reg ( .D(
        new_AGEMA_signal_4068), .CK(clk), .Q(new_AGEMA_signal_4069), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1795_s_current_state_reg ( .D(
        new_AGEMA_signal_4072), .CK(clk), .Q(new_AGEMA_signal_4073), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1799_s_current_state_reg ( .D(
        new_AGEMA_signal_4076), .CK(clk), .Q(new_AGEMA_signal_4077), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1803_s_current_state_reg ( .D(
        new_AGEMA_signal_4080), .CK(clk), .Q(new_AGEMA_signal_4081), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1807_s_current_state_reg ( .D(
        new_AGEMA_signal_4084), .CK(clk), .Q(new_AGEMA_signal_4085), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1811_s_current_state_reg ( .D(
        new_AGEMA_signal_4088), .CK(clk), .Q(new_AGEMA_signal_4089), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1815_s_current_state_reg ( .D(
        new_AGEMA_signal_4092), .CK(clk), .Q(new_AGEMA_signal_4093), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1819_s_current_state_reg ( .D(
        new_AGEMA_signal_4096), .CK(clk), .Q(new_AGEMA_signal_4097), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1823_s_current_state_reg ( .D(
        new_AGEMA_signal_4100), .CK(clk), .Q(new_AGEMA_signal_4101), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1827_s_current_state_reg ( .D(
        new_AGEMA_signal_4104), .CK(clk), .Q(new_AGEMA_signal_4105), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1831_s_current_state_reg ( .D(
        new_AGEMA_signal_4108), .CK(clk), .Q(new_AGEMA_signal_4109), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1835_s_current_state_reg ( .D(
        new_AGEMA_signal_4112), .CK(clk), .Q(new_AGEMA_signal_4113), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1839_s_current_state_reg ( .D(
        new_AGEMA_signal_4116), .CK(clk), .Q(new_AGEMA_signal_4117), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1843_s_current_state_reg ( .D(
        new_AGEMA_signal_4120), .CK(clk), .Q(new_AGEMA_signal_4121), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1847_s_current_state_reg ( .D(
        new_AGEMA_signal_4124), .CK(clk), .Q(new_AGEMA_signal_4125), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1851_s_current_state_reg ( .D(
        new_AGEMA_signal_4128), .CK(clk), .Q(new_AGEMA_signal_4129), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1855_s_current_state_reg ( .D(
        new_AGEMA_signal_4132), .CK(clk), .Q(new_AGEMA_signal_4133), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1859_s_current_state_reg ( .D(
        new_AGEMA_signal_4136), .CK(clk), .Q(new_AGEMA_signal_4137), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1863_s_current_state_reg ( .D(
        new_AGEMA_signal_4140), .CK(clk), .Q(new_AGEMA_signal_4141), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1867_s_current_state_reg ( .D(
        new_AGEMA_signal_4144), .CK(clk), .Q(new_AGEMA_signal_4145), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1871_s_current_state_reg ( .D(
        new_AGEMA_signal_4148), .CK(clk), .Q(new_AGEMA_signal_4149), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1875_s_current_state_reg ( .D(
        new_AGEMA_signal_4152), .CK(clk), .Q(new_AGEMA_signal_4153), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1879_s_current_state_reg ( .D(
        new_AGEMA_signal_4156), .CK(clk), .Q(new_AGEMA_signal_4157), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1883_s_current_state_reg ( .D(
        new_AGEMA_signal_4160), .CK(clk), .Q(new_AGEMA_signal_4161), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1887_s_current_state_reg ( .D(
        new_AGEMA_signal_4164), .CK(clk), .Q(new_AGEMA_signal_4165), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1891_s_current_state_reg ( .D(
        new_AGEMA_signal_4168), .CK(clk), .Q(new_AGEMA_signal_4169), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1895_s_current_state_reg ( .D(
        new_AGEMA_signal_4172), .CK(clk), .Q(new_AGEMA_signal_4173), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1899_s_current_state_reg ( .D(
        new_AGEMA_signal_4176), .CK(clk), .Q(new_AGEMA_signal_4177), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1903_s_current_state_reg ( .D(
        new_AGEMA_signal_4180), .CK(clk), .Q(new_AGEMA_signal_4181), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1907_s_current_state_reg ( .D(
        new_AGEMA_signal_4184), .CK(clk), .Q(new_AGEMA_signal_4185), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1911_s_current_state_reg ( .D(
        new_AGEMA_signal_4188), .CK(clk), .Q(new_AGEMA_signal_4189), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1915_s_current_state_reg ( .D(
        new_AGEMA_signal_4192), .CK(clk), .Q(new_AGEMA_signal_4193), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1919_s_current_state_reg ( .D(
        new_AGEMA_signal_4196), .CK(clk), .Q(new_AGEMA_signal_4197), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1923_s_current_state_reg ( .D(
        new_AGEMA_signal_4200), .CK(clk), .Q(new_AGEMA_signal_4201), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1927_s_current_state_reg ( .D(
        new_AGEMA_signal_4204), .CK(clk), .Q(new_AGEMA_signal_4205), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1931_s_current_state_reg ( .D(
        new_AGEMA_signal_4208), .CK(clk), .Q(new_AGEMA_signal_4209), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1935_s_current_state_reg ( .D(
        new_AGEMA_signal_4212), .CK(clk), .Q(new_AGEMA_signal_4213), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1939_s_current_state_reg ( .D(
        new_AGEMA_signal_4216), .CK(clk), .Q(new_AGEMA_signal_4217), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1943_s_current_state_reg ( .D(
        new_AGEMA_signal_4220), .CK(clk), .Q(new_AGEMA_signal_4221), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1947_s_current_state_reg ( .D(
        new_AGEMA_signal_4224), .CK(clk), .Q(new_AGEMA_signal_4225), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1951_s_current_state_reg ( .D(
        new_AGEMA_signal_4228), .CK(clk), .Q(new_AGEMA_signal_4229), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1955_s_current_state_reg ( .D(
        new_AGEMA_signal_4232), .CK(clk), .Q(new_AGEMA_signal_4233), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1959_s_current_state_reg ( .D(
        new_AGEMA_signal_4236), .CK(clk), .Q(new_AGEMA_signal_4237), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1963_s_current_state_reg ( .D(
        new_AGEMA_signal_4240), .CK(clk), .Q(new_AGEMA_signal_4241), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1967_s_current_state_reg ( .D(
        new_AGEMA_signal_4244), .CK(clk), .Q(new_AGEMA_signal_4245), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1971_s_current_state_reg ( .D(
        new_AGEMA_signal_4248), .CK(clk), .Q(new_AGEMA_signal_4249), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1975_s_current_state_reg ( .D(
        new_AGEMA_signal_4252), .CK(clk), .Q(new_AGEMA_signal_4253), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1979_s_current_state_reg ( .D(
        new_AGEMA_signal_4256), .CK(clk), .Q(new_AGEMA_signal_4257), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1983_s_current_state_reg ( .D(
        new_AGEMA_signal_4260), .CK(clk), .Q(new_AGEMA_signal_4261), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1987_s_current_state_reg ( .D(
        new_AGEMA_signal_4264), .CK(clk), .Q(new_AGEMA_signal_4265), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1991_s_current_state_reg ( .D(
        new_AGEMA_signal_4268), .CK(clk), .Q(new_AGEMA_signal_4269), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1995_s_current_state_reg ( .D(
        new_AGEMA_signal_4272), .CK(clk), .Q(new_AGEMA_signal_4273), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_1999_s_current_state_reg ( .D(
        new_AGEMA_signal_4276), .CK(clk), .Q(new_AGEMA_signal_4277), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2003_s_current_state_reg ( .D(
        new_AGEMA_signal_4280), .CK(clk), .Q(new_AGEMA_signal_4281), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2007_s_current_state_reg ( .D(
        new_AGEMA_signal_4284), .CK(clk), .Q(new_AGEMA_signal_4285), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2011_s_current_state_reg ( .D(
        new_AGEMA_signal_4288), .CK(clk), .Q(new_AGEMA_signal_4289), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2015_s_current_state_reg ( .D(
        new_AGEMA_signal_4292), .CK(clk), .Q(new_AGEMA_signal_4293), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2019_s_current_state_reg ( .D(
        new_AGEMA_signal_4296), .CK(clk), .Q(new_AGEMA_signal_4297), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2023_s_current_state_reg ( .D(
        new_AGEMA_signal_4300), .CK(clk), .Q(new_AGEMA_signal_4301), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2027_s_current_state_reg ( .D(
        new_AGEMA_signal_4304), .CK(clk), .Q(new_AGEMA_signal_4305), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2031_s_current_state_reg ( .D(
        new_AGEMA_signal_4308), .CK(clk), .Q(new_AGEMA_signal_4309), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2035_s_current_state_reg ( .D(
        new_AGEMA_signal_4312), .CK(clk), .Q(new_AGEMA_signal_4313), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2039_s_current_state_reg ( .D(
        new_AGEMA_signal_4316), .CK(clk), .Q(new_AGEMA_signal_4317), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2043_s_current_state_reg ( .D(
        new_AGEMA_signal_4320), .CK(clk), .Q(new_AGEMA_signal_4321), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2047_s_current_state_reg ( .D(
        new_AGEMA_signal_4324), .CK(clk), .Q(new_AGEMA_signal_4325), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2051_s_current_state_reg ( .D(
        new_AGEMA_signal_4328), .CK(clk), .Q(new_AGEMA_signal_4329), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2055_s_current_state_reg ( .D(
        new_AGEMA_signal_4332), .CK(clk), .Q(new_AGEMA_signal_4333), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2059_s_current_state_reg ( .D(
        new_AGEMA_signal_4336), .CK(clk), .Q(new_AGEMA_signal_4337), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2063_s_current_state_reg ( .D(
        new_AGEMA_signal_4340), .CK(clk), .Q(new_AGEMA_signal_4341), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2071_s_current_state_reg ( .D(
        new_AGEMA_signal_4348), .CK(clk), .Q(new_AGEMA_signal_4349), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2073_s_current_state_reg ( .D(
        new_AGEMA_signal_4350), .CK(clk), .Q(new_AGEMA_signal_4351), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2075_s_current_state_reg ( .D(
        new_AGEMA_signal_4352), .CK(clk), .Q(new_AGEMA_signal_4353), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2085_s_current_state_reg ( .D(
        new_AGEMA_signal_4362), .CK(clk), .Q(new_AGEMA_signal_4363), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2089_s_current_state_reg ( .D(
        new_AGEMA_signal_4366), .CK(clk), .Q(new_AGEMA_signal_4367), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2093_s_current_state_reg ( .D(
        new_AGEMA_signal_4370), .CK(clk), .Q(new_AGEMA_signal_4371), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2095_s_current_state_reg ( .D(
        new_AGEMA_signal_4372), .CK(clk), .Q(new_AGEMA_signal_4373), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2097_s_current_state_reg ( .D(
        new_AGEMA_signal_4374), .CK(clk), .Q(new_AGEMA_signal_4375), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2099_s_current_state_reg ( .D(
        new_AGEMA_signal_4376), .CK(clk), .Q(new_AGEMA_signal_4377), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2107_s_current_state_reg ( .D(
        new_AGEMA_signal_4384), .CK(clk), .Q(new_AGEMA_signal_4385), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2109_s_current_state_reg ( .D(
        new_AGEMA_signal_4386), .CK(clk), .Q(new_AGEMA_signal_4387), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2111_s_current_state_reg ( .D(
        new_AGEMA_signal_4388), .CK(clk), .Q(new_AGEMA_signal_4389), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2121_s_current_state_reg ( .D(
        new_AGEMA_signal_4398), .CK(clk), .Q(new_AGEMA_signal_4399), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2125_s_current_state_reg ( .D(
        new_AGEMA_signal_4402), .CK(clk), .Q(new_AGEMA_signal_4403), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2129_s_current_state_reg ( .D(
        new_AGEMA_signal_4406), .CK(clk), .Q(new_AGEMA_signal_4407), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2131_s_current_state_reg ( .D(
        new_AGEMA_signal_4408), .CK(clk), .Q(new_AGEMA_signal_4409), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2133_s_current_state_reg ( .D(
        new_AGEMA_signal_4410), .CK(clk), .Q(new_AGEMA_signal_4411), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2135_s_current_state_reg ( .D(
        new_AGEMA_signal_4412), .CK(clk), .Q(new_AGEMA_signal_4413), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2143_s_current_state_reg ( .D(
        new_AGEMA_signal_4420), .CK(clk), .Q(new_AGEMA_signal_4421), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2145_s_current_state_reg ( .D(
        new_AGEMA_signal_4422), .CK(clk), .Q(new_AGEMA_signal_4423), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2147_s_current_state_reg ( .D(
        new_AGEMA_signal_4424), .CK(clk), .Q(new_AGEMA_signal_4425), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2157_s_current_state_reg ( .D(
        new_AGEMA_signal_4434), .CK(clk), .Q(new_AGEMA_signal_4435), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2161_s_current_state_reg ( .D(
        new_AGEMA_signal_4438), .CK(clk), .Q(new_AGEMA_signal_4439), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2165_s_current_state_reg ( .D(
        new_AGEMA_signal_4442), .CK(clk), .Q(new_AGEMA_signal_4443), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2167_s_current_state_reg ( .D(
        new_AGEMA_signal_4444), .CK(clk), .Q(new_AGEMA_signal_4445), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2169_s_current_state_reg ( .D(
        new_AGEMA_signal_4446), .CK(clk), .Q(new_AGEMA_signal_4447), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2171_s_current_state_reg ( .D(
        new_AGEMA_signal_4448), .CK(clk), .Q(new_AGEMA_signal_4449), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2179_s_current_state_reg ( .D(
        new_AGEMA_signal_4456), .CK(clk), .Q(new_AGEMA_signal_4457), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2181_s_current_state_reg ( .D(
        new_AGEMA_signal_4458), .CK(clk), .Q(new_AGEMA_signal_4459), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2183_s_current_state_reg ( .D(
        new_AGEMA_signal_4460), .CK(clk), .Q(new_AGEMA_signal_4461), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2193_s_current_state_reg ( .D(
        new_AGEMA_signal_4470), .CK(clk), .Q(new_AGEMA_signal_4471), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2197_s_current_state_reg ( .D(
        new_AGEMA_signal_4474), .CK(clk), .Q(new_AGEMA_signal_4475), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2201_s_current_state_reg ( .D(
        new_AGEMA_signal_4478), .CK(clk), .Q(new_AGEMA_signal_4479), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2203_s_current_state_reg ( .D(
        new_AGEMA_signal_4480), .CK(clk), .Q(new_AGEMA_signal_4481), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2205_s_current_state_reg ( .D(
        new_AGEMA_signal_4482), .CK(clk), .Q(new_AGEMA_signal_4483), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2207_s_current_state_reg ( .D(
        new_AGEMA_signal_4484), .CK(clk), .Q(new_AGEMA_signal_4485), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2215_s_current_state_reg ( .D(
        new_AGEMA_signal_4492), .CK(clk), .Q(new_AGEMA_signal_4493), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2217_s_current_state_reg ( .D(
        new_AGEMA_signal_4494), .CK(clk), .Q(new_AGEMA_signal_4495), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2219_s_current_state_reg ( .D(
        new_AGEMA_signal_4496), .CK(clk), .Q(new_AGEMA_signal_4497), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2229_s_current_state_reg ( .D(
        new_AGEMA_signal_4506), .CK(clk), .Q(new_AGEMA_signal_4507), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2233_s_current_state_reg ( .D(
        new_AGEMA_signal_4510), .CK(clk), .Q(new_AGEMA_signal_4511), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2237_s_current_state_reg ( .D(
        new_AGEMA_signal_4514), .CK(clk), .Q(new_AGEMA_signal_4515), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2239_s_current_state_reg ( .D(
        new_AGEMA_signal_4516), .CK(clk), .Q(new_AGEMA_signal_4517), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2241_s_current_state_reg ( .D(
        new_AGEMA_signal_4518), .CK(clk), .Q(new_AGEMA_signal_4519), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2243_s_current_state_reg ( .D(
        new_AGEMA_signal_4520), .CK(clk), .Q(new_AGEMA_signal_4521), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2251_s_current_state_reg ( .D(
        new_AGEMA_signal_4528), .CK(clk), .Q(new_AGEMA_signal_4529), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2253_s_current_state_reg ( .D(
        new_AGEMA_signal_4530), .CK(clk), .Q(new_AGEMA_signal_4531), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2255_s_current_state_reg ( .D(
        new_AGEMA_signal_4532), .CK(clk), .Q(new_AGEMA_signal_4533), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2265_s_current_state_reg ( .D(
        new_AGEMA_signal_4542), .CK(clk), .Q(new_AGEMA_signal_4543), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2269_s_current_state_reg ( .D(
        new_AGEMA_signal_4546), .CK(clk), .Q(new_AGEMA_signal_4547), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2273_s_current_state_reg ( .D(
        new_AGEMA_signal_4550), .CK(clk), .Q(new_AGEMA_signal_4551), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2275_s_current_state_reg ( .D(
        new_AGEMA_signal_4552), .CK(clk), .Q(new_AGEMA_signal_4553), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2277_s_current_state_reg ( .D(
        new_AGEMA_signal_4554), .CK(clk), .Q(new_AGEMA_signal_4555), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2279_s_current_state_reg ( .D(
        new_AGEMA_signal_4556), .CK(clk), .Q(new_AGEMA_signal_4557), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2287_s_current_state_reg ( .D(
        new_AGEMA_signal_4564), .CK(clk), .Q(new_AGEMA_signal_4565), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2289_s_current_state_reg ( .D(
        new_AGEMA_signal_4566), .CK(clk), .Q(new_AGEMA_signal_4567), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2291_s_current_state_reg ( .D(
        new_AGEMA_signal_4568), .CK(clk), .Q(new_AGEMA_signal_4569), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2301_s_current_state_reg ( .D(
        new_AGEMA_signal_4578), .CK(clk), .Q(new_AGEMA_signal_4579), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2305_s_current_state_reg ( .D(
        new_AGEMA_signal_4582), .CK(clk), .Q(new_AGEMA_signal_4583), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2309_s_current_state_reg ( .D(
        new_AGEMA_signal_4586), .CK(clk), .Q(new_AGEMA_signal_4587), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2311_s_current_state_reg ( .D(
        new_AGEMA_signal_4588), .CK(clk), .Q(new_AGEMA_signal_4589), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2313_s_current_state_reg ( .D(
        new_AGEMA_signal_4590), .CK(clk), .Q(new_AGEMA_signal_4591), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2315_s_current_state_reg ( .D(
        new_AGEMA_signal_4592), .CK(clk), .Q(new_AGEMA_signal_4593), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2323_s_current_state_reg ( .D(
        new_AGEMA_signal_4600), .CK(clk), .Q(new_AGEMA_signal_4601), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2325_s_current_state_reg ( .D(
        new_AGEMA_signal_4602), .CK(clk), .Q(new_AGEMA_signal_4603), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2327_s_current_state_reg ( .D(
        new_AGEMA_signal_4604), .CK(clk), .Q(new_AGEMA_signal_4605), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2337_s_current_state_reg ( .D(
        new_AGEMA_signal_4614), .CK(clk), .Q(new_AGEMA_signal_4615), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2341_s_current_state_reg ( .D(
        new_AGEMA_signal_4618), .CK(clk), .Q(new_AGEMA_signal_4619), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2345_s_current_state_reg ( .D(
        new_AGEMA_signal_4622), .CK(clk), .Q(new_AGEMA_signal_4623), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2347_s_current_state_reg ( .D(
        new_AGEMA_signal_4624), .CK(clk), .Q(new_AGEMA_signal_4625), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2349_s_current_state_reg ( .D(
        new_AGEMA_signal_4626), .CK(clk), .Q(new_AGEMA_signal_4627), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2351_s_current_state_reg ( .D(
        new_AGEMA_signal_4628), .CK(clk), .Q(new_AGEMA_signal_4629), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2359_s_current_state_reg ( .D(
        new_AGEMA_signal_4636), .CK(clk), .Q(new_AGEMA_signal_4637), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2361_s_current_state_reg ( .D(
        new_AGEMA_signal_4638), .CK(clk), .Q(new_AGEMA_signal_4639), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2363_s_current_state_reg ( .D(
        new_AGEMA_signal_4640), .CK(clk), .Q(new_AGEMA_signal_4641), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2373_s_current_state_reg ( .D(
        new_AGEMA_signal_4650), .CK(clk), .Q(new_AGEMA_signal_4651), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2377_s_current_state_reg ( .D(
        new_AGEMA_signal_4654), .CK(clk), .Q(new_AGEMA_signal_4655), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2381_s_current_state_reg ( .D(
        new_AGEMA_signal_4658), .CK(clk), .Q(new_AGEMA_signal_4659), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2383_s_current_state_reg ( .D(
        new_AGEMA_signal_4660), .CK(clk), .Q(new_AGEMA_signal_4661), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2385_s_current_state_reg ( .D(
        new_AGEMA_signal_4662), .CK(clk), .Q(new_AGEMA_signal_4663), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2387_s_current_state_reg ( .D(
        new_AGEMA_signal_4664), .CK(clk), .Q(new_AGEMA_signal_4665), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2395_s_current_state_reg ( .D(
        new_AGEMA_signal_4672), .CK(clk), .Q(new_AGEMA_signal_4673), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2397_s_current_state_reg ( .D(
        new_AGEMA_signal_4674), .CK(clk), .Q(new_AGEMA_signal_4675), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2399_s_current_state_reg ( .D(
        new_AGEMA_signal_4676), .CK(clk), .Q(new_AGEMA_signal_4677), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2409_s_current_state_reg ( .D(
        new_AGEMA_signal_4686), .CK(clk), .Q(new_AGEMA_signal_4687), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2413_s_current_state_reg ( .D(
        new_AGEMA_signal_4690), .CK(clk), .Q(new_AGEMA_signal_4691), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2417_s_current_state_reg ( .D(
        new_AGEMA_signal_4694), .CK(clk), .Q(new_AGEMA_signal_4695), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2419_s_current_state_reg ( .D(
        new_AGEMA_signal_4696), .CK(clk), .Q(new_AGEMA_signal_4697), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2421_s_current_state_reg ( .D(
        new_AGEMA_signal_4698), .CK(clk), .Q(new_AGEMA_signal_4699), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2423_s_current_state_reg ( .D(
        new_AGEMA_signal_4700), .CK(clk), .Q(new_AGEMA_signal_4701), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2431_s_current_state_reg ( .D(
        new_AGEMA_signal_4708), .CK(clk), .Q(new_AGEMA_signal_4709), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2433_s_current_state_reg ( .D(
        new_AGEMA_signal_4710), .CK(clk), .Q(new_AGEMA_signal_4711), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2435_s_current_state_reg ( .D(
        new_AGEMA_signal_4712), .CK(clk), .Q(new_AGEMA_signal_4713), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2445_s_current_state_reg ( .D(
        new_AGEMA_signal_4722), .CK(clk), .Q(new_AGEMA_signal_4723), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2449_s_current_state_reg ( .D(
        new_AGEMA_signal_4726), .CK(clk), .Q(new_AGEMA_signal_4727), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2453_s_current_state_reg ( .D(
        new_AGEMA_signal_4730), .CK(clk), .Q(new_AGEMA_signal_4731), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2455_s_current_state_reg ( .D(
        new_AGEMA_signal_4732), .CK(clk), .Q(new_AGEMA_signal_4733), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2457_s_current_state_reg ( .D(
        new_AGEMA_signal_4734), .CK(clk), .Q(new_AGEMA_signal_4735), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2459_s_current_state_reg ( .D(
        new_AGEMA_signal_4736), .CK(clk), .Q(new_AGEMA_signal_4737), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2467_s_current_state_reg ( .D(
        new_AGEMA_signal_4744), .CK(clk), .Q(new_AGEMA_signal_4745), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2469_s_current_state_reg ( .D(
        new_AGEMA_signal_4746), .CK(clk), .Q(new_AGEMA_signal_4747), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2471_s_current_state_reg ( .D(
        new_AGEMA_signal_4748), .CK(clk), .Q(new_AGEMA_signal_4749), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2481_s_current_state_reg ( .D(
        new_AGEMA_signal_4758), .CK(clk), .Q(new_AGEMA_signal_4759), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2485_s_current_state_reg ( .D(
        new_AGEMA_signal_4762), .CK(clk), .Q(new_AGEMA_signal_4763), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2489_s_current_state_reg ( .D(
        new_AGEMA_signal_4766), .CK(clk), .Q(new_AGEMA_signal_4767), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2491_s_current_state_reg ( .D(
        new_AGEMA_signal_4768), .CK(clk), .Q(new_AGEMA_signal_4769), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2493_s_current_state_reg ( .D(
        new_AGEMA_signal_4770), .CK(clk), .Q(new_AGEMA_signal_4771), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2495_s_current_state_reg ( .D(
        new_AGEMA_signal_4772), .CK(clk), .Q(new_AGEMA_signal_4773), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2503_s_current_state_reg ( .D(
        new_AGEMA_signal_4780), .CK(clk), .Q(new_AGEMA_signal_4781), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2505_s_current_state_reg ( .D(
        new_AGEMA_signal_4782), .CK(clk), .Q(new_AGEMA_signal_4783), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2507_s_current_state_reg ( .D(
        new_AGEMA_signal_4784), .CK(clk), .Q(new_AGEMA_signal_4785), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2517_s_current_state_reg ( .D(
        new_AGEMA_signal_4794), .CK(clk), .Q(new_AGEMA_signal_4795), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2521_s_current_state_reg ( .D(
        new_AGEMA_signal_4798), .CK(clk), .Q(new_AGEMA_signal_4799), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2525_s_current_state_reg ( .D(
        new_AGEMA_signal_4802), .CK(clk), .Q(new_AGEMA_signal_4803), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2527_s_current_state_reg ( .D(
        new_AGEMA_signal_4804), .CK(clk), .Q(new_AGEMA_signal_4805), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2529_s_current_state_reg ( .D(
        new_AGEMA_signal_4806), .CK(clk), .Q(new_AGEMA_signal_4807), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2531_s_current_state_reg ( .D(
        new_AGEMA_signal_4808), .CK(clk), .Q(new_AGEMA_signal_4809), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2539_s_current_state_reg ( .D(
        new_AGEMA_signal_4816), .CK(clk), .Q(new_AGEMA_signal_4817), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2541_s_current_state_reg ( .D(
        new_AGEMA_signal_4818), .CK(clk), .Q(new_AGEMA_signal_4819), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2543_s_current_state_reg ( .D(
        new_AGEMA_signal_4820), .CK(clk), .Q(new_AGEMA_signal_4821), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2553_s_current_state_reg ( .D(
        new_AGEMA_signal_4830), .CK(clk), .Q(new_AGEMA_signal_4831), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2557_s_current_state_reg ( .D(
        new_AGEMA_signal_4834), .CK(clk), .Q(new_AGEMA_signal_4835), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2561_s_current_state_reg ( .D(
        new_AGEMA_signal_4838), .CK(clk), .Q(new_AGEMA_signal_4839), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2563_s_current_state_reg ( .D(
        new_AGEMA_signal_4840), .CK(clk), .Q(new_AGEMA_signal_4841), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2565_s_current_state_reg ( .D(
        new_AGEMA_signal_4842), .CK(clk), .Q(new_AGEMA_signal_4843), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2567_s_current_state_reg ( .D(
        new_AGEMA_signal_4844), .CK(clk), .Q(new_AGEMA_signal_4845), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2575_s_current_state_reg ( .D(
        new_AGEMA_signal_4852), .CK(clk), .Q(new_AGEMA_signal_4853), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2577_s_current_state_reg ( .D(
        new_AGEMA_signal_4854), .CK(clk), .Q(new_AGEMA_signal_4855), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2579_s_current_state_reg ( .D(
        new_AGEMA_signal_4856), .CK(clk), .Q(new_AGEMA_signal_4857), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2589_s_current_state_reg ( .D(
        new_AGEMA_signal_4866), .CK(clk), .Q(new_AGEMA_signal_4867), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2593_s_current_state_reg ( .D(
        new_AGEMA_signal_4870), .CK(clk), .Q(new_AGEMA_signal_4871), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2597_s_current_state_reg ( .D(
        new_AGEMA_signal_4874), .CK(clk), .Q(new_AGEMA_signal_4875), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2599_s_current_state_reg ( .D(
        new_AGEMA_signal_4876), .CK(clk), .Q(new_AGEMA_signal_4877), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2601_s_current_state_reg ( .D(
        new_AGEMA_signal_4878), .CK(clk), .Q(new_AGEMA_signal_4879), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2603_s_current_state_reg ( .D(
        new_AGEMA_signal_4880), .CK(clk), .Q(new_AGEMA_signal_4881), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2611_s_current_state_reg ( .D(
        new_AGEMA_signal_4888), .CK(clk), .Q(new_AGEMA_signal_4889), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2613_s_current_state_reg ( .D(
        new_AGEMA_signal_4890), .CK(clk), .Q(new_AGEMA_signal_4891), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2615_s_current_state_reg ( .D(
        new_AGEMA_signal_4892), .CK(clk), .Q(new_AGEMA_signal_4893), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2625_s_current_state_reg ( .D(
        new_AGEMA_signal_4902), .CK(clk), .Q(new_AGEMA_signal_4903), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2629_s_current_state_reg ( .D(
        new_AGEMA_signal_4906), .CK(clk), .Q(new_AGEMA_signal_4907), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2633_s_current_state_reg ( .D(
        new_AGEMA_signal_4910), .CK(clk), .Q(new_AGEMA_signal_4911), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2635_s_current_state_reg ( .D(
        new_AGEMA_signal_4912), .CK(clk), .Q(new_AGEMA_signal_4913), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2637_s_current_state_reg ( .D(
        new_AGEMA_signal_4914), .CK(clk), .Q(new_AGEMA_signal_4915), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2639_s_current_state_reg ( .D(
        new_AGEMA_signal_4916), .CK(clk), .Q(new_AGEMA_signal_4917), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2643_s_current_state_reg ( .D(
        new_AGEMA_signal_4920), .CK(clk), .Q(new_AGEMA_signal_4921), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2647_s_current_state_reg ( .D(
        new_AGEMA_signal_4924), .CK(clk), .Q(new_AGEMA_signal_4925), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2651_s_current_state_reg ( .D(
        new_AGEMA_signal_4928), .CK(clk), .Q(new_AGEMA_signal_4929), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2655_s_current_state_reg ( .D(
        new_AGEMA_signal_4932), .CK(clk), .Q(new_AGEMA_signal_4933), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2659_s_current_state_reg ( .D(
        new_AGEMA_signal_4936), .CK(clk), .Q(new_AGEMA_signal_4937), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2663_s_current_state_reg ( .D(
        new_AGEMA_signal_4940), .CK(clk), .Q(new_AGEMA_signal_4941), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2667_s_current_state_reg ( .D(
        new_AGEMA_signal_4944), .CK(clk), .Q(new_AGEMA_signal_4945), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2671_s_current_state_reg ( .D(
        new_AGEMA_signal_4948), .CK(clk), .Q(new_AGEMA_signal_4949), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2675_s_current_state_reg ( .D(
        new_AGEMA_signal_4952), .CK(clk), .Q(new_AGEMA_signal_4953), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2679_s_current_state_reg ( .D(
        new_AGEMA_signal_4956), .CK(clk), .Q(new_AGEMA_signal_4957), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2683_s_current_state_reg ( .D(
        new_AGEMA_signal_4960), .CK(clk), .Q(new_AGEMA_signal_4961), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2687_s_current_state_reg ( .D(
        new_AGEMA_signal_4964), .CK(clk), .Q(new_AGEMA_signal_4965), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2691_s_current_state_reg ( .D(
        new_AGEMA_signal_4968), .CK(clk), .Q(new_AGEMA_signal_4969), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2695_s_current_state_reg ( .D(
        new_AGEMA_signal_4972), .CK(clk), .Q(new_AGEMA_signal_4973), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2699_s_current_state_reg ( .D(
        new_AGEMA_signal_4976), .CK(clk), .Q(new_AGEMA_signal_4977), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2703_s_current_state_reg ( .D(
        new_AGEMA_signal_4980), .CK(clk), .Q(new_AGEMA_signal_4981), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2707_s_current_state_reg ( .D(
        new_AGEMA_signal_4984), .CK(clk), .Q(new_AGEMA_signal_4985), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2711_s_current_state_reg ( .D(
        new_AGEMA_signal_4988), .CK(clk), .Q(new_AGEMA_signal_4989), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2715_s_current_state_reg ( .D(
        new_AGEMA_signal_4992), .CK(clk), .Q(new_AGEMA_signal_4993), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2719_s_current_state_reg ( .D(
        new_AGEMA_signal_4996), .CK(clk), .Q(new_AGEMA_signal_4997), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2723_s_current_state_reg ( .D(
        new_AGEMA_signal_5000), .CK(clk), .Q(new_AGEMA_signal_5001), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2727_s_current_state_reg ( .D(
        new_AGEMA_signal_5004), .CK(clk), .Q(new_AGEMA_signal_5005), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2731_s_current_state_reg ( .D(
        new_AGEMA_signal_5008), .CK(clk), .Q(new_AGEMA_signal_5009), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2735_s_current_state_reg ( .D(
        new_AGEMA_signal_5012), .CK(clk), .Q(new_AGEMA_signal_5013), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2739_s_current_state_reg ( .D(
        new_AGEMA_signal_5016), .CK(clk), .Q(new_AGEMA_signal_5017), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2743_s_current_state_reg ( .D(
        new_AGEMA_signal_5020), .CK(clk), .Q(new_AGEMA_signal_5021), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2747_s_current_state_reg ( .D(
        new_AGEMA_signal_5024), .CK(clk), .Q(new_AGEMA_signal_5025), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2751_s_current_state_reg ( .D(
        new_AGEMA_signal_5028), .CK(clk), .Q(new_AGEMA_signal_5029), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2755_s_current_state_reg ( .D(
        new_AGEMA_signal_5032), .CK(clk), .Q(new_AGEMA_signal_5033), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2759_s_current_state_reg ( .D(
        new_AGEMA_signal_5036), .CK(clk), .Q(new_AGEMA_signal_5037), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2763_s_current_state_reg ( .D(
        new_AGEMA_signal_5040), .CK(clk), .Q(new_AGEMA_signal_5041), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2767_s_current_state_reg ( .D(
        new_AGEMA_signal_5044), .CK(clk), .Q(new_AGEMA_signal_5045), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2771_s_current_state_reg ( .D(
        new_AGEMA_signal_5048), .CK(clk), .Q(new_AGEMA_signal_5049), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2775_s_current_state_reg ( .D(
        new_AGEMA_signal_5052), .CK(clk), .Q(new_AGEMA_signal_5053), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2779_s_current_state_reg ( .D(
        new_AGEMA_signal_5056), .CK(clk), .Q(new_AGEMA_signal_5057), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2783_s_current_state_reg ( .D(
        new_AGEMA_signal_5060), .CK(clk), .Q(new_AGEMA_signal_5061), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2787_s_current_state_reg ( .D(
        new_AGEMA_signal_5064), .CK(clk), .Q(new_AGEMA_signal_5065), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2791_s_current_state_reg ( .D(
        new_AGEMA_signal_5068), .CK(clk), .Q(new_AGEMA_signal_5069), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2795_s_current_state_reg ( .D(
        new_AGEMA_signal_5072), .CK(clk), .Q(new_AGEMA_signal_5073), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2799_s_current_state_reg ( .D(
        new_AGEMA_signal_5076), .CK(clk), .Q(new_AGEMA_signal_5077), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2803_s_current_state_reg ( .D(
        new_AGEMA_signal_5080), .CK(clk), .Q(new_AGEMA_signal_5081), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2807_s_current_state_reg ( .D(
        new_AGEMA_signal_5084), .CK(clk), .Q(new_AGEMA_signal_5085), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2811_s_current_state_reg ( .D(
        new_AGEMA_signal_5088), .CK(clk), .Q(new_AGEMA_signal_5089), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2815_s_current_state_reg ( .D(
        new_AGEMA_signal_5092), .CK(clk), .Q(new_AGEMA_signal_5093), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2819_s_current_state_reg ( .D(
        new_AGEMA_signal_5096), .CK(clk), .Q(new_AGEMA_signal_5097), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2823_s_current_state_reg ( .D(
        new_AGEMA_signal_5100), .CK(clk), .Q(new_AGEMA_signal_5101), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2827_s_current_state_reg ( .D(
        new_AGEMA_signal_5104), .CK(clk), .Q(new_AGEMA_signal_5105), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2831_s_current_state_reg ( .D(
        new_AGEMA_signal_5108), .CK(clk), .Q(new_AGEMA_signal_5109), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2835_s_current_state_reg ( .D(
        new_AGEMA_signal_5112), .CK(clk), .Q(new_AGEMA_signal_5113), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2839_s_current_state_reg ( .D(
        new_AGEMA_signal_5116), .CK(clk), .Q(new_AGEMA_signal_5117), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2843_s_current_state_reg ( .D(
        new_AGEMA_signal_5120), .CK(clk), .Q(new_AGEMA_signal_5121), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2847_s_current_state_reg ( .D(
        new_AGEMA_signal_5124), .CK(clk), .Q(new_AGEMA_signal_5125), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2849_s_current_state_reg ( .D(
        new_AGEMA_signal_5126), .CK(clk), .Q(new_AGEMA_signal_5127), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2851_s_current_state_reg ( .D(
        new_AGEMA_signal_5128), .CK(clk), .Q(new_AGEMA_signal_5129), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2853_s_current_state_reg ( .D(
        new_AGEMA_signal_5130), .CK(clk), .Q(new_AGEMA_signal_5131), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2855_s_current_state_reg ( .D(
        new_AGEMA_signal_5132), .CK(clk), .Q(new_AGEMA_signal_5133), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2857_s_current_state_reg ( .D(
        new_AGEMA_signal_5134), .CK(clk), .Q(new_AGEMA_signal_5135), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2859_s_current_state_reg ( .D(
        new_AGEMA_signal_5136), .CK(clk), .Q(new_AGEMA_signal_5137), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2861_s_current_state_reg ( .D(
        new_AGEMA_signal_5138), .CK(clk), .Q(new_AGEMA_signal_5139), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2863_s_current_state_reg ( .D(
        new_AGEMA_signal_5140), .CK(clk), .Q(new_AGEMA_signal_5141), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2865_s_current_state_reg ( .D(
        new_AGEMA_signal_5142), .CK(clk), .Q(new_AGEMA_signal_5143), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2867_s_current_state_reg ( .D(
        new_AGEMA_signal_5144), .CK(clk), .Q(new_AGEMA_signal_5145), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2869_s_current_state_reg ( .D(
        new_AGEMA_signal_5146), .CK(clk), .Q(new_AGEMA_signal_5147), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2871_s_current_state_reg ( .D(
        new_AGEMA_signal_5148), .CK(clk), .Q(new_AGEMA_signal_5149), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2873_s_current_state_reg ( .D(
        new_AGEMA_signal_5150), .CK(clk), .Q(new_AGEMA_signal_5151), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2875_s_current_state_reg ( .D(
        new_AGEMA_signal_5152), .CK(clk), .Q(new_AGEMA_signal_5153), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2877_s_current_state_reg ( .D(
        new_AGEMA_signal_5154), .CK(clk), .Q(new_AGEMA_signal_5155), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2879_s_current_state_reg ( .D(
        new_AGEMA_signal_5156), .CK(clk), .Q(new_AGEMA_signal_5157), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2881_s_current_state_reg ( .D(
        new_AGEMA_signal_5158), .CK(clk), .Q(new_AGEMA_signal_5159), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2883_s_current_state_reg ( .D(
        new_AGEMA_signal_5160), .CK(clk), .Q(new_AGEMA_signal_5161), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2885_s_current_state_reg ( .D(
        new_AGEMA_signal_5162), .CK(clk), .Q(new_AGEMA_signal_5163), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2887_s_current_state_reg ( .D(
        new_AGEMA_signal_5164), .CK(clk), .Q(new_AGEMA_signal_5165), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2889_s_current_state_reg ( .D(
        new_AGEMA_signal_5166), .CK(clk), .Q(new_AGEMA_signal_5167), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2891_s_current_state_reg ( .D(
        new_AGEMA_signal_5168), .CK(clk), .Q(new_AGEMA_signal_5169), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2893_s_current_state_reg ( .D(
        new_AGEMA_signal_5170), .CK(clk), .Q(new_AGEMA_signal_5171), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2895_s_current_state_reg ( .D(
        new_AGEMA_signal_5172), .CK(clk), .Q(new_AGEMA_signal_5173), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2897_s_current_state_reg ( .D(
        new_AGEMA_signal_5174), .CK(clk), .Q(new_AGEMA_signal_5175), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2899_s_current_state_reg ( .D(
        new_AGEMA_signal_5176), .CK(clk), .Q(new_AGEMA_signal_5177), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2901_s_current_state_reg ( .D(
        new_AGEMA_signal_5178), .CK(clk), .Q(new_AGEMA_signal_5179), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2903_s_current_state_reg ( .D(
        new_AGEMA_signal_5180), .CK(clk), .Q(new_AGEMA_signal_5181), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2905_s_current_state_reg ( .D(
        new_AGEMA_signal_5182), .CK(clk), .Q(new_AGEMA_signal_5183), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2907_s_current_state_reg ( .D(
        new_AGEMA_signal_5184), .CK(clk), .Q(new_AGEMA_signal_5185), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2909_s_current_state_reg ( .D(
        new_AGEMA_signal_5186), .CK(clk), .Q(new_AGEMA_signal_5187), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2911_s_current_state_reg ( .D(
        new_AGEMA_signal_5188), .CK(clk), .Q(new_AGEMA_signal_5189), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2913_s_current_state_reg ( .D(
        new_AGEMA_signal_5190), .CK(clk), .Q(new_AGEMA_signal_5191), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2915_s_current_state_reg ( .D(
        new_AGEMA_signal_5192), .CK(clk), .Q(new_AGEMA_signal_5193), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2917_s_current_state_reg ( .D(
        new_AGEMA_signal_5194), .CK(clk), .Q(new_AGEMA_signal_5195), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2919_s_current_state_reg ( .D(
        new_AGEMA_signal_5196), .CK(clk), .Q(new_AGEMA_signal_5197), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2921_s_current_state_reg ( .D(
        new_AGEMA_signal_5198), .CK(clk), .Q(new_AGEMA_signal_5199), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2923_s_current_state_reg ( .D(
        new_AGEMA_signal_5200), .CK(clk), .Q(new_AGEMA_signal_5201), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2925_s_current_state_reg ( .D(
        new_AGEMA_signal_5202), .CK(clk), .Q(new_AGEMA_signal_5203), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2927_s_current_state_reg ( .D(
        new_AGEMA_signal_5204), .CK(clk), .Q(new_AGEMA_signal_5205), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2929_s_current_state_reg ( .D(
        new_AGEMA_signal_5206), .CK(clk), .Q(new_AGEMA_signal_5207), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2931_s_current_state_reg ( .D(
        new_AGEMA_signal_5208), .CK(clk), .Q(new_AGEMA_signal_5209), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2933_s_current_state_reg ( .D(
        new_AGEMA_signal_5210), .CK(clk), .Q(new_AGEMA_signal_5211), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2935_s_current_state_reg ( .D(
        new_AGEMA_signal_5212), .CK(clk), .Q(new_AGEMA_signal_5213), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2937_s_current_state_reg ( .D(
        new_AGEMA_signal_5214), .CK(clk), .Q(new_AGEMA_signal_5215), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2939_s_current_state_reg ( .D(
        new_AGEMA_signal_5216), .CK(clk), .Q(new_AGEMA_signal_5217), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2941_s_current_state_reg ( .D(
        new_AGEMA_signal_5218), .CK(clk), .Q(new_AGEMA_signal_5219), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2943_s_current_state_reg ( .D(
        new_AGEMA_signal_5220), .CK(clk), .Q(new_AGEMA_signal_5221), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2945_s_current_state_reg ( .D(
        new_AGEMA_signal_5222), .CK(clk), .Q(new_AGEMA_signal_5223), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2947_s_current_state_reg ( .D(
        new_AGEMA_signal_5224), .CK(clk), .Q(new_AGEMA_signal_5225), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2949_s_current_state_reg ( .D(
        new_AGEMA_signal_5226), .CK(clk), .Q(new_AGEMA_signal_5227), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2951_s_current_state_reg ( .D(
        new_AGEMA_signal_5228), .CK(clk), .Q(new_AGEMA_signal_5229), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2953_s_current_state_reg ( .D(
        new_AGEMA_signal_5230), .CK(clk), .Q(new_AGEMA_signal_5231), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2955_s_current_state_reg ( .D(
        new_AGEMA_signal_5232), .CK(clk), .Q(new_AGEMA_signal_5233), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2957_s_current_state_reg ( .D(
        new_AGEMA_signal_5234), .CK(clk), .Q(new_AGEMA_signal_5235), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2959_s_current_state_reg ( .D(
        new_AGEMA_signal_5236), .CK(clk), .Q(new_AGEMA_signal_5237), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2961_s_current_state_reg ( .D(
        new_AGEMA_signal_5238), .CK(clk), .Q(new_AGEMA_signal_5239), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2963_s_current_state_reg ( .D(
        new_AGEMA_signal_5240), .CK(clk), .Q(new_AGEMA_signal_5241), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2965_s_current_state_reg ( .D(
        new_AGEMA_signal_5242), .CK(clk), .Q(new_AGEMA_signal_5243), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2967_s_current_state_reg ( .D(
        new_AGEMA_signal_5244), .CK(clk), .Q(new_AGEMA_signal_5245), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2969_s_current_state_reg ( .D(
        new_AGEMA_signal_5246), .CK(clk), .Q(new_AGEMA_signal_5247), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2971_s_current_state_reg ( .D(
        new_AGEMA_signal_5248), .CK(clk), .Q(new_AGEMA_signal_5249), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2973_s_current_state_reg ( .D(
        new_AGEMA_signal_5250), .CK(clk), .Q(new_AGEMA_signal_5251), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2975_s_current_state_reg ( .D(
        new_AGEMA_signal_5252), .CK(clk), .Q(new_AGEMA_signal_5253), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2977_s_current_state_reg ( .D(
        new_AGEMA_signal_5254), .CK(clk), .Q(new_AGEMA_signal_5255), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2979_s_current_state_reg ( .D(
        new_AGEMA_signal_5256), .CK(clk), .Q(new_AGEMA_signal_5257), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2981_s_current_state_reg ( .D(
        new_AGEMA_signal_5258), .CK(clk), .Q(new_AGEMA_signal_5259), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2983_s_current_state_reg ( .D(
        new_AGEMA_signal_5260), .CK(clk), .Q(new_AGEMA_signal_5261), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2985_s_current_state_reg ( .D(
        new_AGEMA_signal_5262), .CK(clk), .Q(new_AGEMA_signal_5263), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2987_s_current_state_reg ( .D(
        new_AGEMA_signal_5264), .CK(clk), .Q(new_AGEMA_signal_5265), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2989_s_current_state_reg ( .D(
        new_AGEMA_signal_5266), .CK(clk), .Q(new_AGEMA_signal_5267), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2991_s_current_state_reg ( .D(
        new_AGEMA_signal_5268), .CK(clk), .Q(new_AGEMA_signal_5269), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2993_s_current_state_reg ( .D(
        new_AGEMA_signal_5270), .CK(clk), .Q(new_AGEMA_signal_5271), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2995_s_current_state_reg ( .D(
        new_AGEMA_signal_5272), .CK(clk), .Q(new_AGEMA_signal_5273), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2997_s_current_state_reg ( .D(
        new_AGEMA_signal_5274), .CK(clk), .Q(new_AGEMA_signal_5275), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_2999_s_current_state_reg ( .D(
        new_AGEMA_signal_5276), .CK(clk), .Q(new_AGEMA_signal_5277), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3001_s_current_state_reg ( .D(
        new_AGEMA_signal_5278), .CK(clk), .Q(new_AGEMA_signal_5279), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3003_s_current_state_reg ( .D(
        new_AGEMA_signal_5280), .CK(clk), .Q(new_AGEMA_signal_5281), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3005_s_current_state_reg ( .D(
        new_AGEMA_signal_5282), .CK(clk), .Q(new_AGEMA_signal_5283), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3007_s_current_state_reg ( .D(
        new_AGEMA_signal_5284), .CK(clk), .Q(new_AGEMA_signal_5285), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3009_s_current_state_reg ( .D(
        new_AGEMA_signal_5286), .CK(clk), .Q(new_AGEMA_signal_5287), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3011_s_current_state_reg ( .D(
        new_AGEMA_signal_5288), .CK(clk), .Q(new_AGEMA_signal_5289), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3013_s_current_state_reg ( .D(
        new_AGEMA_signal_5290), .CK(clk), .Q(new_AGEMA_signal_5291), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3015_s_current_state_reg ( .D(
        new_AGEMA_signal_5292), .CK(clk), .Q(new_AGEMA_signal_5293), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3017_s_current_state_reg ( .D(
        new_AGEMA_signal_5294), .CK(clk), .Q(new_AGEMA_signal_5295), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3019_s_current_state_reg ( .D(
        new_AGEMA_signal_5296), .CK(clk), .Q(new_AGEMA_signal_5297), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3021_s_current_state_reg ( .D(
        new_AGEMA_signal_5298), .CK(clk), .Q(new_AGEMA_signal_5299), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3023_s_current_state_reg ( .D(
        new_AGEMA_signal_5300), .CK(clk), .Q(new_AGEMA_signal_5301), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3025_s_current_state_reg ( .D(
        new_AGEMA_signal_5302), .CK(clk), .Q(new_AGEMA_signal_5303), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3027_s_current_state_reg ( .D(
        new_AGEMA_signal_5304), .CK(clk), .Q(new_AGEMA_signal_5305), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3029_s_current_state_reg ( .D(
        new_AGEMA_signal_5306), .CK(clk), .Q(new_AGEMA_signal_5307), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3031_s_current_state_reg ( .D(
        new_AGEMA_signal_5308), .CK(clk), .Q(new_AGEMA_signal_5309), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3033_s_current_state_reg ( .D(
        new_AGEMA_signal_5310), .CK(clk), .Q(new_AGEMA_signal_5311), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3035_s_current_state_reg ( .D(
        new_AGEMA_signal_5312), .CK(clk), .Q(new_AGEMA_signal_5313), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3037_s_current_state_reg ( .D(
        new_AGEMA_signal_5314), .CK(clk), .Q(new_AGEMA_signal_5315), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3039_s_current_state_reg ( .D(
        new_AGEMA_signal_5316), .CK(clk), .Q(new_AGEMA_signal_5317), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3043_s_current_state_reg ( .D(
        new_AGEMA_signal_5320), .CK(clk), .Q(new_AGEMA_signal_5321), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3047_s_current_state_reg ( .D(
        new_AGEMA_signal_5324), .CK(clk), .Q(new_AGEMA_signal_5325), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3051_s_current_state_reg ( .D(
        new_AGEMA_signal_5328), .CK(clk), .Q(new_AGEMA_signal_5329), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3055_s_current_state_reg ( .D(
        new_AGEMA_signal_5332), .CK(clk), .Q(new_AGEMA_signal_5333), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3059_s_current_state_reg ( .D(
        new_AGEMA_signal_5336), .CK(clk), .Q(new_AGEMA_signal_5337), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3063_s_current_state_reg ( .D(
        new_AGEMA_signal_5340), .CK(clk), .Q(new_AGEMA_signal_5341), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3067_s_current_state_reg ( .D(
        new_AGEMA_signal_5344), .CK(clk), .Q(new_AGEMA_signal_5345), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3071_s_current_state_reg ( .D(
        new_AGEMA_signal_5348), .CK(clk), .Q(new_AGEMA_signal_5349), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3075_s_current_state_reg ( .D(
        new_AGEMA_signal_5352), .CK(clk), .Q(new_AGEMA_signal_5353), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3079_s_current_state_reg ( .D(
        new_AGEMA_signal_5356), .CK(clk), .Q(new_AGEMA_signal_5357), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3083_s_current_state_reg ( .D(
        new_AGEMA_signal_5360), .CK(clk), .Q(new_AGEMA_signal_5361), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3087_s_current_state_reg ( .D(
        new_AGEMA_signal_5364), .CK(clk), .Q(new_AGEMA_signal_5365), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3091_s_current_state_reg ( .D(
        new_AGEMA_signal_5368), .CK(clk), .Q(new_AGEMA_signal_5369), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3095_s_current_state_reg ( .D(
        new_AGEMA_signal_5372), .CK(clk), .Q(new_AGEMA_signal_5373), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3099_s_current_state_reg ( .D(
        new_AGEMA_signal_5376), .CK(clk), .Q(new_AGEMA_signal_5377), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3103_s_current_state_reg ( .D(
        new_AGEMA_signal_5380), .CK(clk), .Q(new_AGEMA_signal_5381), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3107_s_current_state_reg ( .D(
        new_AGEMA_signal_5384), .CK(clk), .Q(new_AGEMA_signal_5385), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3111_s_current_state_reg ( .D(
        new_AGEMA_signal_5388), .CK(clk), .Q(new_AGEMA_signal_5389), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3115_s_current_state_reg ( .D(
        new_AGEMA_signal_5392), .CK(clk), .Q(new_AGEMA_signal_5393), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3119_s_current_state_reg ( .D(
        new_AGEMA_signal_5396), .CK(clk), .Q(new_AGEMA_signal_5397), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3123_s_current_state_reg ( .D(
        new_AGEMA_signal_5400), .CK(clk), .Q(new_AGEMA_signal_5401), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3127_s_current_state_reg ( .D(
        new_AGEMA_signal_5404), .CK(clk), .Q(new_AGEMA_signal_5405), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3131_s_current_state_reg ( .D(
        new_AGEMA_signal_5408), .CK(clk), .Q(new_AGEMA_signal_5409), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3135_s_current_state_reg ( .D(
        new_AGEMA_signal_5412), .CK(clk), .Q(new_AGEMA_signal_5413), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3139_s_current_state_reg ( .D(
        new_AGEMA_signal_5416), .CK(clk), .Q(new_AGEMA_signal_5417), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3143_s_current_state_reg ( .D(
        new_AGEMA_signal_5420), .CK(clk), .Q(new_AGEMA_signal_5421), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3147_s_current_state_reg ( .D(
        new_AGEMA_signal_5424), .CK(clk), .Q(new_AGEMA_signal_5425), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3151_s_current_state_reg ( .D(
        new_AGEMA_signal_5428), .CK(clk), .Q(new_AGEMA_signal_5429), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3155_s_current_state_reg ( .D(
        new_AGEMA_signal_5432), .CK(clk), .Q(new_AGEMA_signal_5433), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3159_s_current_state_reg ( .D(
        new_AGEMA_signal_5436), .CK(clk), .Q(new_AGEMA_signal_5437), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3163_s_current_state_reg ( .D(
        new_AGEMA_signal_5440), .CK(clk), .Q(new_AGEMA_signal_5441), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3167_s_current_state_reg ( .D(
        new_AGEMA_signal_5444), .CK(clk), .Q(new_AGEMA_signal_5445), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3171_s_current_state_reg ( .D(
        new_AGEMA_signal_5448), .CK(clk), .Q(new_AGEMA_signal_5449), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3175_s_current_state_reg ( .D(
        new_AGEMA_signal_5452), .CK(clk), .Q(new_AGEMA_signal_5453), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3179_s_current_state_reg ( .D(
        new_AGEMA_signal_5456), .CK(clk), .Q(new_AGEMA_signal_5457), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3183_s_current_state_reg ( .D(
        new_AGEMA_signal_5460), .CK(clk), .Q(new_AGEMA_signal_5461), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3187_s_current_state_reg ( .D(
        new_AGEMA_signal_5464), .CK(clk), .Q(new_AGEMA_signal_5465), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3191_s_current_state_reg ( .D(
        new_AGEMA_signal_5468), .CK(clk), .Q(new_AGEMA_signal_5469), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3195_s_current_state_reg ( .D(
        new_AGEMA_signal_5472), .CK(clk), .Q(new_AGEMA_signal_5473), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3199_s_current_state_reg ( .D(
        new_AGEMA_signal_5476), .CK(clk), .Q(new_AGEMA_signal_5477), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3203_s_current_state_reg ( .D(
        new_AGEMA_signal_5480), .CK(clk), .Q(new_AGEMA_signal_5481), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3207_s_current_state_reg ( .D(
        new_AGEMA_signal_5484), .CK(clk), .Q(new_AGEMA_signal_5485), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3211_s_current_state_reg ( .D(
        new_AGEMA_signal_5488), .CK(clk), .Q(new_AGEMA_signal_5489), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3215_s_current_state_reg ( .D(
        new_AGEMA_signal_5492), .CK(clk), .Q(new_AGEMA_signal_5493), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3219_s_current_state_reg ( .D(
        new_AGEMA_signal_5496), .CK(clk), .Q(new_AGEMA_signal_5497), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3223_s_current_state_reg ( .D(
        new_AGEMA_signal_5500), .CK(clk), .Q(new_AGEMA_signal_5501), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3227_s_current_state_reg ( .D(
        new_AGEMA_signal_5504), .CK(clk), .Q(new_AGEMA_signal_5505), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3231_s_current_state_reg ( .D(
        new_AGEMA_signal_5508), .CK(clk), .Q(new_AGEMA_signal_5509), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3235_s_current_state_reg ( .D(
        new_AGEMA_signal_5512), .CK(clk), .Q(new_AGEMA_signal_5513), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3239_s_current_state_reg ( .D(
        new_AGEMA_signal_5516), .CK(clk), .Q(new_AGEMA_signal_5517), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3243_s_current_state_reg ( .D(
        new_AGEMA_signal_5520), .CK(clk), .Q(new_AGEMA_signal_5521), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3247_s_current_state_reg ( .D(
        new_AGEMA_signal_5524), .CK(clk), .Q(new_AGEMA_signal_5525), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3251_s_current_state_reg ( .D(
        new_AGEMA_signal_5528), .CK(clk), .Q(new_AGEMA_signal_5529), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3255_s_current_state_reg ( .D(
        new_AGEMA_signal_5532), .CK(clk), .Q(new_AGEMA_signal_5533), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3259_s_current_state_reg ( .D(
        new_AGEMA_signal_5536), .CK(clk), .Q(new_AGEMA_signal_5537), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3263_s_current_state_reg ( .D(
        new_AGEMA_signal_5540), .CK(clk), .Q(new_AGEMA_signal_5541), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3267_s_current_state_reg ( .D(
        new_AGEMA_signal_5544), .CK(clk), .Q(new_AGEMA_signal_5545), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3271_s_current_state_reg ( .D(
        new_AGEMA_signal_5548), .CK(clk), .Q(new_AGEMA_signal_5549), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3275_s_current_state_reg ( .D(
        new_AGEMA_signal_5552), .CK(clk), .Q(new_AGEMA_signal_5553), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3279_s_current_state_reg ( .D(
        new_AGEMA_signal_5556), .CK(clk), .Q(new_AGEMA_signal_5557), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3283_s_current_state_reg ( .D(
        new_AGEMA_signal_5560), .CK(clk), .Q(new_AGEMA_signal_5561), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3287_s_current_state_reg ( .D(
        new_AGEMA_signal_5564), .CK(clk), .Q(new_AGEMA_signal_5565), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3291_s_current_state_reg ( .D(
        new_AGEMA_signal_5568), .CK(clk), .Q(new_AGEMA_signal_5569), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3295_s_current_state_reg ( .D(
        new_AGEMA_signal_5572), .CK(clk), .Q(new_AGEMA_signal_5573), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3299_s_current_state_reg ( .D(
        new_AGEMA_signal_5576), .CK(clk), .Q(new_AGEMA_signal_5577), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3303_s_current_state_reg ( .D(
        new_AGEMA_signal_5580), .CK(clk), .Q(new_AGEMA_signal_5581), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3307_s_current_state_reg ( .D(
        new_AGEMA_signal_5584), .CK(clk), .Q(new_AGEMA_signal_5585), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3311_s_current_state_reg ( .D(
        new_AGEMA_signal_5588), .CK(clk), .Q(new_AGEMA_signal_5589), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3315_s_current_state_reg ( .D(
        new_AGEMA_signal_5592), .CK(clk), .Q(new_AGEMA_signal_5593), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3319_s_current_state_reg ( .D(
        new_AGEMA_signal_5596), .CK(clk), .Q(new_AGEMA_signal_5597), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3323_s_current_state_reg ( .D(
        new_AGEMA_signal_5600), .CK(clk), .Q(new_AGEMA_signal_5601), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3327_s_current_state_reg ( .D(
        new_AGEMA_signal_5604), .CK(clk), .Q(new_AGEMA_signal_5605), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3331_s_current_state_reg ( .D(
        new_AGEMA_signal_5608), .CK(clk), .Q(new_AGEMA_signal_5609), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3335_s_current_state_reg ( .D(
        new_AGEMA_signal_5612), .CK(clk), .Q(new_AGEMA_signal_5613), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3339_s_current_state_reg ( .D(
        new_AGEMA_signal_5616), .CK(clk), .Q(new_AGEMA_signal_5617), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3343_s_current_state_reg ( .D(
        new_AGEMA_signal_5620), .CK(clk), .Q(new_AGEMA_signal_5621), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3347_s_current_state_reg ( .D(
        new_AGEMA_signal_5624), .CK(clk), .Q(new_AGEMA_signal_5625), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3351_s_current_state_reg ( .D(
        new_AGEMA_signal_5628), .CK(clk), .Q(new_AGEMA_signal_5629), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3355_s_current_state_reg ( .D(
        new_AGEMA_signal_5632), .CK(clk), .Q(new_AGEMA_signal_5633), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3359_s_current_state_reg ( .D(
        new_AGEMA_signal_5636), .CK(clk), .Q(new_AGEMA_signal_5637), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3363_s_current_state_reg ( .D(
        new_AGEMA_signal_5640), .CK(clk), .Q(new_AGEMA_signal_5641), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3367_s_current_state_reg ( .D(
        new_AGEMA_signal_5644), .CK(clk), .Q(new_AGEMA_signal_5645), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3371_s_current_state_reg ( .D(
        new_AGEMA_signal_5648), .CK(clk), .Q(new_AGEMA_signal_5649), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3375_s_current_state_reg ( .D(
        new_AGEMA_signal_5652), .CK(clk), .Q(new_AGEMA_signal_5653), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3379_s_current_state_reg ( .D(
        new_AGEMA_signal_5656), .CK(clk), .Q(new_AGEMA_signal_5657), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3383_s_current_state_reg ( .D(
        new_AGEMA_signal_5660), .CK(clk), .Q(new_AGEMA_signal_5661), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3387_s_current_state_reg ( .D(
        new_AGEMA_signal_5664), .CK(clk), .Q(new_AGEMA_signal_5665), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3391_s_current_state_reg ( .D(
        new_AGEMA_signal_5668), .CK(clk), .Q(new_AGEMA_signal_5669), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3395_s_current_state_reg ( .D(
        new_AGEMA_signal_5672), .CK(clk), .Q(new_AGEMA_signal_5673), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3399_s_current_state_reg ( .D(
        new_AGEMA_signal_5676), .CK(clk), .Q(new_AGEMA_signal_5677), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3403_s_current_state_reg ( .D(
        new_AGEMA_signal_5680), .CK(clk), .Q(new_AGEMA_signal_5681), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3407_s_current_state_reg ( .D(
        new_AGEMA_signal_5684), .CK(clk), .Q(new_AGEMA_signal_5685), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3411_s_current_state_reg ( .D(
        new_AGEMA_signal_5688), .CK(clk), .Q(new_AGEMA_signal_5689), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3415_s_current_state_reg ( .D(
        new_AGEMA_signal_5692), .CK(clk), .Q(new_AGEMA_signal_5693), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3419_s_current_state_reg ( .D(
        new_AGEMA_signal_5696), .CK(clk), .Q(new_AGEMA_signal_5697), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3423_s_current_state_reg ( .D(
        new_AGEMA_signal_5700), .CK(clk), .Q(new_AGEMA_signal_5701), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3427_s_current_state_reg ( .D(
        new_AGEMA_signal_5704), .CK(clk), .Q(new_AGEMA_signal_5705), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3431_s_current_state_reg ( .D(
        new_AGEMA_signal_5708), .CK(clk), .Q(new_AGEMA_signal_5709), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3435_s_current_state_reg ( .D(
        new_AGEMA_signal_5712), .CK(clk), .Q(new_AGEMA_signal_5713), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3439_s_current_state_reg ( .D(
        new_AGEMA_signal_5716), .CK(clk), .Q(new_AGEMA_signal_5717), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3443_s_current_state_reg ( .D(
        new_AGEMA_signal_5720), .CK(clk), .Q(new_AGEMA_signal_5721), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3447_s_current_state_reg ( .D(
        new_AGEMA_signal_5724), .CK(clk), .Q(new_AGEMA_signal_5725), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3451_s_current_state_reg ( .D(
        new_AGEMA_signal_5728), .CK(clk), .Q(new_AGEMA_signal_5729), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3455_s_current_state_reg ( .D(
        new_AGEMA_signal_5732), .CK(clk), .Q(new_AGEMA_signal_5733), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3459_s_current_state_reg ( .D(
        new_AGEMA_signal_5736), .CK(clk), .Q(new_AGEMA_signal_5737), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3463_s_current_state_reg ( .D(
        new_AGEMA_signal_5740), .CK(clk), .Q(new_AGEMA_signal_5741), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3467_s_current_state_reg ( .D(
        new_AGEMA_signal_5744), .CK(clk), .Q(new_AGEMA_signal_5745), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3471_s_current_state_reg ( .D(
        new_AGEMA_signal_5748), .CK(clk), .Q(new_AGEMA_signal_5749), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3475_s_current_state_reg ( .D(
        new_AGEMA_signal_5752), .CK(clk), .Q(new_AGEMA_signal_5753), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3479_s_current_state_reg ( .D(
        new_AGEMA_signal_5756), .CK(clk), .Q(new_AGEMA_signal_5757), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3483_s_current_state_reg ( .D(
        new_AGEMA_signal_5760), .CK(clk), .Q(new_AGEMA_signal_5761), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3487_s_current_state_reg ( .D(
        new_AGEMA_signal_5764), .CK(clk), .Q(new_AGEMA_signal_5765), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3491_s_current_state_reg ( .D(
        new_AGEMA_signal_5768), .CK(clk), .Q(new_AGEMA_signal_5769), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3495_s_current_state_reg ( .D(
        new_AGEMA_signal_5772), .CK(clk), .Q(new_AGEMA_signal_5773), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3499_s_current_state_reg ( .D(
        new_AGEMA_signal_5776), .CK(clk), .Q(new_AGEMA_signal_5777), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3503_s_current_state_reg ( .D(
        new_AGEMA_signal_5780), .CK(clk), .Q(new_AGEMA_signal_5781), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3507_s_current_state_reg ( .D(
        new_AGEMA_signal_5784), .CK(clk), .Q(new_AGEMA_signal_5785), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3511_s_current_state_reg ( .D(
        new_AGEMA_signal_5788), .CK(clk), .Q(new_AGEMA_signal_5789), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3515_s_current_state_reg ( .D(
        new_AGEMA_signal_5792), .CK(clk), .Q(new_AGEMA_signal_5793), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3519_s_current_state_reg ( .D(
        new_AGEMA_signal_5796), .CK(clk), .Q(new_AGEMA_signal_5797), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3523_s_current_state_reg ( .D(
        new_AGEMA_signal_5800), .CK(clk), .Q(new_AGEMA_signal_5801), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3527_s_current_state_reg ( .D(
        new_AGEMA_signal_5804), .CK(clk), .Q(new_AGEMA_signal_5805), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3531_s_current_state_reg ( .D(
        new_AGEMA_signal_5808), .CK(clk), .Q(new_AGEMA_signal_5809), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3535_s_current_state_reg ( .D(
        new_AGEMA_signal_5812), .CK(clk), .Q(new_AGEMA_signal_5813), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3539_s_current_state_reg ( .D(
        new_AGEMA_signal_5816), .CK(clk), .Q(new_AGEMA_signal_5817), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3543_s_current_state_reg ( .D(
        new_AGEMA_signal_5820), .CK(clk), .Q(new_AGEMA_signal_5821), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3547_s_current_state_reg ( .D(
        new_AGEMA_signal_5824), .CK(clk), .Q(new_AGEMA_signal_5825), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3551_s_current_state_reg ( .D(
        new_AGEMA_signal_5828), .CK(clk), .Q(new_AGEMA_signal_5829), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3555_s_current_state_reg ( .D(
        new_AGEMA_signal_5832), .CK(clk), .Q(new_AGEMA_signal_5833), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3559_s_current_state_reg ( .D(
        new_AGEMA_signal_5836), .CK(clk), .Q(new_AGEMA_signal_5837), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3563_s_current_state_reg ( .D(
        new_AGEMA_signal_5840), .CK(clk), .Q(new_AGEMA_signal_5841), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3567_s_current_state_reg ( .D(
        new_AGEMA_signal_5844), .CK(clk), .Q(new_AGEMA_signal_5845), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3571_s_current_state_reg ( .D(
        new_AGEMA_signal_5848), .CK(clk), .Q(new_AGEMA_signal_5849), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3575_s_current_state_reg ( .D(
        new_AGEMA_signal_5852), .CK(clk), .Q(new_AGEMA_signal_5853), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3579_s_current_state_reg ( .D(
        new_AGEMA_signal_5856), .CK(clk), .Q(new_AGEMA_signal_5857), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3583_s_current_state_reg ( .D(
        new_AGEMA_signal_5860), .CK(clk), .Q(new_AGEMA_signal_5861), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3587_s_current_state_reg ( .D(
        new_AGEMA_signal_5864), .CK(clk), .Q(new_AGEMA_signal_5865), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3591_s_current_state_reg ( .D(
        new_AGEMA_signal_5868), .CK(clk), .Q(new_AGEMA_signal_5869), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3595_s_current_state_reg ( .D(
        new_AGEMA_signal_5872), .CK(clk), .Q(new_AGEMA_signal_5873), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3599_s_current_state_reg ( .D(
        new_AGEMA_signal_5876), .CK(clk), .Q(new_AGEMA_signal_5877), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3603_s_current_state_reg ( .D(
        new_AGEMA_signal_5880), .CK(clk), .Q(new_AGEMA_signal_5881), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3607_s_current_state_reg ( .D(
        new_AGEMA_signal_5884), .CK(clk), .Q(new_AGEMA_signal_5885), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3611_s_current_state_reg ( .D(
        new_AGEMA_signal_5888), .CK(clk), .Q(new_AGEMA_signal_5889), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3615_s_current_state_reg ( .D(
        new_AGEMA_signal_5892), .CK(clk), .Q(new_AGEMA_signal_5893), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3619_s_current_state_reg ( .D(
        new_AGEMA_signal_5896), .CK(clk), .Q(new_AGEMA_signal_5897), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3623_s_current_state_reg ( .D(
        new_AGEMA_signal_5900), .CK(clk), .Q(new_AGEMA_signal_5901), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3627_s_current_state_reg ( .D(
        new_AGEMA_signal_5904), .CK(clk), .Q(new_AGEMA_signal_5905), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3631_s_current_state_reg ( .D(
        new_AGEMA_signal_5908), .CK(clk), .Q(new_AGEMA_signal_5909), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3635_s_current_state_reg ( .D(
        new_AGEMA_signal_5912), .CK(clk), .Q(new_AGEMA_signal_5913), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3639_s_current_state_reg ( .D(
        new_AGEMA_signal_5916), .CK(clk), .Q(new_AGEMA_signal_5917), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3643_s_current_state_reg ( .D(
        new_AGEMA_signal_5920), .CK(clk), .Q(new_AGEMA_signal_5921), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3647_s_current_state_reg ( .D(
        new_AGEMA_signal_5924), .CK(clk), .Q(new_AGEMA_signal_5925), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3651_s_current_state_reg ( .D(
        new_AGEMA_signal_5928), .CK(clk), .Q(new_AGEMA_signal_5929), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3655_s_current_state_reg ( .D(
        new_AGEMA_signal_5932), .CK(clk), .Q(new_AGEMA_signal_5933), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3659_s_current_state_reg ( .D(
        new_AGEMA_signal_5936), .CK(clk), .Q(new_AGEMA_signal_5937), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3663_s_current_state_reg ( .D(
        new_AGEMA_signal_5940), .CK(clk), .Q(new_AGEMA_signal_5941), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3667_s_current_state_reg ( .D(
        new_AGEMA_signal_5944), .CK(clk), .Q(new_AGEMA_signal_5945), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3671_s_current_state_reg ( .D(
        new_AGEMA_signal_5948), .CK(clk), .Q(new_AGEMA_signal_5949), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3675_s_current_state_reg ( .D(
        new_AGEMA_signal_5952), .CK(clk), .Q(new_AGEMA_signal_5953), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3679_s_current_state_reg ( .D(
        new_AGEMA_signal_5956), .CK(clk), .Q(new_AGEMA_signal_5957), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3683_s_current_state_reg ( .D(
        new_AGEMA_signal_5960), .CK(clk), .Q(new_AGEMA_signal_5961), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3687_s_current_state_reg ( .D(
        new_AGEMA_signal_5964), .CK(clk), .Q(new_AGEMA_signal_5965), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3691_s_current_state_reg ( .D(
        new_AGEMA_signal_5968), .CK(clk), .Q(new_AGEMA_signal_5969), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3695_s_current_state_reg ( .D(
        new_AGEMA_signal_5972), .CK(clk), .Q(new_AGEMA_signal_5973), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3699_s_current_state_reg ( .D(
        new_AGEMA_signal_5976), .CK(clk), .Q(new_AGEMA_signal_5977), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3703_s_current_state_reg ( .D(
        new_AGEMA_signal_5980), .CK(clk), .Q(new_AGEMA_signal_5981), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3707_s_current_state_reg ( .D(
        new_AGEMA_signal_5984), .CK(clk), .Q(new_AGEMA_signal_5985), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3711_s_current_state_reg ( .D(
        new_AGEMA_signal_5988), .CK(clk), .Q(new_AGEMA_signal_5989), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3715_s_current_state_reg ( .D(
        new_AGEMA_signal_5992), .CK(clk), .Q(new_AGEMA_signal_5993), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3719_s_current_state_reg ( .D(
        new_AGEMA_signal_5996), .CK(clk), .Q(new_AGEMA_signal_5997), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3723_s_current_state_reg ( .D(
        new_AGEMA_signal_6000), .CK(clk), .Q(new_AGEMA_signal_6001), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3727_s_current_state_reg ( .D(
        new_AGEMA_signal_6004), .CK(clk), .Q(new_AGEMA_signal_6005), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3731_s_current_state_reg ( .D(
        new_AGEMA_signal_6008), .CK(clk), .Q(new_AGEMA_signal_6009), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3735_s_current_state_reg ( .D(
        new_AGEMA_signal_6012), .CK(clk), .Q(new_AGEMA_signal_6013), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3739_s_current_state_reg ( .D(
        new_AGEMA_signal_6016), .CK(clk), .Q(new_AGEMA_signal_6017), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3743_s_current_state_reg ( .D(
        new_AGEMA_signal_6020), .CK(clk), .Q(new_AGEMA_signal_6021), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3747_s_current_state_reg ( .D(
        new_AGEMA_signal_6024), .CK(clk), .Q(new_AGEMA_signal_6025), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3751_s_current_state_reg ( .D(
        new_AGEMA_signal_6028), .CK(clk), .Q(new_AGEMA_signal_6029), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3755_s_current_state_reg ( .D(
        new_AGEMA_signal_6032), .CK(clk), .Q(new_AGEMA_signal_6033), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3759_s_current_state_reg ( .D(
        new_AGEMA_signal_6036), .CK(clk), .Q(new_AGEMA_signal_6037), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3763_s_current_state_reg ( .D(
        new_AGEMA_signal_6040), .CK(clk), .Q(new_AGEMA_signal_6041), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3767_s_current_state_reg ( .D(
        new_AGEMA_signal_6044), .CK(clk), .Q(new_AGEMA_signal_6045), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3771_s_current_state_reg ( .D(
        new_AGEMA_signal_6048), .CK(clk), .Q(new_AGEMA_signal_6049), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3775_s_current_state_reg ( .D(
        new_AGEMA_signal_6052), .CK(clk), .Q(new_AGEMA_signal_6053), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3779_s_current_state_reg ( .D(
        new_AGEMA_signal_6056), .CK(clk), .Q(new_AGEMA_signal_6057), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3783_s_current_state_reg ( .D(
        new_AGEMA_signal_6060), .CK(clk), .Q(new_AGEMA_signal_6061), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3787_s_current_state_reg ( .D(
        new_AGEMA_signal_6064), .CK(clk), .Q(new_AGEMA_signal_6065), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3791_s_current_state_reg ( .D(
        new_AGEMA_signal_6068), .CK(clk), .Q(new_AGEMA_signal_6069), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3795_s_current_state_reg ( .D(
        new_AGEMA_signal_6072), .CK(clk), .Q(new_AGEMA_signal_6073), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3799_s_current_state_reg ( .D(
        new_AGEMA_signal_6076), .CK(clk), .Q(new_AGEMA_signal_6077), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3803_s_current_state_reg ( .D(
        new_AGEMA_signal_6080), .CK(clk), .Q(new_AGEMA_signal_6081), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3807_s_current_state_reg ( .D(
        new_AGEMA_signal_6084), .CK(clk), .Q(new_AGEMA_signal_6085), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3811_s_current_state_reg ( .D(
        new_AGEMA_signal_6088), .CK(clk), .Q(new_AGEMA_signal_6089), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3815_s_current_state_reg ( .D(
        new_AGEMA_signal_6092), .CK(clk), .Q(new_AGEMA_signal_6093), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3819_s_current_state_reg ( .D(
        new_AGEMA_signal_6096), .CK(clk), .Q(new_AGEMA_signal_6097), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3823_s_current_state_reg ( .D(
        new_AGEMA_signal_6100), .CK(clk), .Q(new_AGEMA_signal_6101), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3827_s_current_state_reg ( .D(
        new_AGEMA_signal_6104), .CK(clk), .Q(new_AGEMA_signal_6105), .QN() );
  DFF_X1 new_AGEMA_reg_buffer_3831_s_current_state_reg ( .D(
        new_AGEMA_signal_6108), .CK(clk), .Q(new_AGEMA_signal_6109), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5127), .CK(clk), .Q(Ciphertext_s0[63]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5129), .CK(clk), .Q(Ciphertext_s1[63]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5131), .CK(clk), .Q(Ciphertext_s2[63]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5133), .CK(clk), .Q(Ciphertext_s0[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5135), .CK(clk), .Q(Ciphertext_s1[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5137), .CK(clk), .Q(Ciphertext_s2[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[61]), .CK(clk), .Q(Ciphertext_s0[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3084), .CK(clk), .Q(Ciphertext_s1[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3085), .CK(clk), .Q(Ciphertext_s2[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[60]), .CK(clk), .Q(Ciphertext_s0[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3066), .CK(clk), .Q(Ciphertext_s1[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3067), .CK(clk), .Q(Ciphertext_s2[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5139), .CK(clk), .Q(Ciphertext_s0[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5141), .CK(clk), .Q(Ciphertext_s1[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5143), .CK(clk), .Q(Ciphertext_s2[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5145), .CK(clk), .Q(Ciphertext_s0[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5147), .CK(clk), .Q(Ciphertext_s1[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5149), .CK(clk), .Q(Ciphertext_s2[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[57]), .CK(clk), .Q(Ciphertext_s0[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3038), .CK(clk), .Q(Ciphertext_s1[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3039), .CK(clk), .Q(Ciphertext_s2[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[56]), .CK(clk), .Q(Ciphertext_s0[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2952), .CK(clk), .Q(Ciphertext_s1[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2953), .CK(clk), .Q(Ciphertext_s2[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5151), .CK(clk), .Q(Ciphertext_s0[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5153), .CK(clk), .Q(Ciphertext_s1[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5155), .CK(clk), .Q(Ciphertext_s2[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5157), .CK(clk), .Q(Ciphertext_s0[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5159), .CK(clk), .Q(Ciphertext_s1[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5161), .CK(clk), .Q(Ciphertext_s2[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[53]), .CK(clk), .Q(Ciphertext_s0[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3034), .CK(clk), .Q(Ciphertext_s1[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3035), .CK(clk), .Q(Ciphertext_s2[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[52]), .CK(clk), .Q(Ciphertext_s0[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2948), .CK(clk), .Q(Ciphertext_s1[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2949), .CK(clk), .Q(Ciphertext_s2[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5163), .CK(clk), .Q(Ciphertext_s0[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5165), .CK(clk), .Q(Ciphertext_s1[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5167), .CK(clk), .Q(Ciphertext_s2[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5169), .CK(clk), .Q(Ciphertext_s0[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5171), .CK(clk), .Q(Ciphertext_s1[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5173), .CK(clk), .Q(Ciphertext_s2[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[49]), .CK(clk), .Q(Ciphertext_s0[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3030), .CK(clk), .Q(Ciphertext_s1[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3031), .CK(clk), .Q(Ciphertext_s2[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[48]), .CK(clk), .Q(Ciphertext_s0[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2944), .CK(clk), .Q(Ciphertext_s1[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2945), .CK(clk), .Q(Ciphertext_s2[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5175), .CK(clk), .Q(Ciphertext_s0[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5177), .CK(clk), .Q(Ciphertext_s1[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5179), .CK(clk), .Q(Ciphertext_s2[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5181), .CK(clk), .Q(Ciphertext_s0[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5183), .CK(clk), .Q(Ciphertext_s1[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5185), .CK(clk), .Q(Ciphertext_s2[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[45]), .CK(clk), .Q(Ciphertext_s0[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3026), .CK(clk), .Q(Ciphertext_s1[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3027), .CK(clk), .Q(Ciphertext_s2[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[44]), .CK(clk), .Q(Ciphertext_s0[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2940), .CK(clk), .Q(Ciphertext_s1[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2941), .CK(clk), .Q(Ciphertext_s2[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5187), .CK(clk), .Q(Ciphertext_s0[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5189), .CK(clk), .Q(Ciphertext_s1[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5191), .CK(clk), .Q(Ciphertext_s2[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5193), .CK(clk), .Q(Ciphertext_s0[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5195), .CK(clk), .Q(Ciphertext_s1[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5197), .CK(clk), .Q(Ciphertext_s2[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[41]), .CK(clk), .Q(Ciphertext_s0[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2832), .CK(clk), .Q(Ciphertext_s1[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2833), .CK(clk), .Q(Ciphertext_s2[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[40]), .CK(clk), .Q(Ciphertext_s0[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2712), .CK(clk), .Q(Ciphertext_s1[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2713), .CK(clk), .Q(Ciphertext_s2[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5199), .CK(clk), .Q(Ciphertext_s0[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5201), .CK(clk), .Q(Ciphertext_s1[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5203), .CK(clk), .Q(Ciphertext_s2[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5205), .CK(clk), .Q(Ciphertext_s0[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5207), .CK(clk), .Q(Ciphertext_s1[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5209), .CK(clk), .Q(Ciphertext_s2[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[37]), .CK(clk), .Q(Ciphertext_s0[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2828), .CK(clk), .Q(Ciphertext_s1[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2829), .CK(clk), .Q(Ciphertext_s2[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[36]), .CK(clk), .Q(Ciphertext_s0[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2708), .CK(clk), .Q(Ciphertext_s1[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2709), .CK(clk), .Q(Ciphertext_s2[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5211), .CK(clk), .Q(Ciphertext_s0[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5213), .CK(clk), .Q(Ciphertext_s1[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5215), .CK(clk), .Q(Ciphertext_s2[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5217), .CK(clk), .Q(Ciphertext_s0[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5219), .CK(clk), .Q(Ciphertext_s1[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5221), .CK(clk), .Q(Ciphertext_s2[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[33]), .CK(clk), .Q(Ciphertext_s0[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2824), .CK(clk), .Q(Ciphertext_s1[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2825), .CK(clk), .Q(Ciphertext_s2[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[32]), .CK(clk), .Q(Ciphertext_s0[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2704), .CK(clk), .Q(Ciphertext_s1[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2705), .CK(clk), .Q(Ciphertext_s2[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5223), .CK(clk), .Q(Ciphertext_s0[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5225), .CK(clk), .Q(Ciphertext_s1[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5227), .CK(clk), .Q(Ciphertext_s2[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5229), .CK(clk), .Q(Ciphertext_s0[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5231), .CK(clk), .Q(Ciphertext_s1[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5233), .CK(clk), .Q(Ciphertext_s2[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[29]), .CK(clk), .Q(Ciphertext_s0[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3022), .CK(clk), .Q(Ciphertext_s1[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3023), .CK(clk), .Q(Ciphertext_s2[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[28]), .CK(clk), .Q(Ciphertext_s0[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2936), .CK(clk), .Q(Ciphertext_s1[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2937), .CK(clk), .Q(Ciphertext_s2[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5235), .CK(clk), .Q(Ciphertext_s0[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5237), .CK(clk), .Q(Ciphertext_s1[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5239), .CK(clk), .Q(Ciphertext_s2[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5241), .CK(clk), .Q(Ciphertext_s0[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5243), .CK(clk), .Q(Ciphertext_s1[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5245), .CK(clk), .Q(Ciphertext_s2[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[25]), .CK(clk), .Q(Ciphertext_s0[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3080), .CK(clk), .Q(Ciphertext_s1[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3081), .CK(clk), .Q(Ciphertext_s2[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[24]), .CK(clk), .Q(Ciphertext_s0[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3062), .CK(clk), .Q(Ciphertext_s1[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3063), .CK(clk), .Q(Ciphertext_s2[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5247), .CK(clk), .Q(Ciphertext_s0[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5249), .CK(clk), .Q(Ciphertext_s1[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5251), .CK(clk), .Q(Ciphertext_s2[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5253), .CK(clk), .Q(Ciphertext_s0[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5255), .CK(clk), .Q(Ciphertext_s1[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5257), .CK(clk), .Q(Ciphertext_s2[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[21]), .CK(clk), .Q(Ciphertext_s0[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3014), .CK(clk), .Q(Ciphertext_s1[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3015), .CK(clk), .Q(Ciphertext_s2[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[20]), .CK(clk), .Q(Ciphertext_s0[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2928), .CK(clk), .Q(Ciphertext_s1[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2929), .CK(clk), .Q(Ciphertext_s2[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5259), .CK(clk), .Q(Ciphertext_s0[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5261), .CK(clk), .Q(Ciphertext_s1[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5263), .CK(clk), .Q(Ciphertext_s2[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5265), .CK(clk), .Q(Ciphertext_s0[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5267), .CK(clk), .Q(Ciphertext_s1[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5269), .CK(clk), .Q(Ciphertext_s2[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[17]), .CK(clk), .Q(Ciphertext_s0[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3010), .CK(clk), .Q(Ciphertext_s1[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3011), .CK(clk), .Q(Ciphertext_s2[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[16]), .CK(clk), .Q(Ciphertext_s0[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2924), .CK(clk), .Q(Ciphertext_s1[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2925), .CK(clk), .Q(Ciphertext_s2[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5271), .CK(clk), .Q(Ciphertext_s0[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5273), .CK(clk), .Q(Ciphertext_s1[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5275), .CK(clk), .Q(Ciphertext_s2[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5277), .CK(clk), .Q(Ciphertext_s0[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5279), .CK(clk), .Q(Ciphertext_s1[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5281), .CK(clk), .Q(Ciphertext_s2[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[13]), .CK(clk), .Q(Ciphertext_s0[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3076), .CK(clk), .Q(Ciphertext_s1[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3077), .CK(clk), .Q(Ciphertext_s2[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[12]), .CK(clk), .Q(Ciphertext_s0[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3058), .CK(clk), .Q(Ciphertext_s1[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3059), .CK(clk), .Q(Ciphertext_s2[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5283), .CK(clk), .Q(Ciphertext_s0[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5285), .CK(clk), .Q(Ciphertext_s1[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5287), .CK(clk), .Q(Ciphertext_s2[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5289), .CK(clk), .Q(Ciphertext_s0[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5291), .CK(clk), .Q(Ciphertext_s1[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5293), .CK(clk), .Q(Ciphertext_s2[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[9]), .CK(clk), .Q(Ciphertext_s0[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_3002), .CK(clk), .Q(Ciphertext_s1[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_3003), .CK(clk), .Q(Ciphertext_s2[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[8]), .CK(clk), .Q(Ciphertext_s0[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2916), .CK(clk), .Q(Ciphertext_s1[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2917), .CK(clk), .Q(Ciphertext_s2[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5295), .CK(clk), .Q(Ciphertext_s0[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5297), .CK(clk), .Q(Ciphertext_s1[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5299), .CK(clk), .Q(Ciphertext_s2[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5301), .CK(clk), .Q(Ciphertext_s0[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5303), .CK(clk), .Q(Ciphertext_s1[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5305), .CK(clk), .Q(Ciphertext_s2[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[5]), .CK(clk), .Q(Ciphertext_s0[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2998), .CK(clk), .Q(Ciphertext_s1[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2999), .CK(clk), .Q(Ciphertext_s2[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[4]), .CK(clk), .Q(Ciphertext_s0[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2912), .CK(clk), .Q(Ciphertext_s1[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2913), .CK(clk), .Q(Ciphertext_s2[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5307), .CK(clk), .Q(Ciphertext_s0[3]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5309), .CK(clk), .Q(Ciphertext_s1[3]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5311), .CK(clk), .Q(Ciphertext_s2[3]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5313), .CK(clk), .Q(Ciphertext_s0[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5315), .CK(clk), .Q(Ciphertext_s1[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5317), .CK(clk), .Q(Ciphertext_s2[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[1]), .CK(clk), .Q(Ciphertext_s0[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2994), .CK(clk), .Q(Ciphertext_s1[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2995), .CK(clk), .Q(Ciphertext_s2[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_0__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[0]), .CK(clk), .Q(Ciphertext_s0[0]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_0__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2908), .CK(clk), .Q(Ciphertext_s1[0]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_0__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_2909), .CK(clk), .Q(Ciphertext_s2[0]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5321), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[31]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5325), .CK(clk), .Q(new_AGEMA_signal_1542), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5329), .CK(clk), .Q(new_AGEMA_signal_1543), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5333), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[30]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5337), .CK(clk), .Q(new_AGEMA_signal_1536), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5341), .CK(clk), .Q(new_AGEMA_signal_1537), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5345), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[29]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5349), .CK(clk), .Q(new_AGEMA_signal_1530), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5353), .CK(clk), .Q(new_AGEMA_signal_1531), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5357), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[28]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5361), .CK(clk), .Q(new_AGEMA_signal_1524), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5365), .CK(clk), .Q(new_AGEMA_signal_1525), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5369), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[27]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5373), .CK(clk), .Q(new_AGEMA_signal_1518), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5377), .CK(clk), .Q(new_AGEMA_signal_1519), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5381), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[26]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5385), .CK(clk), .Q(new_AGEMA_signal_1512), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5389), .CK(clk), .Q(new_AGEMA_signal_1513), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5393), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[25]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5397), .CK(clk), .Q(new_AGEMA_signal_1506), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5401), .CK(clk), .Q(new_AGEMA_signal_1507), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5405), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[24]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5409), .CK(clk), .Q(new_AGEMA_signal_1500), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5413), .CK(clk), .Q(new_AGEMA_signal_1501), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5417), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[23]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5421), .CK(clk), .Q(new_AGEMA_signal_1494), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5425), .CK(clk), .Q(new_AGEMA_signal_1495), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5429), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[22]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5433), .CK(clk), .Q(new_AGEMA_signal_1488), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5437), .CK(clk), .Q(new_AGEMA_signal_1489), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5441), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[21]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5445), .CK(clk), .Q(new_AGEMA_signal_1482), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5449), .CK(clk), .Q(new_AGEMA_signal_1483), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5453), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[20]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5457), .CK(clk), .Q(new_AGEMA_signal_1476), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5461), .CK(clk), .Q(new_AGEMA_signal_1477), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5465), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[19]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5469), .CK(clk), .Q(new_AGEMA_signal_1470), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5473), .CK(clk), .Q(new_AGEMA_signal_1471), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5477), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[18]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5481), .CK(clk), .Q(new_AGEMA_signal_1464), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5485), .CK(clk), .Q(new_AGEMA_signal_1465), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5489), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[17]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5493), .CK(clk), .Q(new_AGEMA_signal_1458), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5497), .CK(clk), .Q(new_AGEMA_signal_1459), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5501), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[16]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5505), .CK(clk), .Q(new_AGEMA_signal_1452), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5509), .CK(clk), .Q(new_AGEMA_signal_1453), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5513), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[15]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5517), .CK(clk), .Q(new_AGEMA_signal_1446), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5521), .CK(clk), .Q(new_AGEMA_signal_1447), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5525), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[14]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5529), .CK(clk), .Q(new_AGEMA_signal_1440), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5533), .CK(clk), .Q(new_AGEMA_signal_1441), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5537), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[13]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5541), .CK(clk), .Q(new_AGEMA_signal_1434), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5545), .CK(clk), .Q(new_AGEMA_signal_1435), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5549), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[12]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5553), .CK(clk), .Q(new_AGEMA_signal_1428), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5557), .CK(clk), .Q(new_AGEMA_signal_1429), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5561), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[11]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5565), .CK(clk), .Q(new_AGEMA_signal_1422), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5569), .CK(clk), .Q(new_AGEMA_signal_1423), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5573), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[10]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5577), .CK(clk), .Q(new_AGEMA_signal_1416), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5581), .CK(clk), .Q(new_AGEMA_signal_1417), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5585), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[9]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5589), .CK(clk), .Q(new_AGEMA_signal_1410), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5593), .CK(clk), .Q(new_AGEMA_signal_1411), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5597), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[8]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5601), .CK(clk), .Q(new_AGEMA_signal_1404), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5605), .CK(clk), .Q(new_AGEMA_signal_1405), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5609), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[7]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5613), .CK(clk), .Q(new_AGEMA_signal_1398), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5617), .CK(clk), .Q(new_AGEMA_signal_1399), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5621), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[6]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5625), .CK(clk), .Q(new_AGEMA_signal_1392), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5629), .CK(clk), .Q(new_AGEMA_signal_1393), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5633), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[5]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5637), .CK(clk), .Q(new_AGEMA_signal_1386), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5641), .CK(clk), .Q(new_AGEMA_signal_1387), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5645), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[4]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5649), .CK(clk), .Q(new_AGEMA_signal_1380), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5653), .CK(clk), .Q(new_AGEMA_signal_1381), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5657), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[3]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5661), .CK(clk), .Q(new_AGEMA_signal_1374), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5665), .CK(clk), .Q(new_AGEMA_signal_1375), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5669), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[2]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5673), .CK(clk), .Q(new_AGEMA_signal_1368), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5677), .CK(clk), .Q(new_AGEMA_signal_1369), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5681), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[1]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5685), .CK(clk), .Q(new_AGEMA_signal_1362), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5689), .CK(clk), .Q(new_AGEMA_signal_1363), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5693), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[0]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5697), .CK(clk), .Q(new_AGEMA_signal_1356), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5701), .CK(clk), .Q(new_AGEMA_signal_1357), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5705), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[55]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5709), .CK(clk), .Q(new_AGEMA_signal_1686), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5713), .CK(clk), .Q(new_AGEMA_signal_1687), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5717), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[54]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5721), .CK(clk), .Q(new_AGEMA_signal_1680), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5725), .CK(clk), .Q(new_AGEMA_signal_1681), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5729), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[53]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5733), .CK(clk), .Q(new_AGEMA_signal_1674), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5737), .CK(clk), .Q(new_AGEMA_signal_1675), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5741), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[52]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5745), .CK(clk), .Q(new_AGEMA_signal_1668), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5749), .CK(clk), .Q(new_AGEMA_signal_1669), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5753), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[63]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5757), .CK(clk), .Q(new_AGEMA_signal_1734), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5761), .CK(clk), .Q(new_AGEMA_signal_1735), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5765), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[62]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5769), .CK(clk), .Q(new_AGEMA_signal_1728), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5773), .CK(clk), .Q(new_AGEMA_signal_1729), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5777), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[61]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5781), .CK(clk), .Q(new_AGEMA_signal_1722), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5785), .CK(clk), .Q(new_AGEMA_signal_1723), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5789), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[60]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5793), .CK(clk), .Q(new_AGEMA_signal_1716), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5797), .CK(clk), .Q(new_AGEMA_signal_1717), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5801), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[47]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5805), .CK(clk), .Q(new_AGEMA_signal_1638), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5809), .CK(clk), .Q(new_AGEMA_signal_1639), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5813), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[46]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5817), .CK(clk), .Q(new_AGEMA_signal_1632), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5821), .CK(clk), .Q(new_AGEMA_signal_1633), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5825), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[45]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5829), .CK(clk), .Q(new_AGEMA_signal_1626), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5833), .CK(clk), .Q(new_AGEMA_signal_1627), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5837), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[44]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5841), .CK(clk), .Q(new_AGEMA_signal_1620), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5845), .CK(clk), .Q(new_AGEMA_signal_1621), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5849), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[35]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5853), .CK(clk), .Q(new_AGEMA_signal_1566), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5857), .CK(clk), .Q(new_AGEMA_signal_1567), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5861), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[34]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5865), .CK(clk), .Q(new_AGEMA_signal_1560), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5869), .CK(clk), .Q(new_AGEMA_signal_1561), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5873), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[33]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5877), .CK(clk), .Q(new_AGEMA_signal_1554), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5881), .CK(clk), .Q(new_AGEMA_signal_1555), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5885), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[32]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5889), .CK(clk), .Q(new_AGEMA_signal_1548), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5893), .CK(clk), .Q(new_AGEMA_signal_1549), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5897), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[39]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5901), .CK(clk), .Q(new_AGEMA_signal_1590), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5905), .CK(clk), .Q(new_AGEMA_signal_1591), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5909), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[38]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5913), .CK(clk), .Q(new_AGEMA_signal_1584), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5917), .CK(clk), .Q(new_AGEMA_signal_1585), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5921), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[37]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5925), .CK(clk), .Q(new_AGEMA_signal_1578), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5929), .CK(clk), .Q(new_AGEMA_signal_1579), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5933), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[36]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5937), .CK(clk), .Q(new_AGEMA_signal_1572), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5941), .CK(clk), .Q(new_AGEMA_signal_1573), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5945), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[51]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5949), .CK(clk), .Q(new_AGEMA_signal_1662), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5953), .CK(clk), .Q(new_AGEMA_signal_1663), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5957), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[50]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5961), .CK(clk), .Q(new_AGEMA_signal_1656), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5965), .CK(clk), .Q(new_AGEMA_signal_1657), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5969), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[49]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5973), .CK(clk), .Q(new_AGEMA_signal_1650), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5977), .CK(clk), .Q(new_AGEMA_signal_1651), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5981), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[48]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5985), .CK(clk), .Q(new_AGEMA_signal_1644), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_5989), .CK(clk), .Q(new_AGEMA_signal_1645), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_5993), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[43]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_5997), .CK(clk), .Q(new_AGEMA_signal_1614), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6001), .CK(clk), .Q(new_AGEMA_signal_1615), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6005), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[42]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6009), .CK(clk), .Q(new_AGEMA_signal_1608), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6013), .CK(clk), .Q(new_AGEMA_signal_1609), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6017), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[41]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6021), .CK(clk), .Q(new_AGEMA_signal_1602), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6025), .CK(clk), .Q(new_AGEMA_signal_1603), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6029), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[40]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6033), .CK(clk), .Q(new_AGEMA_signal_1596), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6037), .CK(clk), .Q(new_AGEMA_signal_1597), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6041), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[59]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6045), .CK(clk), .Q(new_AGEMA_signal_1710), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6049), .CK(clk), .Q(new_AGEMA_signal_1711), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6053), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[58]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6057), .CK(clk), .Q(new_AGEMA_signal_1704), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6061), .CK(clk), .Q(new_AGEMA_signal_1705), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6065), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[57]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6069), .CK(clk), .Q(new_AGEMA_signal_1698), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6073), .CK(clk), .Q(new_AGEMA_signal_1699), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(new_AGEMA_signal_6077), .CK(clk), .Q(
        TweakeyGeneration_key_Feedback[56]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_6081), .CK(clk), .Q(new_AGEMA_signal_1692), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF_s_reg_2_s_current_state_reg ( 
        .D(new_AGEMA_signal_6085), .CK(clk), .Q(new_AGEMA_signal_1693), .QN()
         );
endmodule

