////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module AES in file /AGEMA/Designs/AES_serial/AGEMA/sbox_opt3/AES.v */
/* clock gating is added to the circuit, the latency increased 4 time(s)  */

module AES_HPC3_ClockGating_d1 (plaintext_s0, key_s0, clk, start, plaintext_s1, key_s1, Fresh, ciphertext_s0, done, ciphertext_s1, Synch);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input start ;
    input [127:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [67:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output Synch ;
    wire nReset ;
    wire selMC ;
    wire selSR ;
    wire selXOR ;
    wire enRCon ;
    wire finalStep ;
    wire intFinal ;
    wire intselXOR ;
    wire notFirst ;
    wire n10 ;
    wire n9 ;
    wire n12 ;
    wire n13 ;
    wire ctrl_n16 ;
    wire ctrl_n15 ;
    wire ctrl_n14 ;
    wire ctrl_n11 ;
    wire ctrl_n10 ;
    wire ctrl_n9 ;
    wire ctrl_n8 ;
    wire ctrl_n7 ;
    wire ctrl_n5 ;
    wire ctrl_n4 ;
    wire ctrl_n2 ;
    wire ctrl_n12 ;
    wire ctrl_n6 ;
    wire ctrl_N14 ;
    wire ctrl_seq4Out_1_ ;
    wire ctrl_seq4In_1_ ;
    wire ctrl_nRstSeq4 ;
    wire ctrl_n13 ;
    wire ctrl_seq6Out_4_ ;
    wire ctrl_seq6In_1_ ;
    wire ctrl_seq6In_2_ ;
    wire ctrl_seq6In_3_ ;
    wire ctrl_seq6In_4_ ;
    wire ctrl_seq6_SFF_0_QD ;
    wire ctrl_seq6_SFF_1_QD ;
    wire ctrl_seq6_SFF_2_QD ;
    wire ctrl_seq6_SFF_3_QD ;
    wire ctrl_seq6_SFF_4_QD ;
    wire ctrl_seq4_SFF_0_QD ;
    wire ctrl_seq4_SFF_1_QD ;
    wire stateArray_n33 ;
    wire stateArray_n32 ;
    wire stateArray_n31 ;
    wire stateArray_n30 ;
    wire stateArray_n29 ;
    wire stateArray_n28 ;
    wire stateArray_n27 ;
    wire stateArray_n26 ;
    wire stateArray_n25 ;
    wire stateArray_n24 ;
    wire stateArray_n23 ;
    wire stateArray_n22 ;
    wire stateArray_n21 ;
    wire stateArray_n20 ;
    wire stateArray_n19 ;
    wire stateArray_n18 ;
    wire stateArray_n17 ;
    wire stateArray_n16 ;
    wire stateArray_n15 ;
    wire stateArray_n14 ;
    wire stateArray_n13 ;
    wire stateArray_S00reg_gff_1_SFF_0_QD ;
    wire stateArray_S00reg_gff_1_SFF_1_QD ;
    wire stateArray_S00reg_gff_1_SFF_2_QD ;
    wire stateArray_S00reg_gff_1_SFF_3_QD ;
    wire stateArray_S00reg_gff_1_SFF_4_QD ;
    wire stateArray_S00reg_gff_1_SFF_5_QD ;
    wire stateArray_S00reg_gff_1_SFF_6_QD ;
    wire stateArray_S00reg_gff_1_SFF_7_QD ;
    wire stateArray_S01reg_gff_1_SFF_0_QD ;
    wire stateArray_S01reg_gff_1_SFF_1_QD ;
    wire stateArray_S01reg_gff_1_SFF_2_QD ;
    wire stateArray_S01reg_gff_1_SFF_3_QD ;
    wire stateArray_S01reg_gff_1_SFF_4_QD ;
    wire stateArray_S01reg_gff_1_SFF_5_QD ;
    wire stateArray_S01reg_gff_1_SFF_6_QD ;
    wire stateArray_S01reg_gff_1_SFF_7_QD ;
    wire stateArray_S02reg_gff_1_SFF_0_QD ;
    wire stateArray_S02reg_gff_1_SFF_1_QD ;
    wire stateArray_S02reg_gff_1_SFF_2_QD ;
    wire stateArray_S02reg_gff_1_SFF_3_QD ;
    wire stateArray_S02reg_gff_1_SFF_4_QD ;
    wire stateArray_S02reg_gff_1_SFF_5_QD ;
    wire stateArray_S02reg_gff_1_SFF_6_QD ;
    wire stateArray_S02reg_gff_1_SFF_7_QD ;
    wire stateArray_S03reg_gff_1_SFF_0_QD ;
    wire stateArray_S03reg_gff_1_SFF_1_QD ;
    wire stateArray_S03reg_gff_1_SFF_2_QD ;
    wire stateArray_S03reg_gff_1_SFF_3_QD ;
    wire stateArray_S03reg_gff_1_SFF_4_QD ;
    wire stateArray_S03reg_gff_1_SFF_5_QD ;
    wire stateArray_S03reg_gff_1_SFF_6_QD ;
    wire stateArray_S03reg_gff_1_SFF_7_QD ;
    wire stateArray_S10reg_gff_1_SFF_0_QD ;
    wire stateArray_S10reg_gff_1_SFF_1_QD ;
    wire stateArray_S10reg_gff_1_SFF_2_QD ;
    wire stateArray_S10reg_gff_1_SFF_3_QD ;
    wire stateArray_S10reg_gff_1_SFF_4_QD ;
    wire stateArray_S10reg_gff_1_SFF_5_QD ;
    wire stateArray_S10reg_gff_1_SFF_6_QD ;
    wire stateArray_S10reg_gff_1_SFF_7_QD ;
    wire stateArray_S11reg_gff_1_SFF_0_QD ;
    wire stateArray_S11reg_gff_1_SFF_1_QD ;
    wire stateArray_S11reg_gff_1_SFF_2_QD ;
    wire stateArray_S11reg_gff_1_SFF_3_QD ;
    wire stateArray_S11reg_gff_1_SFF_4_QD ;
    wire stateArray_S11reg_gff_1_SFF_5_QD ;
    wire stateArray_S11reg_gff_1_SFF_6_QD ;
    wire stateArray_S11reg_gff_1_SFF_7_QD ;
    wire stateArray_S12reg_gff_1_SFF_0_QD ;
    wire stateArray_S12reg_gff_1_SFF_1_QD ;
    wire stateArray_S12reg_gff_1_SFF_2_QD ;
    wire stateArray_S12reg_gff_1_SFF_3_QD ;
    wire stateArray_S12reg_gff_1_SFF_4_QD ;
    wire stateArray_S12reg_gff_1_SFF_5_QD ;
    wire stateArray_S12reg_gff_1_SFF_6_QD ;
    wire stateArray_S12reg_gff_1_SFF_7_QD ;
    wire stateArray_S13reg_gff_1_SFF_0_QD ;
    wire stateArray_S13reg_gff_1_SFF_1_QD ;
    wire stateArray_S13reg_gff_1_SFF_2_QD ;
    wire stateArray_S13reg_gff_1_SFF_3_QD ;
    wire stateArray_S13reg_gff_1_SFF_4_QD ;
    wire stateArray_S13reg_gff_1_SFF_5_QD ;
    wire stateArray_S13reg_gff_1_SFF_6_QD ;
    wire stateArray_S13reg_gff_1_SFF_7_QD ;
    wire stateArray_S20reg_gff_1_SFF_0_QD ;
    wire stateArray_S20reg_gff_1_SFF_1_QD ;
    wire stateArray_S20reg_gff_1_SFF_2_QD ;
    wire stateArray_S20reg_gff_1_SFF_3_QD ;
    wire stateArray_S20reg_gff_1_SFF_4_QD ;
    wire stateArray_S20reg_gff_1_SFF_5_QD ;
    wire stateArray_S20reg_gff_1_SFF_6_QD ;
    wire stateArray_S20reg_gff_1_SFF_7_QD ;
    wire stateArray_S21reg_gff_1_SFF_0_QD ;
    wire stateArray_S21reg_gff_1_SFF_1_QD ;
    wire stateArray_S21reg_gff_1_SFF_2_QD ;
    wire stateArray_S21reg_gff_1_SFF_3_QD ;
    wire stateArray_S21reg_gff_1_SFF_4_QD ;
    wire stateArray_S21reg_gff_1_SFF_5_QD ;
    wire stateArray_S21reg_gff_1_SFF_6_QD ;
    wire stateArray_S21reg_gff_1_SFF_7_QD ;
    wire stateArray_S22reg_gff_1_SFF_0_QD ;
    wire stateArray_S22reg_gff_1_SFF_1_QD ;
    wire stateArray_S22reg_gff_1_SFF_2_QD ;
    wire stateArray_S22reg_gff_1_SFF_3_QD ;
    wire stateArray_S22reg_gff_1_SFF_4_QD ;
    wire stateArray_S22reg_gff_1_SFF_5_QD ;
    wire stateArray_S22reg_gff_1_SFF_6_QD ;
    wire stateArray_S22reg_gff_1_SFF_7_QD ;
    wire stateArray_S23reg_gff_1_SFF_0_QD ;
    wire stateArray_S23reg_gff_1_SFF_1_QD ;
    wire stateArray_S23reg_gff_1_SFF_2_QD ;
    wire stateArray_S23reg_gff_1_SFF_3_QD ;
    wire stateArray_S23reg_gff_1_SFF_4_QD ;
    wire stateArray_S23reg_gff_1_SFF_5_QD ;
    wire stateArray_S23reg_gff_1_SFF_6_QD ;
    wire stateArray_S23reg_gff_1_SFF_7_QD ;
    wire stateArray_S30reg_gff_1_SFF_0_QD ;
    wire stateArray_S30reg_gff_1_SFF_1_QD ;
    wire stateArray_S30reg_gff_1_SFF_2_QD ;
    wire stateArray_S30reg_gff_1_SFF_3_QD ;
    wire stateArray_S30reg_gff_1_SFF_4_QD ;
    wire stateArray_S30reg_gff_1_SFF_5_QD ;
    wire stateArray_S30reg_gff_1_SFF_6_QD ;
    wire stateArray_S30reg_gff_1_SFF_7_QD ;
    wire stateArray_S31reg_gff_1_SFF_0_QD ;
    wire stateArray_S31reg_gff_1_SFF_1_QD ;
    wire stateArray_S31reg_gff_1_SFF_2_QD ;
    wire stateArray_S31reg_gff_1_SFF_3_QD ;
    wire stateArray_S31reg_gff_1_SFF_4_QD ;
    wire stateArray_S31reg_gff_1_SFF_5_QD ;
    wire stateArray_S31reg_gff_1_SFF_6_QD ;
    wire stateArray_S31reg_gff_1_SFF_7_QD ;
    wire stateArray_S32reg_gff_1_SFF_0_QD ;
    wire stateArray_S32reg_gff_1_SFF_1_QD ;
    wire stateArray_S32reg_gff_1_SFF_2_QD ;
    wire stateArray_S32reg_gff_1_SFF_3_QD ;
    wire stateArray_S32reg_gff_1_SFF_4_QD ;
    wire stateArray_S32reg_gff_1_SFF_5_QD ;
    wire stateArray_S32reg_gff_1_SFF_6_QD ;
    wire stateArray_S32reg_gff_1_SFF_7_QD ;
    wire stateArray_S33reg_gff_1_SFF_0_QD ;
    wire stateArray_S33reg_gff_1_SFF_1_QD ;
    wire stateArray_S33reg_gff_1_SFF_2_QD ;
    wire stateArray_S33reg_gff_1_SFF_3_QD ;
    wire stateArray_S33reg_gff_1_SFF_4_QD ;
    wire stateArray_S33reg_gff_1_SFF_5_QD ;
    wire stateArray_S33reg_gff_1_SFF_6_QD ;
    wire stateArray_S33reg_gff_1_SFF_7_QD ;
    wire MUX_StateInMC_n7 ;
    wire MUX_StateInMC_n6 ;
    wire MUX_StateInMC_n5 ;
    wire KeyArray_n55 ;
    wire KeyArray_n54 ;
    wire KeyArray_n53 ;
    wire KeyArray_n52 ;
    wire KeyArray_n51 ;
    wire KeyArray_n50 ;
    wire KeyArray_n49 ;
    wire KeyArray_n48 ;
    wire KeyArray_n47 ;
    wire KeyArray_n46 ;
    wire KeyArray_n45 ;
    wire KeyArray_n44 ;
    wire KeyArray_n43 ;
    wire KeyArray_n42 ;
    wire KeyArray_n41 ;
    wire KeyArray_n40 ;
    wire KeyArray_n39 ;
    wire KeyArray_n38 ;
    wire KeyArray_n37 ;
    wire KeyArray_n36 ;
    wire KeyArray_n35 ;
    wire KeyArray_n34 ;
    wire KeyArray_n33 ;
    wire KeyArray_n32 ;
    wire KeyArray_n31 ;
    wire KeyArray_n30 ;
    wire KeyArray_n29 ;
    wire KeyArray_n28 ;
    wire KeyArray_n27 ;
    wire KeyArray_n26 ;
    wire KeyArray_n25 ;
    wire KeyArray_n24 ;
    wire KeyArray_n23 ;
    wire KeyArray_n22 ;
    wire KeyArray_outS01ser_0_ ;
    wire KeyArray_outS01ser_1_ ;
    wire KeyArray_outS01ser_2_ ;
    wire KeyArray_outS01ser_3_ ;
    wire KeyArray_outS01ser_4_ ;
    wire KeyArray_outS01ser_5_ ;
    wire KeyArray_outS01ser_6_ ;
    wire KeyArray_outS01ser_7_ ;
    wire KeyArray_S00reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S00reg_gff_1_SFF_0_QD ;
    wire KeyArray_S00reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_1_QD ;
    wire KeyArray_S00reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_2_QD ;
    wire KeyArray_S00reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_3_QD ;
    wire KeyArray_S00reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_4_QD ;
    wire KeyArray_S00reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_5_QD ;
    wire KeyArray_S00reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_6_QD ;
    wire KeyArray_S00reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_7_QD ;
    wire KeyArray_S01reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_0_QD ;
    wire KeyArray_S01reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_1_QD ;
    wire KeyArray_S01reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_2_QD ;
    wire KeyArray_S01reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_3_QD ;
    wire KeyArray_S01reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_4_QD ;
    wire KeyArray_S01reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_5_QD ;
    wire KeyArray_S01reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_6_QD ;
    wire KeyArray_S01reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_7_QD ;
    wire KeyArray_S02reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_0_QD ;
    wire KeyArray_S02reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_1_QD ;
    wire KeyArray_S02reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_2_QD ;
    wire KeyArray_S02reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_3_QD ;
    wire KeyArray_S02reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_4_QD ;
    wire KeyArray_S02reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_5_QD ;
    wire KeyArray_S02reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_6_QD ;
    wire KeyArray_S02reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_7_QD ;
    wire KeyArray_S03reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_0_QD ;
    wire KeyArray_S03reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_1_QD ;
    wire KeyArray_S03reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_2_QD ;
    wire KeyArray_S03reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_3_QD ;
    wire KeyArray_S03reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_4_QD ;
    wire KeyArray_S03reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S03reg_gff_1_SFF_5_QD ;
    wire KeyArray_S03reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S03reg_gff_1_SFF_6_QD ;
    wire KeyArray_S03reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S03reg_gff_1_SFF_7_QD ;
    wire KeyArray_S10reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_0_QD ;
    wire KeyArray_S10reg_gff_1_SFF_1_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_1_QD ;
    wire KeyArray_S10reg_gff_1_SFF_2_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_2_QD ;
    wire KeyArray_S10reg_gff_1_SFF_3_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_3_QD ;
    wire KeyArray_S10reg_gff_1_SFF_4_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_4_QD ;
    wire KeyArray_S10reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_5_QD ;
    wire KeyArray_S10reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_6_QD ;
    wire KeyArray_S10reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_7_QD ;
    wire KeyArray_S11reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_0_QD ;
    wire KeyArray_S11reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_1_QD ;
    wire KeyArray_S11reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_2_QD ;
    wire KeyArray_S11reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_3_QD ;
    wire KeyArray_S11reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_4_QD ;
    wire KeyArray_S11reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_5_QD ;
    wire KeyArray_S11reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_6_QD ;
    wire KeyArray_S11reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_7_QD ;
    wire KeyArray_S12reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_0_QD ;
    wire KeyArray_S12reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_1_QD ;
    wire KeyArray_S12reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_2_QD ;
    wire KeyArray_S12reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_3_QD ;
    wire KeyArray_S12reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_4_QD ;
    wire KeyArray_S12reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_5_QD ;
    wire KeyArray_S12reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_6_QD ;
    wire KeyArray_S12reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_7_QD ;
    wire KeyArray_S13reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_0_QD ;
    wire KeyArray_S13reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_1_QD ;
    wire KeyArray_S13reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_2_QD ;
    wire KeyArray_S13reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_3_QD ;
    wire KeyArray_S13reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_4_QD ;
    wire KeyArray_S13reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S13reg_gff_1_SFF_5_QD ;
    wire KeyArray_S13reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S13reg_gff_1_SFF_6_QD ;
    wire KeyArray_S13reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S13reg_gff_1_SFF_7_QD ;
    wire KeyArray_S20reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_0_QD ;
    wire KeyArray_S20reg_gff_1_SFF_1_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_1_QD ;
    wire KeyArray_S20reg_gff_1_SFF_2_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_2_QD ;
    wire KeyArray_S20reg_gff_1_SFF_3_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_3_QD ;
    wire KeyArray_S20reg_gff_1_SFF_4_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_4_QD ;
    wire KeyArray_S20reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_5_QD ;
    wire KeyArray_S20reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_6_QD ;
    wire KeyArray_S20reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_7_QD ;
    wire KeyArray_S21reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_0_QD ;
    wire KeyArray_S21reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_1_QD ;
    wire KeyArray_S21reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_2_QD ;
    wire KeyArray_S21reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_3_QD ;
    wire KeyArray_S21reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_4_QD ;
    wire KeyArray_S21reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_5_QD ;
    wire KeyArray_S21reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_6_QD ;
    wire KeyArray_S21reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_7_QD ;
    wire KeyArray_S22reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_0_QD ;
    wire KeyArray_S22reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_1_QD ;
    wire KeyArray_S22reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_2_QD ;
    wire KeyArray_S22reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_3_QD ;
    wire KeyArray_S22reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_4_QD ;
    wire KeyArray_S22reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_5_QD ;
    wire KeyArray_S22reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_6_QD ;
    wire KeyArray_S22reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_7_QD ;
    wire KeyArray_S23reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_0_QD ;
    wire KeyArray_S23reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_1_QD ;
    wire KeyArray_S23reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_2_QD ;
    wire KeyArray_S23reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_3_QD ;
    wire KeyArray_S23reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_4_QD ;
    wire KeyArray_S23reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S23reg_gff_1_SFF_5_QD ;
    wire KeyArray_S23reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S23reg_gff_1_SFF_6_QD ;
    wire KeyArray_S23reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S23reg_gff_1_SFF_7_QD ;
    wire KeyArray_S30reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_0_QD ;
    wire KeyArray_S30reg_gff_1_SFF_1_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_1_QD ;
    wire KeyArray_S30reg_gff_1_SFF_2_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_2_QD ;
    wire KeyArray_S30reg_gff_1_SFF_3_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_3_QD ;
    wire KeyArray_S30reg_gff_1_SFF_4_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_4_QD ;
    wire KeyArray_S30reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_5_QD ;
    wire KeyArray_S30reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_6_QD ;
    wire KeyArray_S30reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_7_QD ;
    wire KeyArray_S31reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_0_QD ;
    wire KeyArray_S31reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_1_QD ;
    wire KeyArray_S31reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_2_QD ;
    wire KeyArray_S31reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_3_QD ;
    wire KeyArray_S31reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_4_QD ;
    wire KeyArray_S31reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_5_QD ;
    wire KeyArray_S31reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_6_QD ;
    wire KeyArray_S31reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_7_QD ;
    wire KeyArray_S32reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_0_QD ;
    wire KeyArray_S32reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_1_QD ;
    wire KeyArray_S32reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_2_QD ;
    wire KeyArray_S32reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_3_QD ;
    wire KeyArray_S32reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_4_QD ;
    wire KeyArray_S32reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_5_QD ;
    wire KeyArray_S32reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S32reg_gff_1_SFF_6_QD ;
    wire KeyArray_S32reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S32reg_gff_1_SFF_7_QD ;
    wire KeyArray_S33reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_0_QD ;
    wire KeyArray_S33reg_gff_1_SFF_1_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_1_QD ;
    wire KeyArray_S33reg_gff_1_SFF_2_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_2_QD ;
    wire KeyArray_S33reg_gff_1_SFF_3_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_3_QD ;
    wire KeyArray_S33reg_gff_1_SFF_4_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_4_QD ;
    wire KeyArray_S33reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_5_QD ;
    wire KeyArray_S33reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_6_QD ;
    wire KeyArray_S33reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_7_QD ;
    wire MixColumns_line0_n16 ;
    wire MixColumns_line0_n15 ;
    wire MixColumns_line0_n14 ;
    wire MixColumns_line0_n13 ;
    wire MixColumns_line0_n12 ;
    wire MixColumns_line0_n11 ;
    wire MixColumns_line0_n10 ;
    wire MixColumns_line0_n9 ;
    wire MixColumns_line0_n8 ;
    wire MixColumns_line0_n7 ;
    wire MixColumns_line0_n6 ;
    wire MixColumns_line0_n5 ;
    wire MixColumns_line0_n4 ;
    wire MixColumns_line0_n3 ;
    wire MixColumns_line0_n2 ;
    wire MixColumns_line0_n1 ;
    wire MixColumns_line1_n16 ;
    wire MixColumns_line1_n15 ;
    wire MixColumns_line1_n14 ;
    wire MixColumns_line1_n13 ;
    wire MixColumns_line1_n12 ;
    wire MixColumns_line1_n11 ;
    wire MixColumns_line1_n10 ;
    wire MixColumns_line1_n9 ;
    wire MixColumns_line1_n8 ;
    wire MixColumns_line1_n7 ;
    wire MixColumns_line1_n6 ;
    wire MixColumns_line1_n5 ;
    wire MixColumns_line1_n4 ;
    wire MixColumns_line1_n3 ;
    wire MixColumns_line1_n2 ;
    wire MixColumns_line1_n1 ;
    wire MixColumns_line1_S02_1_ ;
    wire MixColumns_line1_S02_3_ ;
    wire MixColumns_line1_S02_4_ ;
    wire MixColumns_line2_n16 ;
    wire MixColumns_line2_n15 ;
    wire MixColumns_line2_n14 ;
    wire MixColumns_line2_n13 ;
    wire MixColumns_line2_n12 ;
    wire MixColumns_line2_n11 ;
    wire MixColumns_line2_n10 ;
    wire MixColumns_line2_n9 ;
    wire MixColumns_line2_n8 ;
    wire MixColumns_line2_n7 ;
    wire MixColumns_line2_n6 ;
    wire MixColumns_line2_n5 ;
    wire MixColumns_line2_n4 ;
    wire MixColumns_line2_n3 ;
    wire MixColumns_line2_n2 ;
    wire MixColumns_line2_n1 ;
    wire MixColumns_line2_S02_1_ ;
    wire MixColumns_line2_S02_3_ ;
    wire MixColumns_line2_S02_4_ ;
    wire MixColumns_line3_n16 ;
    wire MixColumns_line3_n15 ;
    wire MixColumns_line3_n14 ;
    wire MixColumns_line3_n13 ;
    wire MixColumns_line3_n12 ;
    wire MixColumns_line3_n11 ;
    wire MixColumns_line3_n10 ;
    wire MixColumns_line3_n9 ;
    wire MixColumns_line3_n8 ;
    wire MixColumns_line3_n7 ;
    wire MixColumns_line3_n6 ;
    wire MixColumns_line3_n5 ;
    wire MixColumns_line3_n4 ;
    wire MixColumns_line3_n3 ;
    wire MixColumns_line3_n2 ;
    wire MixColumns_line3_n1 ;
    wire MixColumns_line3_S02_1_ ;
    wire MixColumns_line3_S02_3_ ;
    wire MixColumns_line3_S02_4_ ;
    wire MixColumns_line3_timesTHREE_input2_1_ ;
    wire MixColumns_line3_timesTHREE_input2_3_ ;
    wire MixColumns_line3_timesTHREE_input2_4_ ;
    wire calcRCon_n38 ;
    wire calcRCon_n37 ;
    wire calcRCon_n36 ;
    wire calcRCon_n35 ;
    wire calcRCon_n34 ;
    wire calcRCon_n33 ;
    wire calcRCon_n32 ;
    wire calcRCon_n31 ;
    wire calcRCon_n30 ;
    wire calcRCon_n29 ;
    wire calcRCon_n28 ;
    wire calcRCon_n27 ;
    wire calcRCon_n26 ;
    wire calcRCon_n25 ;
    wire calcRCon_n24 ;
    wire calcRCon_n23 ;
    wire calcRCon_n22 ;
    wire calcRCon_n21 ;
    wire calcRCon_n20 ;
    wire calcRCon_n19 ;
    wire calcRCon_n18 ;
    wire calcRCon_n17 ;
    wire calcRCon_n10 ;
    wire calcRCon_n9 ;
    wire calcRCon_n8 ;
    wire calcRCon_n7 ;
    wire calcRCon_n6 ;
    wire calcRCon_n5 ;
    wire calcRCon_n3 ;
    wire calcRCon_n11 ;
    wire calcRCon_n44 ;
    wire calcRCon_n16 ;
    wire calcRCon_n45 ;
    wire calcRCon_n46 ;
    wire calcRCon_n47 ;
    wire calcRCon_n15 ;
    wire calcRCon_n48 ;
    wire calcRCon_n12 ;
    wire calcRCon_n49 ;
    wire calcRCon_n14 ;
    wire calcRCon_n50 ;
    wire calcRCon_n13 ;
    wire calcRCon_s_current_state_0_ ;
    wire calcRCon_s_current_state_1_ ;
    wire calcRCon_s_current_state_2_ ;
    wire calcRCon_s_current_state_3_ ;
    wire calcRCon_s_current_state_4_ ;
    wire calcRCon_s_current_state_5_ ;
    wire calcRCon_s_current_state_6_ ;
    wire calcRCon_n51 ;
    wire Inst_bSbox_L29 ;
    wire Inst_bSbox_L28 ;
    wire Inst_bSbox_L27 ;
    wire Inst_bSbox_L26 ;
    wire Inst_bSbox_L25 ;
    wire Inst_bSbox_L24 ;
    wire Inst_bSbox_L23 ;
    wire Inst_bSbox_L22 ;
    wire Inst_bSbox_L21 ;
    wire Inst_bSbox_L20 ;
    wire Inst_bSbox_L19 ;
    wire Inst_bSbox_L18 ;
    wire Inst_bSbox_L17 ;
    wire Inst_bSbox_L16 ;
    wire Inst_bSbox_L15 ;
    wire Inst_bSbox_L14 ;
    wire Inst_bSbox_L13 ;
    wire Inst_bSbox_L12 ;
    wire Inst_bSbox_L11 ;
    wire Inst_bSbox_L10 ;
    wire Inst_bSbox_L9 ;
    wire Inst_bSbox_L8 ;
    wire Inst_bSbox_L7 ;
    wire Inst_bSbox_L6 ;
    wire Inst_bSbox_L5 ;
    wire Inst_bSbox_L4 ;
    wire Inst_bSbox_L3 ;
    wire Inst_bSbox_L2 ;
    wire Inst_bSbox_L1 ;
    wire Inst_bSbox_L0 ;
    wire Inst_bSbox_M63 ;
    wire Inst_bSbox_M62 ;
    wire Inst_bSbox_M61 ;
    wire Inst_bSbox_M60 ;
    wire Inst_bSbox_M59 ;
    wire Inst_bSbox_M58 ;
    wire Inst_bSbox_M57 ;
    wire Inst_bSbox_M56 ;
    wire Inst_bSbox_M55 ;
    wire Inst_bSbox_M54 ;
    wire Inst_bSbox_M53 ;
    wire Inst_bSbox_M52 ;
    wire Inst_bSbox_M51 ;
    wire Inst_bSbox_M50 ;
    wire Inst_bSbox_M49 ;
    wire Inst_bSbox_M48 ;
    wire Inst_bSbox_M47 ;
    wire Inst_bSbox_M46 ;
    wire Inst_bSbox_M45 ;
    wire Inst_bSbox_M44 ;
    wire Inst_bSbox_M43 ;
    wire Inst_bSbox_M42 ;
    wire Inst_bSbox_M41 ;
    wire Inst_bSbox_M40 ;
    wire Inst_bSbox_M39 ;
    wire Inst_bSbox_M38 ;
    wire Inst_bSbox_M37 ;
    wire Inst_bSbox_M36 ;
    wire Inst_bSbox_M35 ;
    wire Inst_bSbox_M34 ;
    wire Inst_bSbox_M33 ;
    wire Inst_bSbox_M32 ;
    wire Inst_bSbox_M31 ;
    wire Inst_bSbox_M30 ;
    wire Inst_bSbox_M29 ;
    wire Inst_bSbox_M28 ;
    wire Inst_bSbox_M27 ;
    wire Inst_bSbox_M26 ;
    wire Inst_bSbox_M25 ;
    wire Inst_bSbox_M24 ;
    wire Inst_bSbox_M23 ;
    wire Inst_bSbox_M22 ;
    wire Inst_bSbox_M21 ;
    wire Inst_bSbox_M20 ;
    wire Inst_bSbox_M19 ;
    wire Inst_bSbox_M18 ;
    wire Inst_bSbox_M17 ;
    wire Inst_bSbox_M16 ;
    wire Inst_bSbox_M15 ;
    wire Inst_bSbox_M14 ;
    wire Inst_bSbox_M13 ;
    wire Inst_bSbox_M12 ;
    wire Inst_bSbox_M11 ;
    wire Inst_bSbox_M10 ;
    wire Inst_bSbox_M9 ;
    wire Inst_bSbox_M8 ;
    wire Inst_bSbox_M7 ;
    wire Inst_bSbox_M6 ;
    wire Inst_bSbox_M5 ;
    wire Inst_bSbox_M4 ;
    wire Inst_bSbox_M3 ;
    wire Inst_bSbox_M2 ;
    wire Inst_bSbox_M1 ;
    wire Inst_bSbox_T27 ;
    wire Inst_bSbox_T26 ;
    wire Inst_bSbox_T25 ;
    wire Inst_bSbox_T24 ;
    wire Inst_bSbox_T23 ;
    wire Inst_bSbox_T22 ;
    wire Inst_bSbox_T21 ;
    wire Inst_bSbox_T20 ;
    wire Inst_bSbox_T19 ;
    wire Inst_bSbox_T18 ;
    wire Inst_bSbox_T17 ;
    wire Inst_bSbox_T16 ;
    wire Inst_bSbox_T15 ;
    wire Inst_bSbox_T14 ;
    wire Inst_bSbox_T13 ;
    wire Inst_bSbox_T12 ;
    wire Inst_bSbox_T11 ;
    wire Inst_bSbox_T10 ;
    wire Inst_bSbox_T9 ;
    wire Inst_bSbox_T8 ;
    wire Inst_bSbox_T7 ;
    wire Inst_bSbox_T6 ;
    wire Inst_bSbox_T5 ;
    wire Inst_bSbox_T4 ;
    wire Inst_bSbox_T3 ;
    wire Inst_bSbox_T2 ;
    wire Inst_bSbox_T1 ;
    wire [7:0] SboxOut ;
    wire [7:0] StateOutXORroundKey ;
    wire [7:0] StateIn ;
    wire [31:0] StateInMC ;
    wire [31:0] MCout ;
    wire [7:0] keyStateIn ;
    wire [7:0] roundConstant ;
    wire [7:0] keySBIn ;
    wire [7:0] SboxIn ;
    wire [7:0] stateArray_input_MC ;
    wire [7:0] stateArray_outS30ser_MC ;
    wire [7:0] stateArray_outS20ser_MC ;
    wire [7:0] stateArray_outS10ser_MC ;
    wire [7:0] stateArray_inS33ser ;
    wire [7:0] stateArray_inS32ser ;
    wire [7:0] stateArray_inS31ser ;
    wire [7:0] stateArray_inS30ser ;
    wire [7:0] stateArray_inS23ser ;
    wire [7:0] stateArray_inS22ser ;
    wire [7:0] stateArray_inS21ser ;
    wire [7:0] stateArray_inS20ser ;
    wire [7:0] stateArray_inS13ser ;
    wire [7:0] stateArray_inS12ser ;
    wire [7:0] stateArray_inS11ser ;
    wire [7:0] stateArray_inS10ser ;
    wire [7:0] stateArray_inS03ser ;
    wire [7:0] stateArray_inS02ser ;
    wire [7:0] stateArray_inS01ser ;
    wire [7:0] stateArray_inS00ser ;
    wire [7:0] KeyArray_outS01ser_p ;
    wire [7:0] KeyArray_outS01ser_XOR_00 ;
    wire [7:0] KeyArray_outS33ser ;
    wire [7:0] KeyArray_inS33ser ;
    wire [7:0] KeyArray_outS32ser ;
    wire [7:0] KeyArray_inS32ser ;
    wire [7:0] KeyArray_outS31ser ;
    wire [7:0] KeyArray_inS31ser ;
    wire [7:0] KeyArray_outS30ser ;
    wire [7:0] KeyArray_inS30par ;
    wire [7:0] KeyArray_inS30ser ;
    wire [7:0] KeyArray_outS23ser ;
    wire [7:0] KeyArray_inS23ser ;
    wire [7:0] KeyArray_outS22ser ;
    wire [7:0] KeyArray_inS22ser ;
    wire [7:0] KeyArray_outS21ser ;
    wire [7:0] KeyArray_inS21ser ;
    wire [7:0] KeyArray_outS20ser ;
    wire [7:0] KeyArray_inS20ser ;
    wire [7:0] KeyArray_inS13ser ;
    wire [7:0] KeyArray_outS12ser ;
    wire [7:0] KeyArray_inS12ser ;
    wire [7:0] KeyArray_outS11ser ;
    wire [7:0] KeyArray_inS11ser ;
    wire [7:0] KeyArray_outS10ser ;
    wire [7:0] KeyArray_inS10ser ;
    wire [7:0] KeyArray_outS03ser ;
    wire [7:0] KeyArray_inS03ser ;
    wire [7:0] KeyArray_outS02ser ;
    wire [7:0] KeyArray_inS02ser ;
    wire [7:0] KeyArray_inS01ser ;
    wire [7:0] KeyArray_inS00ser ;
    wire [7:0] MixColumns_line0_S13 ;
    wire [4:1] MixColumns_line0_S02 ;
    wire [4:1] MixColumns_line0_timesTHREE_input2 ;
    wire [7:0] MixColumns_line1_S13 ;
    wire [4:1] MixColumns_line1_timesTHREE_input2 ;
    wire [7:0] MixColumns_line2_S13 ;
    wire [4:1] MixColumns_line2_timesTHREE_input2 ;
    wire [7:0] MixColumns_line3_S13 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire clk_gated ;

    /* cells in depth 0 */
    INV_X1 U28 ( .A (selSR), .ZN (n12) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) U29 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_1983, keyStateIn[0]}), .c ({new_AGEMA_signal_1984, StateOutXORroundKey[0]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) U30 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_1986, keyStateIn[1]}), .c ({new_AGEMA_signal_1987, StateOutXORroundKey[1]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) U31 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({new_AGEMA_signal_1989, keyStateIn[2]}), .c ({new_AGEMA_signal_1990, StateOutXORroundKey[2]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) U32 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({new_AGEMA_signal_1992, keyStateIn[3]}), .c ({new_AGEMA_signal_1993, StateOutXORroundKey[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) U33 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_1995, keyStateIn[4]}), .c ({new_AGEMA_signal_1996, StateOutXORroundKey[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) U34 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({new_AGEMA_signal_1998, keyStateIn[5]}), .c ({new_AGEMA_signal_1999, StateOutXORroundKey[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) U35 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({new_AGEMA_signal_2001, keyStateIn[6]}), .c ({new_AGEMA_signal_2002, StateOutXORroundKey[6]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) U36 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2004, keyStateIn[7]}), .c ({new_AGEMA_signal_2005, StateOutXORroundKey[7]}) ) ;
    NAND2_X1 U37 ( .A1 (intFinal), .A2 (finalStep), .ZN (n13) ) ;
    NOR2_X1 U38 ( .A1 (n10), .A2 (n13), .ZN (done) ) ;
    AND2_X1 U39 ( .A1 (notFirst), .A2 (selXOR), .ZN (intselXOR) ) ;
    INV_X1 U40 ( .A (start), .ZN (n9) ) ;
    NOR2_X1 ctrl_U20 ( .A1 (ctrl_n16), .A2 (ctrl_n4), .ZN (ctrl_nRstSeq4) ) ;
    XNOR2_X1 ctrl_U19 ( .A (ctrl_seq6Out_4_), .B (ctrl_seq6In_1_), .ZN (ctrl_n13) ) ;
    NOR2_X1 ctrl_U18 ( .A1 (ctrl_n15), .A2 (ctrl_n14), .ZN (finalStep) ) ;
    NAND2_X1 ctrl_U17 ( .A1 (ctrl_seq4In_1_), .A2 (ctrl_n2), .ZN (ctrl_n14) ) ;
    INV_X1 ctrl_U16 ( .A (ctrl_n16), .ZN (ctrl_n15) ) ;
    INV_X1 ctrl_U15 ( .A (ctrl_seq4Out_1_), .ZN (ctrl_n2) ) ;
    NAND2_X1 ctrl_U14 ( .A1 (ctrl_n11), .A2 (ctrl_n10), .ZN (ctrl_N14) ) ;
    NAND2_X1 ctrl_U13 ( .A1 (selXOR), .A2 (ctrl_n6), .ZN (ctrl_n11) ) ;
    NOR2_X1 ctrl_U12 ( .A1 (ctrl_seq6In_3_), .A2 (ctrl_seq6Out_4_), .ZN (ctrl_n7) ) ;
    NOR2_X1 ctrl_U11 ( .A1 (ctrl_seq6In_1_), .A2 (ctrl_seq6In_4_), .ZN (ctrl_n8) ) ;
    NOR2_X1 ctrl_U10 ( .A1 (ctrl_n4), .A2 (ctrl_n5), .ZN (selXOR) ) ;
    NOR2_X1 ctrl_U9 ( .A1 (ctrl_seq4Out_1_), .A2 (ctrl_seq4In_1_), .ZN (ctrl_n5) ) ;
    INV_X1 ctrl_U8 ( .A (nReset), .ZN (ctrl_n4) ) ;
    NAND2_X1 ctrl_U7 ( .A1 (ctrl_n8), .A2 (ctrl_n7), .ZN (ctrl_n9) ) ;
    NOR2_X1 ctrl_U6 ( .A1 (ctrl_seq6In_2_), .A2 (ctrl_n9), .ZN (ctrl_n16) ) ;
    NAND2_X1 ctrl_U5 ( .A1 (nReset), .A2 (ctrl_n16), .ZN (ctrl_n10) ) ;
    INV_X1 ctrl_U4 ( .A (ctrl_n10), .ZN (selSR) ) ;
    NOR2_X1 ctrl_U3 ( .A1 (ctrl_n12), .A2 (ctrl_n4), .ZN (selMC) ) ;
    MUX2_X1 ctrl_seq6_SFF_0_MUXInst_U1 ( .S (nReset), .A (1'b1), .B (ctrl_n13), .Z (ctrl_seq6_SFF_0_QD) ) ;
    MUX2_X1 ctrl_seq6_SFF_1_MUXInst_U1 ( .S (nReset), .A (1'b0), .B (ctrl_seq6In_1_), .Z (ctrl_seq6_SFF_1_QD) ) ;
    MUX2_X1 ctrl_seq6_SFF_2_MUXInst_U1 ( .S (nReset), .A (1'b1), .B (ctrl_seq6In_2_), .Z (ctrl_seq6_SFF_2_QD) ) ;
    MUX2_X1 ctrl_seq6_SFF_3_MUXInst_U1 ( .S (nReset), .A (1'b0), .B (ctrl_seq6In_3_), .Z (ctrl_seq6_SFF_3_QD) ) ;
    MUX2_X1 ctrl_seq6_SFF_4_MUXInst_U1 ( .S (nReset), .A (1'b1), .B (ctrl_seq6In_4_), .Z (ctrl_seq6_SFF_4_QD) ) ;
    MUX2_X1 ctrl_seq4_SFF_0_MUXInst_U1 ( .S (ctrl_nRstSeq4), .A (1'b1), .B (ctrl_n2), .Z (ctrl_seq4_SFF_0_QD) ) ;
    MUX2_X1 ctrl_seq4_SFF_1_MUXInst_U1 ( .S (ctrl_nRstSeq4), .A (1'b0), .B (ctrl_seq4In_1_), .Z (ctrl_seq4_SFF_1_QD) ) ;
    INV_X1 ctrl_CSselMC_reg_U1 ( .A (ctrl_n6), .ZN (ctrl_n12) ) ;
    INV_X1 stateArray_U21 ( .A (selMC), .ZN (stateArray_n24) ) ;
    INV_X1 stateArray_U20 ( .A (stateArray_n24), .ZN (stateArray_n22) ) ;
    INV_X1 stateArray_U19 ( .A (nReset), .ZN (stateArray_n33) ) ;
    INV_X1 stateArray_U18 ( .A (stateArray_n33), .ZN (stateArray_n25) ) ;
    INV_X1 stateArray_U17 ( .A (stateArray_n21), .ZN (stateArray_n13) ) ;
    INV_X1 stateArray_U16 ( .A (stateArray_n24), .ZN (stateArray_n23) ) ;
    INV_X1 stateArray_U15 ( .A (stateArray_n33), .ZN (stateArray_n29) ) ;
    INV_X1 stateArray_U14 ( .A (stateArray_n21), .ZN (stateArray_n17) ) ;
    INV_X1 stateArray_U13 ( .A (stateArray_n33), .ZN (stateArray_n31) ) ;
    INV_X1 stateArray_U12 ( .A (stateArray_n21), .ZN (stateArray_n19) ) ;
    INV_X1 stateArray_U11 ( .A (stateArray_n33), .ZN (stateArray_n27) ) ;
    INV_X1 stateArray_U10 ( .A (stateArray_n21), .ZN (stateArray_n15) ) ;
    INV_X1 stateArray_U9 ( .A (stateArray_n33), .ZN (stateArray_n32) ) ;
    INV_X1 stateArray_U8 ( .A (stateArray_n21), .ZN (stateArray_n20) ) ;
    INV_X1 stateArray_U7 ( .A (stateArray_n33), .ZN (stateArray_n30) ) ;
    INV_X1 stateArray_U6 ( .A (stateArray_n21), .ZN (stateArray_n18) ) ;
    INV_X1 stateArray_U5 ( .A (stateArray_n33), .ZN (stateArray_n28) ) ;
    INV_X1 stateArray_U4 ( .A (stateArray_n21), .ZN (stateArray_n16) ) ;
    INV_X1 stateArray_U3 ( .A (stateArray_n33), .ZN (stateArray_n26) ) ;
    INV_X1 stateArray_U2 ( .A (stateArray_n21), .ZN (stateArray_n14) ) ;
    INV_X1 stateArray_U1 ( .A (selSR), .ZN (stateArray_n21) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S00reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2156, stateArray_inS00ser[0]}), .a ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_3126, stateArray_S00reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S00reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2159, stateArray_inS00ser[1]}), .a ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_3127, stateArray_S00reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S00reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2162, stateArray_inS00ser[2]}), .a ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_3128, stateArray_S00reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S00reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2165, stateArray_inS00ser[3]}), .a ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_3129, stateArray_S00reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S00reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2168, stateArray_inS00ser[4]}), .a ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_3130, stateArray_S00reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S00reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2171, stateArray_inS00ser[5]}), .a ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_3131, stateArray_S00reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S00reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2174, stateArray_inS00ser[6]}), .a ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({new_AGEMA_signal_3132, stateArray_S00reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S00reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2177, stateArray_inS00ser[7]}), .a ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({new_AGEMA_signal_3133, stateArray_S00reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S01reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2180, stateArray_inS01ser[0]}), .a ({ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_3134, stateArray_S01reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S01reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2183, stateArray_inS01ser[1]}), .a ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_3135, stateArray_S01reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S01reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2186, stateArray_inS01ser[2]}), .a ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_3136, stateArray_S01reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S01reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2189, stateArray_inS01ser[3]}), .a ({ciphertext_s1[115], ciphertext_s0[115]}), .c ({new_AGEMA_signal_3137, stateArray_S01reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S01reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2192, stateArray_inS01ser[4]}), .a ({ciphertext_s1[116], ciphertext_s0[116]}), .c ({new_AGEMA_signal_3138, stateArray_S01reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S01reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2195, stateArray_inS01ser[5]}), .a ({ciphertext_s1[117], ciphertext_s0[117]}), .c ({new_AGEMA_signal_3139, stateArray_S01reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S01reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2198, stateArray_inS01ser[6]}), .a ({ciphertext_s1[118], ciphertext_s0[118]}), .c ({new_AGEMA_signal_3140, stateArray_S01reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S01reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n20), .b ({new_AGEMA_signal_2201, stateArray_inS01ser[7]}), .a ({ciphertext_s1[119], ciphertext_s0[119]}), .c ({new_AGEMA_signal_3141, stateArray_S01reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S02reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2204, stateArray_inS02ser[0]}), .a ({ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_3142, stateArray_S02reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S02reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2207, stateArray_inS02ser[1]}), .a ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_3143, stateArray_S02reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S02reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2210, stateArray_inS02ser[2]}), .a ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_3144, stateArray_S02reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S02reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2213, stateArray_inS02ser[3]}), .a ({ciphertext_s1[107], ciphertext_s0[107]}), .c ({new_AGEMA_signal_3145, stateArray_S02reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S02reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2216, stateArray_inS02ser[4]}), .a ({ciphertext_s1[108], ciphertext_s0[108]}), .c ({new_AGEMA_signal_3146, stateArray_S02reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S02reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2219, stateArray_inS02ser[5]}), .a ({ciphertext_s1[109], ciphertext_s0[109]}), .c ({new_AGEMA_signal_3147, stateArray_S02reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S02reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2222, stateArray_inS02ser[6]}), .a ({ciphertext_s1[110], ciphertext_s0[110]}), .c ({new_AGEMA_signal_3148, stateArray_S02reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S02reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_2225, stateArray_inS02ser[7]}), .a ({ciphertext_s1[111], ciphertext_s0[111]}), .c ({new_AGEMA_signal_3149, stateArray_S02reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S03reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_3046, stateArray_inS03ser[0]}), .a ({ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_3150, stateArray_S03reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S03reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_3048, stateArray_inS03ser[1]}), .a ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_3151, stateArray_S03reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S03reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_3050, stateArray_inS03ser[2]}), .a ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_3152, stateArray_S03reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S03reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_3052, stateArray_inS03ser[3]}), .a ({ciphertext_s1[99], ciphertext_s0[99]}), .c ({new_AGEMA_signal_3153, stateArray_S03reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S03reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_3054, stateArray_inS03ser[4]}), .a ({ciphertext_s1[100], ciphertext_s0[100]}), .c ({new_AGEMA_signal_3154, stateArray_S03reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S03reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_3056, stateArray_inS03ser[5]}), .a ({ciphertext_s1[101], ciphertext_s0[101]}), .c ({new_AGEMA_signal_3155, stateArray_S03reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S03reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_3058, stateArray_inS03ser[6]}), .a ({ciphertext_s1[102], ciphertext_s0[102]}), .c ({new_AGEMA_signal_3156, stateArray_S03reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S03reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n19), .b ({new_AGEMA_signal_3060, stateArray_inS03ser[7]}), .a ({ciphertext_s1[103], ciphertext_s0[103]}), .c ({new_AGEMA_signal_3157, stateArray_S03reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S10reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2228, stateArray_inS10ser[0]}), .a ({ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_3158, stateArray_S10reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S10reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2231, stateArray_inS10ser[1]}), .a ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_3159, stateArray_S10reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S10reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2234, stateArray_inS10ser[2]}), .a ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_3160, stateArray_S10reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S10reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2237, stateArray_inS10ser[3]}), .a ({ciphertext_s1[83], ciphertext_s0[83]}), .c ({new_AGEMA_signal_3161, stateArray_S10reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S10reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2240, stateArray_inS10ser[4]}), .a ({ciphertext_s1[84], ciphertext_s0[84]}), .c ({new_AGEMA_signal_3162, stateArray_S10reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S10reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2243, stateArray_inS10ser[5]}), .a ({ciphertext_s1[85], ciphertext_s0[85]}), .c ({new_AGEMA_signal_3163, stateArray_S10reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S10reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2246, stateArray_inS10ser[6]}), .a ({ciphertext_s1[86], ciphertext_s0[86]}), .c ({new_AGEMA_signal_3164, stateArray_S10reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S10reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2249, stateArray_inS10ser[7]}), .a ({ciphertext_s1[87], ciphertext_s0[87]}), .c ({new_AGEMA_signal_3165, stateArray_S10reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S11reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2252, stateArray_inS11ser[0]}), .a ({ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_3166, stateArray_S11reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S11reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2255, stateArray_inS11ser[1]}), .a ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_3167, stateArray_S11reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S11reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2258, stateArray_inS11ser[2]}), .a ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_3168, stateArray_S11reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S11reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2261, stateArray_inS11ser[3]}), .a ({ciphertext_s1[75], ciphertext_s0[75]}), .c ({new_AGEMA_signal_3169, stateArray_S11reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S11reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2264, stateArray_inS11ser[4]}), .a ({ciphertext_s1[76], ciphertext_s0[76]}), .c ({new_AGEMA_signal_3170, stateArray_S11reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S11reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2267, stateArray_inS11ser[5]}), .a ({ciphertext_s1[77], ciphertext_s0[77]}), .c ({new_AGEMA_signal_3171, stateArray_S11reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S11reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2270, stateArray_inS11ser[6]}), .a ({ciphertext_s1[78], ciphertext_s0[78]}), .c ({new_AGEMA_signal_3172, stateArray_S11reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S11reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n18), .b ({new_AGEMA_signal_2273, stateArray_inS11ser[7]}), .a ({ciphertext_s1[79], ciphertext_s0[79]}), .c ({new_AGEMA_signal_3173, stateArray_S11reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S12reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2276, stateArray_inS12ser[0]}), .a ({ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_3174, stateArray_S12reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S12reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2279, stateArray_inS12ser[1]}), .a ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_3175, stateArray_S12reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S12reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2282, stateArray_inS12ser[2]}), .a ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_3176, stateArray_S12reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S12reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2285, stateArray_inS12ser[3]}), .a ({ciphertext_s1[67], ciphertext_s0[67]}), .c ({new_AGEMA_signal_3177, stateArray_S12reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S12reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2288, stateArray_inS12ser[4]}), .a ({ciphertext_s1[68], ciphertext_s0[68]}), .c ({new_AGEMA_signal_3178, stateArray_S12reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S12reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2291, stateArray_inS12ser[5]}), .a ({ciphertext_s1[69], ciphertext_s0[69]}), .c ({new_AGEMA_signal_3179, stateArray_S12reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S12reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2294, stateArray_inS12ser[6]}), .a ({ciphertext_s1[70], ciphertext_s0[70]}), .c ({new_AGEMA_signal_3180, stateArray_S12reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S12reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_2297, stateArray_inS12ser[7]}), .a ({ciphertext_s1[71], ciphertext_s0[71]}), .c ({new_AGEMA_signal_3181, stateArray_S12reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S13reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_3062, stateArray_inS13ser[0]}), .a ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_3182, stateArray_S13reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S13reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_3064, stateArray_inS13ser[1]}), .a ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_3183, stateArray_S13reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S13reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_3066, stateArray_inS13ser[2]}), .a ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_3184, stateArray_S13reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S13reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_3068, stateArray_inS13ser[3]}), .a ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_3185, stateArray_S13reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S13reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_3070, stateArray_inS13ser[4]}), .a ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_3186, stateArray_S13reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S13reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_3072, stateArray_inS13ser[5]}), .a ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_3187, stateArray_S13reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S13reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_3074, stateArray_inS13ser[6]}), .a ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({new_AGEMA_signal_3188, stateArray_S13reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S13reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n17), .b ({new_AGEMA_signal_3076, stateArray_inS13ser[7]}), .a ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({new_AGEMA_signal_3189, stateArray_S13reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S20reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2300, stateArray_inS20ser[0]}), .a ({ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_3190, stateArray_S20reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S20reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2303, stateArray_inS20ser[1]}), .a ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_3191, stateArray_S20reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S20reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2306, stateArray_inS20ser[2]}), .a ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_3192, stateArray_S20reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S20reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2309, stateArray_inS20ser[3]}), .a ({ciphertext_s1[43], ciphertext_s0[43]}), .c ({new_AGEMA_signal_3193, stateArray_S20reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S20reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2312, stateArray_inS20ser[4]}), .a ({ciphertext_s1[44], ciphertext_s0[44]}), .c ({new_AGEMA_signal_3194, stateArray_S20reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S20reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2315, stateArray_inS20ser[5]}), .a ({ciphertext_s1[45], ciphertext_s0[45]}), .c ({new_AGEMA_signal_3195, stateArray_S20reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S20reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2318, stateArray_inS20ser[6]}), .a ({ciphertext_s1[46], ciphertext_s0[46]}), .c ({new_AGEMA_signal_3196, stateArray_S20reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S20reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2321, stateArray_inS20ser[7]}), .a ({ciphertext_s1[47], ciphertext_s0[47]}), .c ({new_AGEMA_signal_3197, stateArray_S20reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S21reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2324, stateArray_inS21ser[0]}), .a ({ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_3198, stateArray_S21reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S21reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2327, stateArray_inS21ser[1]}), .a ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_3199, stateArray_S21reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S21reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2330, stateArray_inS21ser[2]}), .a ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_3200, stateArray_S21reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S21reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2333, stateArray_inS21ser[3]}), .a ({ciphertext_s1[35], ciphertext_s0[35]}), .c ({new_AGEMA_signal_3201, stateArray_S21reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S21reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2336, stateArray_inS21ser[4]}), .a ({ciphertext_s1[36], ciphertext_s0[36]}), .c ({new_AGEMA_signal_3202, stateArray_S21reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S21reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2339, stateArray_inS21ser[5]}), .a ({ciphertext_s1[37], ciphertext_s0[37]}), .c ({new_AGEMA_signal_3203, stateArray_S21reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S21reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2342, stateArray_inS21ser[6]}), .a ({ciphertext_s1[38], ciphertext_s0[38]}), .c ({new_AGEMA_signal_3204, stateArray_S21reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S21reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n16), .b ({new_AGEMA_signal_2345, stateArray_inS21ser[7]}), .a ({ciphertext_s1[39], ciphertext_s0[39]}), .c ({new_AGEMA_signal_3205, stateArray_S21reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S22reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_2348, stateArray_inS22ser[0]}), .a ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_3206, stateArray_S22reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S22reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_2351, stateArray_inS22ser[1]}), .a ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_3207, stateArray_S22reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S22reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_2354, stateArray_inS22ser[2]}), .a ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_3208, stateArray_S22reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S22reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_2357, stateArray_inS22ser[3]}), .a ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_3209, stateArray_S22reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S22reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_2360, stateArray_inS22ser[4]}), .a ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_3210, stateArray_S22reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S22reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_2363, stateArray_inS22ser[5]}), .a ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_3211, stateArray_S22reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S22reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_2366, stateArray_inS22ser[6]}), .a ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({new_AGEMA_signal_3212, stateArray_S22reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S22reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_2369, stateArray_inS22ser[7]}), .a ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({new_AGEMA_signal_3213, stateArray_S22reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S23reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3078, stateArray_inS23ser[0]}), .a ({ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_3214, stateArray_S23reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S23reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3080, stateArray_inS23ser[1]}), .a ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_3215, stateArray_S23reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S23reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3082, stateArray_inS23ser[2]}), .a ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_3216, stateArray_S23reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S23reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3084, stateArray_inS23ser[3]}), .a ({ciphertext_s1[51], ciphertext_s0[51]}), .c ({new_AGEMA_signal_3217, stateArray_S23reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S23reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3086, stateArray_inS23ser[4]}), .a ({ciphertext_s1[52], ciphertext_s0[52]}), .c ({new_AGEMA_signal_3218, stateArray_S23reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S23reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3088, stateArray_inS23ser[5]}), .a ({ciphertext_s1[53], ciphertext_s0[53]}), .c ({new_AGEMA_signal_3219, stateArray_S23reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S23reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3090, stateArray_inS23ser[6]}), .a ({ciphertext_s1[54], ciphertext_s0[54]}), .c ({new_AGEMA_signal_3220, stateArray_S23reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S23reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n15), .b ({new_AGEMA_signal_3092, stateArray_inS23ser[7]}), .a ({ciphertext_s1[55], ciphertext_s0[55]}), .c ({new_AGEMA_signal_3221, stateArray_S23reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S30reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2372, stateArray_inS30ser[0]}), .a ({ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_3222, stateArray_S30reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S30reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2375, stateArray_inS30ser[1]}), .a ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_3223, stateArray_S30reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S30reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2378, stateArray_inS30ser[2]}), .a ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_3224, stateArray_S30reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S30reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2381, stateArray_inS30ser[3]}), .a ({ciphertext_s1[3], ciphertext_s0[3]}), .c ({new_AGEMA_signal_3225, stateArray_S30reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S30reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2384, stateArray_inS30ser[4]}), .a ({ciphertext_s1[4], ciphertext_s0[4]}), .c ({new_AGEMA_signal_3226, stateArray_S30reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S30reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2387, stateArray_inS30ser[5]}), .a ({ciphertext_s1[5], ciphertext_s0[5]}), .c ({new_AGEMA_signal_3227, stateArray_S30reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S30reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2390, stateArray_inS30ser[6]}), .a ({ciphertext_s1[6], ciphertext_s0[6]}), .c ({new_AGEMA_signal_3228, stateArray_S30reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S30reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2393, stateArray_inS30ser[7]}), .a ({ciphertext_s1[7], ciphertext_s0[7]}), .c ({new_AGEMA_signal_3229, stateArray_S30reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S31reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2396, stateArray_inS31ser[0]}), .a ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_3230, stateArray_S31reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S31reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2399, stateArray_inS31ser[1]}), .a ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_3231, stateArray_S31reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S31reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2402, stateArray_inS31ser[2]}), .a ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_3232, stateArray_S31reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S31reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2405, stateArray_inS31ser[3]}), .a ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_3233, stateArray_S31reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S31reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2408, stateArray_inS31ser[4]}), .a ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_3234, stateArray_S31reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S31reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2411, stateArray_inS31ser[5]}), .a ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_3235, stateArray_S31reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S31reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2414, stateArray_inS31ser[6]}), .a ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({new_AGEMA_signal_3236, stateArray_S31reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S31reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n14), .b ({new_AGEMA_signal_2417, stateArray_inS31ser[7]}), .a ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({new_AGEMA_signal_3237, stateArray_S31reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S32reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_2420, stateArray_inS32ser[0]}), .a ({ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_3238, stateArray_S32reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S32reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_2423, stateArray_inS32ser[1]}), .a ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_3239, stateArray_S32reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S32reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_2426, stateArray_inS32ser[2]}), .a ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_3240, stateArray_S32reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S32reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_2429, stateArray_inS32ser[3]}), .a ({ciphertext_s1[19], ciphertext_s0[19]}), .c ({new_AGEMA_signal_3241, stateArray_S32reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S32reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_2432, stateArray_inS32ser[4]}), .a ({ciphertext_s1[20], ciphertext_s0[20]}), .c ({new_AGEMA_signal_3242, stateArray_S32reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S32reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_2435, stateArray_inS32ser[5]}), .a ({ciphertext_s1[21], ciphertext_s0[21]}), .c ({new_AGEMA_signal_3243, stateArray_S32reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S32reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_2438, stateArray_inS32ser[6]}), .a ({ciphertext_s1[22], ciphertext_s0[22]}), .c ({new_AGEMA_signal_3244, stateArray_S32reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S32reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_2441, stateArray_inS32ser[7]}), .a ({ciphertext_s1[23], ciphertext_s0[23]}), .c ({new_AGEMA_signal_3245, stateArray_S32reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS00ser_mux_inst_0_U1 ( .s (stateArray_n32), .b ({plaintext_s1[120], plaintext_s0[120]}), .a ({ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_2156, stateArray_inS00ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS00ser_mux_inst_1_U1 ( .s (stateArray_n32), .b ({plaintext_s1[121], plaintext_s0[121]}), .a ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_2159, stateArray_inS00ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS00ser_mux_inst_2_U1 ( .s (stateArray_n32), .b ({plaintext_s1[122], plaintext_s0[122]}), .a ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_2162, stateArray_inS00ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS00ser_mux_inst_3_U1 ( .s (stateArray_n32), .b ({plaintext_s1[123], plaintext_s0[123]}), .a ({ciphertext_s1[115], ciphertext_s0[115]}), .c ({new_AGEMA_signal_2165, stateArray_inS00ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS00ser_mux_inst_4_U1 ( .s (stateArray_n32), .b ({plaintext_s1[124], plaintext_s0[124]}), .a ({ciphertext_s1[116], ciphertext_s0[116]}), .c ({new_AGEMA_signal_2168, stateArray_inS00ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS00ser_mux_inst_5_U1 ( .s (stateArray_n32), .b ({plaintext_s1[125], plaintext_s0[125]}), .a ({ciphertext_s1[117], ciphertext_s0[117]}), .c ({new_AGEMA_signal_2171, stateArray_inS00ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS00ser_mux_inst_6_U1 ( .s (stateArray_n32), .b ({plaintext_s1[126], plaintext_s0[126]}), .a ({ciphertext_s1[118], ciphertext_s0[118]}), .c ({new_AGEMA_signal_2174, stateArray_inS00ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS00ser_mux_inst_7_U1 ( .s (stateArray_n32), .b ({plaintext_s1[127], plaintext_s0[127]}), .a ({ciphertext_s1[119], ciphertext_s0[119]}), .c ({new_AGEMA_signal_2177, stateArray_inS00ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS01ser_mux_inst_0_U1 ( .s (stateArray_n32), .b ({plaintext_s1[112], plaintext_s0[112]}), .a ({ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_2180, stateArray_inS01ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS01ser_mux_inst_1_U1 ( .s (stateArray_n32), .b ({plaintext_s1[113], plaintext_s0[113]}), .a ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_2183, stateArray_inS01ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS01ser_mux_inst_2_U1 ( .s (stateArray_n32), .b ({plaintext_s1[114], plaintext_s0[114]}), .a ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_2186, stateArray_inS01ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS01ser_mux_inst_3_U1 ( .s (stateArray_n32), .b ({plaintext_s1[115], plaintext_s0[115]}), .a ({ciphertext_s1[107], ciphertext_s0[107]}), .c ({new_AGEMA_signal_2189, stateArray_inS01ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS01ser_mux_inst_4_U1 ( .s (stateArray_n32), .b ({plaintext_s1[116], plaintext_s0[116]}), .a ({ciphertext_s1[108], ciphertext_s0[108]}), .c ({new_AGEMA_signal_2192, stateArray_inS01ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS01ser_mux_inst_5_U1 ( .s (stateArray_n32), .b ({plaintext_s1[117], plaintext_s0[117]}), .a ({ciphertext_s1[109], ciphertext_s0[109]}), .c ({new_AGEMA_signal_2195, stateArray_inS01ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS01ser_mux_inst_6_U1 ( .s (stateArray_n32), .b ({plaintext_s1[118], plaintext_s0[118]}), .a ({ciphertext_s1[110], ciphertext_s0[110]}), .c ({new_AGEMA_signal_2198, stateArray_inS01ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS01ser_mux_inst_7_U1 ( .s (stateArray_n32), .b ({plaintext_s1[119], plaintext_s0[119]}), .a ({ciphertext_s1[111], ciphertext_s0[111]}), .c ({new_AGEMA_signal_2201, stateArray_inS01ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS02ser_mux_inst_0_U1 ( .s (stateArray_n31), .b ({plaintext_s1[104], plaintext_s0[104]}), .a ({ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_2204, stateArray_inS02ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS02ser_mux_inst_1_U1 ( .s (stateArray_n31), .b ({plaintext_s1[105], plaintext_s0[105]}), .a ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_2207, stateArray_inS02ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS02ser_mux_inst_2_U1 ( .s (stateArray_n31), .b ({plaintext_s1[106], plaintext_s0[106]}), .a ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_2210, stateArray_inS02ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS02ser_mux_inst_3_U1 ( .s (stateArray_n31), .b ({plaintext_s1[107], plaintext_s0[107]}), .a ({ciphertext_s1[99], ciphertext_s0[99]}), .c ({new_AGEMA_signal_2213, stateArray_inS02ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS02ser_mux_inst_4_U1 ( .s (stateArray_n31), .b ({plaintext_s1[108], plaintext_s0[108]}), .a ({ciphertext_s1[100], ciphertext_s0[100]}), .c ({new_AGEMA_signal_2216, stateArray_inS02ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS02ser_mux_inst_5_U1 ( .s (stateArray_n31), .b ({plaintext_s1[109], plaintext_s0[109]}), .a ({ciphertext_s1[101], ciphertext_s0[101]}), .c ({new_AGEMA_signal_2219, stateArray_inS02ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS02ser_mux_inst_6_U1 ( .s (stateArray_n31), .b ({plaintext_s1[110], plaintext_s0[110]}), .a ({ciphertext_s1[102], ciphertext_s0[102]}), .c ({new_AGEMA_signal_2222, stateArray_inS02ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS02ser_mux_inst_7_U1 ( .s (stateArray_n31), .b ({plaintext_s1[111], plaintext_s0[111]}), .a ({ciphertext_s1[103], ciphertext_s0[103]}), .c ({new_AGEMA_signal_2225, stateArray_inS02ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS10_MC_mux_inst_0_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .a ({new_AGEMA_signal_2880, StateInMC[24]}), .c ({new_AGEMA_signal_3008, stateArray_outS10ser_MC[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS10_MC_mux_inst_1_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .a ({new_AGEMA_signal_2881, StateInMC[25]}), .c ({new_AGEMA_signal_3009, stateArray_outS10ser_MC[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS10_MC_mux_inst_2_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .a ({new_AGEMA_signal_2882, StateInMC[26]}), .c ({new_AGEMA_signal_3010, stateArray_outS10ser_MC[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS10_MC_mux_inst_3_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .a ({new_AGEMA_signal_2883, StateInMC[27]}), .c ({new_AGEMA_signal_3011, stateArray_outS10ser_MC[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS10_MC_mux_inst_4_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .a ({new_AGEMA_signal_2884, StateInMC[28]}), .c ({new_AGEMA_signal_3012, stateArray_outS10ser_MC[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS10_MC_mux_inst_5_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .a ({new_AGEMA_signal_2885, StateInMC[29]}), .c ({new_AGEMA_signal_3013, stateArray_outS10ser_MC[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS10_MC_mux_inst_6_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .a ({new_AGEMA_signal_2886, StateInMC[30]}), .c ({new_AGEMA_signal_3014, stateArray_outS10ser_MC[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS10_MC_mux_inst_7_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .a ({new_AGEMA_signal_2887, StateInMC[31]}), .c ({new_AGEMA_signal_3015, stateArray_outS10ser_MC[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS03ser_mux_inst_0_U1 ( .s (stateArray_n31), .b ({plaintext_s1[96], plaintext_s0[96]}), .a ({new_AGEMA_signal_3008, stateArray_outS10ser_MC[0]}), .c ({new_AGEMA_signal_3046, stateArray_inS03ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS03ser_mux_inst_1_U1 ( .s (stateArray_n31), .b ({plaintext_s1[97], plaintext_s0[97]}), .a ({new_AGEMA_signal_3009, stateArray_outS10ser_MC[1]}), .c ({new_AGEMA_signal_3048, stateArray_inS03ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS03ser_mux_inst_2_U1 ( .s (stateArray_n31), .b ({plaintext_s1[98], plaintext_s0[98]}), .a ({new_AGEMA_signal_3010, stateArray_outS10ser_MC[2]}), .c ({new_AGEMA_signal_3050, stateArray_inS03ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS03ser_mux_inst_3_U1 ( .s (stateArray_n31), .b ({plaintext_s1[99], plaintext_s0[99]}), .a ({new_AGEMA_signal_3011, stateArray_outS10ser_MC[3]}), .c ({new_AGEMA_signal_3052, stateArray_inS03ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS03ser_mux_inst_4_U1 ( .s (stateArray_n31), .b ({plaintext_s1[100], plaintext_s0[100]}), .a ({new_AGEMA_signal_3012, stateArray_outS10ser_MC[4]}), .c ({new_AGEMA_signal_3054, stateArray_inS03ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS03ser_mux_inst_5_U1 ( .s (stateArray_n31), .b ({plaintext_s1[101], plaintext_s0[101]}), .a ({new_AGEMA_signal_3013, stateArray_outS10ser_MC[5]}), .c ({new_AGEMA_signal_3056, stateArray_inS03ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS03ser_mux_inst_6_U1 ( .s (stateArray_n31), .b ({plaintext_s1[102], plaintext_s0[102]}), .a ({new_AGEMA_signal_3014, stateArray_outS10ser_MC[6]}), .c ({new_AGEMA_signal_3058, stateArray_inS03ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS03ser_mux_inst_7_U1 ( .s (stateArray_n31), .b ({plaintext_s1[103], plaintext_s0[103]}), .a ({new_AGEMA_signal_3015, stateArray_outS10ser_MC[7]}), .c ({new_AGEMA_signal_3060, stateArray_inS03ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS10ser_mux_inst_0_U1 ( .s (stateArray_n30), .b ({plaintext_s1[88], plaintext_s0[88]}), .a ({ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_2228, stateArray_inS10ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS10ser_mux_inst_1_U1 ( .s (stateArray_n30), .b ({plaintext_s1[89], plaintext_s0[89]}), .a ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_2231, stateArray_inS10ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS10ser_mux_inst_2_U1 ( .s (stateArray_n30), .b ({plaintext_s1[90], plaintext_s0[90]}), .a ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_2234, stateArray_inS10ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS10ser_mux_inst_3_U1 ( .s (stateArray_n30), .b ({plaintext_s1[91], plaintext_s0[91]}), .a ({ciphertext_s1[83], ciphertext_s0[83]}), .c ({new_AGEMA_signal_2237, stateArray_inS10ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS10ser_mux_inst_4_U1 ( .s (stateArray_n30), .b ({plaintext_s1[92], plaintext_s0[92]}), .a ({ciphertext_s1[84], ciphertext_s0[84]}), .c ({new_AGEMA_signal_2240, stateArray_inS10ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS10ser_mux_inst_5_U1 ( .s (stateArray_n30), .b ({plaintext_s1[93], plaintext_s0[93]}), .a ({ciphertext_s1[85], ciphertext_s0[85]}), .c ({new_AGEMA_signal_2243, stateArray_inS10ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS10ser_mux_inst_6_U1 ( .s (stateArray_n30), .b ({plaintext_s1[94], plaintext_s0[94]}), .a ({ciphertext_s1[86], ciphertext_s0[86]}), .c ({new_AGEMA_signal_2246, stateArray_inS10ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS10ser_mux_inst_7_U1 ( .s (stateArray_n30), .b ({plaintext_s1[95], plaintext_s0[95]}), .a ({ciphertext_s1[87], ciphertext_s0[87]}), .c ({new_AGEMA_signal_2249, stateArray_inS10ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS11ser_mux_inst_0_U1 ( .s (stateArray_n30), .b ({plaintext_s1[80], plaintext_s0[80]}), .a ({ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_2252, stateArray_inS11ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS11ser_mux_inst_1_U1 ( .s (stateArray_n30), .b ({plaintext_s1[81], plaintext_s0[81]}), .a ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_2255, stateArray_inS11ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS11ser_mux_inst_2_U1 ( .s (stateArray_n30), .b ({plaintext_s1[82], plaintext_s0[82]}), .a ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_2258, stateArray_inS11ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS11ser_mux_inst_3_U1 ( .s (stateArray_n30), .b ({plaintext_s1[83], plaintext_s0[83]}), .a ({ciphertext_s1[75], ciphertext_s0[75]}), .c ({new_AGEMA_signal_2261, stateArray_inS11ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS11ser_mux_inst_4_U1 ( .s (stateArray_n30), .b ({plaintext_s1[84], plaintext_s0[84]}), .a ({ciphertext_s1[76], ciphertext_s0[76]}), .c ({new_AGEMA_signal_2264, stateArray_inS11ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS11ser_mux_inst_5_U1 ( .s (stateArray_n30), .b ({plaintext_s1[85], plaintext_s0[85]}), .a ({ciphertext_s1[77], ciphertext_s0[77]}), .c ({new_AGEMA_signal_2267, stateArray_inS11ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS11ser_mux_inst_6_U1 ( .s (stateArray_n30), .b ({plaintext_s1[86], plaintext_s0[86]}), .a ({ciphertext_s1[78], ciphertext_s0[78]}), .c ({new_AGEMA_signal_2270, stateArray_inS11ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS11ser_mux_inst_7_U1 ( .s (stateArray_n30), .b ({plaintext_s1[87], plaintext_s0[87]}), .a ({ciphertext_s1[79], ciphertext_s0[79]}), .c ({new_AGEMA_signal_2273, stateArray_inS11ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS12ser_mux_inst_0_U1 ( .s (stateArray_n29), .b ({plaintext_s1[72], plaintext_s0[72]}), .a ({ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_2276, stateArray_inS12ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS12ser_mux_inst_1_U1 ( .s (stateArray_n29), .b ({plaintext_s1[73], plaintext_s0[73]}), .a ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_2279, stateArray_inS12ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS12ser_mux_inst_2_U1 ( .s (stateArray_n29), .b ({plaintext_s1[74], plaintext_s0[74]}), .a ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_2282, stateArray_inS12ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS12ser_mux_inst_3_U1 ( .s (stateArray_n29), .b ({plaintext_s1[75], plaintext_s0[75]}), .a ({ciphertext_s1[67], ciphertext_s0[67]}), .c ({new_AGEMA_signal_2285, stateArray_inS12ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS12ser_mux_inst_4_U1 ( .s (stateArray_n29), .b ({plaintext_s1[76], plaintext_s0[76]}), .a ({ciphertext_s1[68], ciphertext_s0[68]}), .c ({new_AGEMA_signal_2288, stateArray_inS12ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS12ser_mux_inst_5_U1 ( .s (stateArray_n29), .b ({plaintext_s1[77], plaintext_s0[77]}), .a ({ciphertext_s1[69], ciphertext_s0[69]}), .c ({new_AGEMA_signal_2291, stateArray_inS12ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS12ser_mux_inst_6_U1 ( .s (stateArray_n29), .b ({plaintext_s1[78], plaintext_s0[78]}), .a ({ciphertext_s1[70], ciphertext_s0[70]}), .c ({new_AGEMA_signal_2294, stateArray_inS12ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS12ser_mux_inst_7_U1 ( .s (stateArray_n29), .b ({plaintext_s1[79], plaintext_s0[79]}), .a ({ciphertext_s1[71], ciphertext_s0[71]}), .c ({new_AGEMA_signal_2297, stateArray_inS12ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS20_MC_mux_inst_0_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .a ({new_AGEMA_signal_2872, StateInMC[16]}), .c ({new_AGEMA_signal_3016, stateArray_outS20ser_MC[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS20_MC_mux_inst_1_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .a ({new_AGEMA_signal_2873, StateInMC[17]}), .c ({new_AGEMA_signal_3017, stateArray_outS20ser_MC[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS20_MC_mux_inst_2_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .a ({new_AGEMA_signal_2874, StateInMC[18]}), .c ({new_AGEMA_signal_3018, stateArray_outS20ser_MC[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS20_MC_mux_inst_3_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .a ({new_AGEMA_signal_2875, StateInMC[19]}), .c ({new_AGEMA_signal_3019, stateArray_outS20ser_MC[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS20_MC_mux_inst_4_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .a ({new_AGEMA_signal_2876, StateInMC[20]}), .c ({new_AGEMA_signal_3020, stateArray_outS20ser_MC[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS20_MC_mux_inst_5_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .a ({new_AGEMA_signal_2877, StateInMC[21]}), .c ({new_AGEMA_signal_3021, stateArray_outS20ser_MC[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS20_MC_mux_inst_6_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .a ({new_AGEMA_signal_2878, StateInMC[22]}), .c ({new_AGEMA_signal_3022, stateArray_outS20ser_MC[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS20_MC_mux_inst_7_U1 ( .s (stateArray_n23), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .a ({new_AGEMA_signal_2879, StateInMC[23]}), .c ({new_AGEMA_signal_3023, stateArray_outS20ser_MC[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS13ser_mux_inst_0_U1 ( .s (stateArray_n29), .b ({plaintext_s1[64], plaintext_s0[64]}), .a ({new_AGEMA_signal_3016, stateArray_outS20ser_MC[0]}), .c ({new_AGEMA_signal_3062, stateArray_inS13ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS13ser_mux_inst_1_U1 ( .s (stateArray_n29), .b ({plaintext_s1[65], plaintext_s0[65]}), .a ({new_AGEMA_signal_3017, stateArray_outS20ser_MC[1]}), .c ({new_AGEMA_signal_3064, stateArray_inS13ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS13ser_mux_inst_2_U1 ( .s (stateArray_n29), .b ({plaintext_s1[66], plaintext_s0[66]}), .a ({new_AGEMA_signal_3018, stateArray_outS20ser_MC[2]}), .c ({new_AGEMA_signal_3066, stateArray_inS13ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS13ser_mux_inst_3_U1 ( .s (stateArray_n29), .b ({plaintext_s1[67], plaintext_s0[67]}), .a ({new_AGEMA_signal_3019, stateArray_outS20ser_MC[3]}), .c ({new_AGEMA_signal_3068, stateArray_inS13ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS13ser_mux_inst_4_U1 ( .s (stateArray_n29), .b ({plaintext_s1[68], plaintext_s0[68]}), .a ({new_AGEMA_signal_3020, stateArray_outS20ser_MC[4]}), .c ({new_AGEMA_signal_3070, stateArray_inS13ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS13ser_mux_inst_5_U1 ( .s (stateArray_n29), .b ({plaintext_s1[69], plaintext_s0[69]}), .a ({new_AGEMA_signal_3021, stateArray_outS20ser_MC[5]}), .c ({new_AGEMA_signal_3072, stateArray_inS13ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS13ser_mux_inst_6_U1 ( .s (stateArray_n29), .b ({plaintext_s1[70], plaintext_s0[70]}), .a ({new_AGEMA_signal_3022, stateArray_outS20ser_MC[6]}), .c ({new_AGEMA_signal_3074, stateArray_inS13ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS13ser_mux_inst_7_U1 ( .s (stateArray_n29), .b ({plaintext_s1[71], plaintext_s0[71]}), .a ({new_AGEMA_signal_3023, stateArray_outS20ser_MC[7]}), .c ({new_AGEMA_signal_3076, stateArray_inS13ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS20ser_mux_inst_0_U1 ( .s (stateArray_n28), .b ({plaintext_s1[56], plaintext_s0[56]}), .a ({ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_2300, stateArray_inS20ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS20ser_mux_inst_1_U1 ( .s (stateArray_n28), .b ({plaintext_s1[57], plaintext_s0[57]}), .a ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_2303, stateArray_inS20ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS20ser_mux_inst_2_U1 ( .s (stateArray_n28), .b ({plaintext_s1[58], plaintext_s0[58]}), .a ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_2306, stateArray_inS20ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS20ser_mux_inst_3_U1 ( .s (stateArray_n28), .b ({plaintext_s1[59], plaintext_s0[59]}), .a ({ciphertext_s1[51], ciphertext_s0[51]}), .c ({new_AGEMA_signal_2309, stateArray_inS20ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS20ser_mux_inst_4_U1 ( .s (stateArray_n28), .b ({plaintext_s1[60], plaintext_s0[60]}), .a ({ciphertext_s1[52], ciphertext_s0[52]}), .c ({new_AGEMA_signal_2312, stateArray_inS20ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS20ser_mux_inst_5_U1 ( .s (stateArray_n28), .b ({plaintext_s1[61], plaintext_s0[61]}), .a ({ciphertext_s1[53], ciphertext_s0[53]}), .c ({new_AGEMA_signal_2315, stateArray_inS20ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS20ser_mux_inst_6_U1 ( .s (stateArray_n28), .b ({plaintext_s1[62], plaintext_s0[62]}), .a ({ciphertext_s1[54], ciphertext_s0[54]}), .c ({new_AGEMA_signal_2318, stateArray_inS20ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS20ser_mux_inst_7_U1 ( .s (stateArray_n28), .b ({plaintext_s1[63], plaintext_s0[63]}), .a ({ciphertext_s1[55], ciphertext_s0[55]}), .c ({new_AGEMA_signal_2321, stateArray_inS20ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS21ser_mux_inst_0_U1 ( .s (stateArray_n28), .b ({plaintext_s1[48], plaintext_s0[48]}), .a ({ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_2324, stateArray_inS21ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS21ser_mux_inst_1_U1 ( .s (stateArray_n28), .b ({plaintext_s1[49], plaintext_s0[49]}), .a ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_2327, stateArray_inS21ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS21ser_mux_inst_2_U1 ( .s (stateArray_n28), .b ({plaintext_s1[50], plaintext_s0[50]}), .a ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_2330, stateArray_inS21ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS21ser_mux_inst_3_U1 ( .s (stateArray_n28), .b ({plaintext_s1[51], plaintext_s0[51]}), .a ({ciphertext_s1[43], ciphertext_s0[43]}), .c ({new_AGEMA_signal_2333, stateArray_inS21ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS21ser_mux_inst_4_U1 ( .s (stateArray_n28), .b ({plaintext_s1[52], plaintext_s0[52]}), .a ({ciphertext_s1[44], ciphertext_s0[44]}), .c ({new_AGEMA_signal_2336, stateArray_inS21ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS21ser_mux_inst_5_U1 ( .s (stateArray_n28), .b ({plaintext_s1[53], plaintext_s0[53]}), .a ({ciphertext_s1[45], ciphertext_s0[45]}), .c ({new_AGEMA_signal_2339, stateArray_inS21ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS21ser_mux_inst_6_U1 ( .s (stateArray_n28), .b ({plaintext_s1[54], plaintext_s0[54]}), .a ({ciphertext_s1[46], ciphertext_s0[46]}), .c ({new_AGEMA_signal_2342, stateArray_inS21ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS21ser_mux_inst_7_U1 ( .s (stateArray_n28), .b ({plaintext_s1[55], plaintext_s0[55]}), .a ({ciphertext_s1[47], ciphertext_s0[47]}), .c ({new_AGEMA_signal_2345, stateArray_inS21ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS22ser_mux_inst_0_U1 ( .s (stateArray_n27), .b ({plaintext_s1[40], plaintext_s0[40]}), .a ({ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_2348, stateArray_inS22ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS22ser_mux_inst_1_U1 ( .s (stateArray_n27), .b ({plaintext_s1[41], plaintext_s0[41]}), .a ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_2351, stateArray_inS22ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS22ser_mux_inst_2_U1 ( .s (stateArray_n27), .b ({plaintext_s1[42], plaintext_s0[42]}), .a ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_2354, stateArray_inS22ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS22ser_mux_inst_3_U1 ( .s (stateArray_n27), .b ({plaintext_s1[43], plaintext_s0[43]}), .a ({ciphertext_s1[35], ciphertext_s0[35]}), .c ({new_AGEMA_signal_2357, stateArray_inS22ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS22ser_mux_inst_4_U1 ( .s (stateArray_n27), .b ({plaintext_s1[44], plaintext_s0[44]}), .a ({ciphertext_s1[36], ciphertext_s0[36]}), .c ({new_AGEMA_signal_2360, stateArray_inS22ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS22ser_mux_inst_5_U1 ( .s (stateArray_n27), .b ({plaintext_s1[45], plaintext_s0[45]}), .a ({ciphertext_s1[37], ciphertext_s0[37]}), .c ({new_AGEMA_signal_2363, stateArray_inS22ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS22ser_mux_inst_6_U1 ( .s (stateArray_n27), .b ({plaintext_s1[46], plaintext_s0[46]}), .a ({ciphertext_s1[38], ciphertext_s0[38]}), .c ({new_AGEMA_signal_2366, stateArray_inS22ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS22ser_mux_inst_7_U1 ( .s (stateArray_n27), .b ({plaintext_s1[47], plaintext_s0[47]}), .a ({ciphertext_s1[39], ciphertext_s0[39]}), .c ({new_AGEMA_signal_2369, stateArray_inS22ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS30_MC_mux_inst_0_U1 ( .s (stateArray_n22), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .a ({new_AGEMA_signal_2864, StateInMC[8]}), .c ({new_AGEMA_signal_3024, stateArray_outS30ser_MC[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS30_MC_mux_inst_1_U1 ( .s (stateArray_n22), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .a ({new_AGEMA_signal_2865, StateInMC[9]}), .c ({new_AGEMA_signal_3025, stateArray_outS30ser_MC[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS30_MC_mux_inst_2_U1 ( .s (stateArray_n22), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .a ({new_AGEMA_signal_2866, StateInMC[10]}), .c ({new_AGEMA_signal_3026, stateArray_outS30ser_MC[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS30_MC_mux_inst_3_U1 ( .s (stateArray_n22), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .a ({new_AGEMA_signal_2867, StateInMC[11]}), .c ({new_AGEMA_signal_3027, stateArray_outS30ser_MC[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS30_MC_mux_inst_4_U1 ( .s (stateArray_n22), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .a ({new_AGEMA_signal_2868, StateInMC[12]}), .c ({new_AGEMA_signal_3028, stateArray_outS30ser_MC[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS30_MC_mux_inst_5_U1 ( .s (stateArray_n22), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .a ({new_AGEMA_signal_2869, StateInMC[13]}), .c ({new_AGEMA_signal_3029, stateArray_outS30ser_MC[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS30_MC_mux_inst_6_U1 ( .s (stateArray_n22), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .a ({new_AGEMA_signal_2870, StateInMC[14]}), .c ({new_AGEMA_signal_3030, stateArray_outS30ser_MC[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_outS30_MC_mux_inst_7_U1 ( .s (stateArray_n22), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .a ({new_AGEMA_signal_2871, StateInMC[15]}), .c ({new_AGEMA_signal_3031, stateArray_outS30ser_MC[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS23ser_mux_inst_0_U1 ( .s (stateArray_n27), .b ({plaintext_s1[32], plaintext_s0[32]}), .a ({new_AGEMA_signal_3024, stateArray_outS30ser_MC[0]}), .c ({new_AGEMA_signal_3078, stateArray_inS23ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS23ser_mux_inst_1_U1 ( .s (stateArray_n27), .b ({plaintext_s1[33], plaintext_s0[33]}), .a ({new_AGEMA_signal_3025, stateArray_outS30ser_MC[1]}), .c ({new_AGEMA_signal_3080, stateArray_inS23ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS23ser_mux_inst_2_U1 ( .s (stateArray_n27), .b ({plaintext_s1[34], plaintext_s0[34]}), .a ({new_AGEMA_signal_3026, stateArray_outS30ser_MC[2]}), .c ({new_AGEMA_signal_3082, stateArray_inS23ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS23ser_mux_inst_3_U1 ( .s (stateArray_n27), .b ({plaintext_s1[35], plaintext_s0[35]}), .a ({new_AGEMA_signal_3027, stateArray_outS30ser_MC[3]}), .c ({new_AGEMA_signal_3084, stateArray_inS23ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS23ser_mux_inst_4_U1 ( .s (stateArray_n27), .b ({plaintext_s1[36], plaintext_s0[36]}), .a ({new_AGEMA_signal_3028, stateArray_outS30ser_MC[4]}), .c ({new_AGEMA_signal_3086, stateArray_inS23ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS23ser_mux_inst_5_U1 ( .s (stateArray_n27), .b ({plaintext_s1[37], plaintext_s0[37]}), .a ({new_AGEMA_signal_3029, stateArray_outS30ser_MC[5]}), .c ({new_AGEMA_signal_3088, stateArray_inS23ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS23ser_mux_inst_6_U1 ( .s (stateArray_n27), .b ({plaintext_s1[38], plaintext_s0[38]}), .a ({new_AGEMA_signal_3030, stateArray_outS30ser_MC[6]}), .c ({new_AGEMA_signal_3090, stateArray_inS23ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS23ser_mux_inst_7_U1 ( .s (stateArray_n27), .b ({plaintext_s1[39], plaintext_s0[39]}), .a ({new_AGEMA_signal_3031, stateArray_outS30ser_MC[7]}), .c ({new_AGEMA_signal_3092, stateArray_inS23ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS30ser_mux_inst_0_U1 ( .s (stateArray_n26), .b ({plaintext_s1[24], plaintext_s0[24]}), .a ({ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_2372, stateArray_inS30ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS30ser_mux_inst_1_U1 ( .s (stateArray_n26), .b ({plaintext_s1[25], plaintext_s0[25]}), .a ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_2375, stateArray_inS30ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS30ser_mux_inst_2_U1 ( .s (stateArray_n26), .b ({plaintext_s1[26], plaintext_s0[26]}), .a ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_2378, stateArray_inS30ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS30ser_mux_inst_3_U1 ( .s (stateArray_n26), .b ({plaintext_s1[27], plaintext_s0[27]}), .a ({ciphertext_s1[19], ciphertext_s0[19]}), .c ({new_AGEMA_signal_2381, stateArray_inS30ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS30ser_mux_inst_4_U1 ( .s (stateArray_n26), .b ({plaintext_s1[28], plaintext_s0[28]}), .a ({ciphertext_s1[20], ciphertext_s0[20]}), .c ({new_AGEMA_signal_2384, stateArray_inS30ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS30ser_mux_inst_5_U1 ( .s (stateArray_n26), .b ({plaintext_s1[29], plaintext_s0[29]}), .a ({ciphertext_s1[21], ciphertext_s0[21]}), .c ({new_AGEMA_signal_2387, stateArray_inS30ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS30ser_mux_inst_6_U1 ( .s (stateArray_n26), .b ({plaintext_s1[30], plaintext_s0[30]}), .a ({ciphertext_s1[22], ciphertext_s0[22]}), .c ({new_AGEMA_signal_2390, stateArray_inS30ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS30ser_mux_inst_7_U1 ( .s (stateArray_n26), .b ({plaintext_s1[31], plaintext_s0[31]}), .a ({ciphertext_s1[23], ciphertext_s0[23]}), .c ({new_AGEMA_signal_2393, stateArray_inS30ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS31ser_mux_inst_0_U1 ( .s (stateArray_n26), .b ({plaintext_s1[16], plaintext_s0[16]}), .a ({ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_2396, stateArray_inS31ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS31ser_mux_inst_1_U1 ( .s (stateArray_n26), .b ({plaintext_s1[17], plaintext_s0[17]}), .a ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_2399, stateArray_inS31ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS31ser_mux_inst_2_U1 ( .s (stateArray_n26), .b ({plaintext_s1[18], plaintext_s0[18]}), .a ({ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_2402, stateArray_inS31ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS31ser_mux_inst_3_U1 ( .s (stateArray_n26), .b ({plaintext_s1[19], plaintext_s0[19]}), .a ({ciphertext_s1[11], ciphertext_s0[11]}), .c ({new_AGEMA_signal_2405, stateArray_inS31ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS31ser_mux_inst_4_U1 ( .s (stateArray_n26), .b ({plaintext_s1[20], plaintext_s0[20]}), .a ({ciphertext_s1[12], ciphertext_s0[12]}), .c ({new_AGEMA_signal_2408, stateArray_inS31ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS31ser_mux_inst_5_U1 ( .s (stateArray_n26), .b ({plaintext_s1[21], plaintext_s0[21]}), .a ({ciphertext_s1[13], ciphertext_s0[13]}), .c ({new_AGEMA_signal_2411, stateArray_inS31ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS31ser_mux_inst_6_U1 ( .s (stateArray_n26), .b ({plaintext_s1[22], plaintext_s0[22]}), .a ({ciphertext_s1[14], ciphertext_s0[14]}), .c ({new_AGEMA_signal_2414, stateArray_inS31ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS31ser_mux_inst_7_U1 ( .s (stateArray_n26), .b ({plaintext_s1[23], plaintext_s0[23]}), .a ({ciphertext_s1[15], ciphertext_s0[15]}), .c ({new_AGEMA_signal_2417, stateArray_inS31ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS32ser_mux_inst_0_U1 ( .s (stateArray_n25), .b ({plaintext_s1[8], plaintext_s0[8]}), .a ({ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_2420, stateArray_inS32ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS32ser_mux_inst_1_U1 ( .s (stateArray_n25), .b ({plaintext_s1[9], plaintext_s0[9]}), .a ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_2423, stateArray_inS32ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS32ser_mux_inst_2_U1 ( .s (stateArray_n25), .b ({plaintext_s1[10], plaintext_s0[10]}), .a ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_2426, stateArray_inS32ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS32ser_mux_inst_3_U1 ( .s (stateArray_n25), .b ({plaintext_s1[11], plaintext_s0[11]}), .a ({ciphertext_s1[3], ciphertext_s0[3]}), .c ({new_AGEMA_signal_2429, stateArray_inS32ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS32ser_mux_inst_4_U1 ( .s (stateArray_n25), .b ({plaintext_s1[12], plaintext_s0[12]}), .a ({ciphertext_s1[4], ciphertext_s0[4]}), .c ({new_AGEMA_signal_2432, stateArray_inS32ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS32ser_mux_inst_5_U1 ( .s (stateArray_n25), .b ({plaintext_s1[13], plaintext_s0[13]}), .a ({ciphertext_s1[5], ciphertext_s0[5]}), .c ({new_AGEMA_signal_2435, stateArray_inS32ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS32ser_mux_inst_6_U1 ( .s (stateArray_n25), .b ({plaintext_s1[14], plaintext_s0[14]}), .a ({ciphertext_s1[6], ciphertext_s0[6]}), .c ({new_AGEMA_signal_2438, stateArray_inS32ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS32ser_mux_inst_7_U1 ( .s (stateArray_n25), .b ({plaintext_s1[15], plaintext_s0[15]}), .a ({ciphertext_s1[7], ciphertext_s0[7]}), .c ({new_AGEMA_signal_2441, stateArray_inS32ser[7]}) ) ;
    INV_X1 MUX_StateInMC_U3 ( .A (intFinal), .ZN (MUX_StateInMC_n7) ) ;
    INV_X1 MUX_StateInMC_U2 ( .A (MUX_StateInMC_n7), .ZN (MUX_StateInMC_n6) ) ;
    INV_X1 MUX_StateInMC_U1 ( .A (MUX_StateInMC_n7), .ZN (MUX_StateInMC_n5) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_0_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2825, MCout[0]}), .a ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_2860, StateInMC[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_1_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2849, MCout[1]}), .a ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_2861, StateInMC[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_2_U1 ( .s (intFinal), .b ({new_AGEMA_signal_2823, MCout[2]}), .a ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_2834, StateInMC[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_3_U1 ( .s (intFinal), .b ({new_AGEMA_signal_2848, MCout[3]}), .a ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_2862, StateInMC[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_4_U1 ( .s (intFinal), .b ({new_AGEMA_signal_2847, MCout[4]}), .a ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_2863, StateInMC[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_5_U1 ( .s (intFinal), .b ({new_AGEMA_signal_2820, MCout[5]}), .a ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_2835, StateInMC[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_6_U1 ( .s (intFinal), .b ({new_AGEMA_signal_2819, MCout[6]}), .a ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({new_AGEMA_signal_2836, StateInMC[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_7_U1 ( .s (intFinal), .b ({new_AGEMA_signal_2818, MCout[7]}), .a ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({new_AGEMA_signal_2837, StateInMC[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_8_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2817, MCout[8]}), .a ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_2864, StateInMC[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_9_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2846, MCout[9]}), .a ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_2865, StateInMC[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_10_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2815, MCout[10]}), .a ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_2866, StateInMC[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_11_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2845, MCout[11]}), .a ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_2867, StateInMC[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_12_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2844, MCout[12]}), .a ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_2868, StateInMC[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_13_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2812, MCout[13]}), .a ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_2869, StateInMC[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_14_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2811, MCout[14]}), .a ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({new_AGEMA_signal_2870, StateInMC[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_15_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2810, MCout[15]}), .a ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({new_AGEMA_signal_2871, StateInMC[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_16_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2809, MCout[16]}), .a ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_2872, StateInMC[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_17_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2843, MCout[17]}), .a ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_2873, StateInMC[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_18_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2807, MCout[18]}), .a ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_2874, StateInMC[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_19_U1 ( .s (MUX_StateInMC_n6), .b ({new_AGEMA_signal_2842, MCout[19]}), .a ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_2875, StateInMC[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_20_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2841, MCout[20]}), .a ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_2876, StateInMC[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_21_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2804, MCout[21]}), .a ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_2877, StateInMC[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_22_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2803, MCout[22]}), .a ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({new_AGEMA_signal_2878, StateInMC[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_23_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2802, MCout[23]}), .a ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({new_AGEMA_signal_2879, StateInMC[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_24_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2801, MCout[24]}), .a ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_2880, StateInMC[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_25_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2840, MCout[25]}), .a ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_2881, StateInMC[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_26_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2799, MCout[26]}), .a ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_2882, StateInMC[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_27_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2839, MCout[27]}), .a ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_2883, StateInMC[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_28_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2838, MCout[28]}), .a ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_2884, StateInMC[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_29_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2796, MCout[29]}), .a ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_2885, StateInMC[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_30_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2795, MCout[30]}), .a ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({new_AGEMA_signal_2886, StateInMC[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateInMC_mux_inst_31_U1 ( .s (MUX_StateInMC_n5), .b ({new_AGEMA_signal_2794, MCout[31]}), .a ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({new_AGEMA_signal_2887, StateInMC[31]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U50 ( .a ({new_AGEMA_signal_2006, KeyArray_outS01ser_7_}), .b ({new_AGEMA_signal_2004, keyStateIn[7]}), .c ({new_AGEMA_signal_2007, KeyArray_outS01ser_XOR_00[7]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U49 ( .a ({new_AGEMA_signal_2008, KeyArray_outS01ser_6_}), .b ({new_AGEMA_signal_2001, keyStateIn[6]}), .c ({new_AGEMA_signal_2009, KeyArray_outS01ser_XOR_00[6]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U48 ( .a ({new_AGEMA_signal_2010, KeyArray_outS01ser_5_}), .b ({new_AGEMA_signal_1998, keyStateIn[5]}), .c ({new_AGEMA_signal_2011, KeyArray_outS01ser_XOR_00[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U47 ( .a ({new_AGEMA_signal_2012, KeyArray_outS01ser_4_}), .b ({new_AGEMA_signal_1995, keyStateIn[4]}), .c ({new_AGEMA_signal_2013, KeyArray_outS01ser_XOR_00[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U46 ( .a ({new_AGEMA_signal_2014, KeyArray_outS01ser_3_}), .b ({new_AGEMA_signal_1992, keyStateIn[3]}), .c ({new_AGEMA_signal_2015, KeyArray_outS01ser_XOR_00[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U45 ( .a ({new_AGEMA_signal_2016, KeyArray_outS01ser_2_}), .b ({new_AGEMA_signal_1989, keyStateIn[2]}), .c ({new_AGEMA_signal_2017, KeyArray_outS01ser_XOR_00[2]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U44 ( .a ({new_AGEMA_signal_2018, KeyArray_outS01ser_1_}), .b ({new_AGEMA_signal_1986, keyStateIn[1]}), .c ({new_AGEMA_signal_2019, KeyArray_outS01ser_XOR_00[1]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U43 ( .a ({new_AGEMA_signal_2020, KeyArray_outS01ser_0_}), .b ({new_AGEMA_signal_1983, keyStateIn[0]}), .c ({new_AGEMA_signal_2021, KeyArray_outS01ser_XOR_00[0]}) ) ;
    INV_X1 KeyArray_U26 ( .A (KeyArray_n47), .ZN (KeyArray_n46) ) ;
    INV_X1 KeyArray_U25 ( .A (KeyArray_n47), .ZN (KeyArray_n45) ) ;
    INV_X1 KeyArray_U24 ( .A (KeyArray_n47), .ZN (KeyArray_n44) ) ;
    INV_X1 KeyArray_U23 ( .A (KeyArray_n47), .ZN (KeyArray_n43) ) ;
    INV_X1 KeyArray_U22 ( .A (KeyArray_n47), .ZN (KeyArray_n42) ) ;
    INV_X1 KeyArray_U21 ( .A (KeyArray_n47), .ZN (KeyArray_n41) ) ;
    INV_X1 KeyArray_U20 ( .A (KeyArray_n47), .ZN (KeyArray_n40) ) ;
    INV_X1 KeyArray_U19 ( .A (KeyArray_n47), .ZN (KeyArray_n39) ) ;
    INV_X1 KeyArray_U18 ( .A (nReset), .ZN (KeyArray_n47) ) ;
    INV_X1 KeyArray_U17 ( .A (KeyArray_n38), .ZN (KeyArray_n31) ) ;
    INV_X1 KeyArray_U16 ( .A (KeyArray_n29), .ZN (KeyArray_n23) ) ;
    INV_X1 KeyArray_U15 ( .A (KeyArray_n38), .ZN (KeyArray_n37) ) ;
    INV_X1 KeyArray_U14 ( .A (KeyArray_n29), .ZN (KeyArray_n28) ) ;
    INV_X1 KeyArray_U13 ( .A (KeyArray_n38), .ZN (KeyArray_n36) ) ;
    INV_X1 KeyArray_U12 ( .A (KeyArray_n29), .ZN (KeyArray_n27) ) ;
    INV_X1 KeyArray_U11 ( .A (KeyArray_n38), .ZN (KeyArray_n35) ) ;
    INV_X1 KeyArray_U10 ( .A (KeyArray_n29), .ZN (KeyArray_n26) ) ;
    INV_X1 KeyArray_U9 ( .A (KeyArray_n38), .ZN (KeyArray_n32) ) ;
    INV_X1 KeyArray_U8 ( .A (KeyArray_n29), .ZN (KeyArray_n24) ) ;
    INV_X1 KeyArray_U7 ( .A (KeyArray_n38), .ZN (KeyArray_n33) ) ;
    INV_X1 KeyArray_U6 ( .A (KeyArray_n29), .ZN (KeyArray_n25) ) ;
    INV_X1 KeyArray_U5 ( .A (KeyArray_n38), .ZN (KeyArray_n30) ) ;
    INV_X1 KeyArray_U4 ( .A (KeyArray_n29), .ZN (KeyArray_n22) ) ;
    INV_X1 KeyArray_U3 ( .A (KeyArray_n38), .ZN (KeyArray_n34) ) ;
    INV_X1 KeyArray_U2 ( .A (selMC), .ZN (KeyArray_n38) ) ;
    INV_X1 KeyArray_U1 ( .A (n12), .ZN (KeyArray_n29) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_0_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_1983, keyStateIn[0]}), .a ({new_AGEMA_signal_3267, KeyArray_S00reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3375, KeyArray_S00reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3247, KeyArray_inS00ser[0]}), .a ({new_AGEMA_signal_2491, KeyArray_outS10ser[0]}), .c ({new_AGEMA_signal_3267, KeyArray_S00reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_1_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_1986, keyStateIn[1]}), .a ({new_AGEMA_signal_3268, KeyArray_S00reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3376, KeyArray_S00reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3249, KeyArray_inS00ser[1]}), .a ({new_AGEMA_signal_2494, KeyArray_outS10ser[1]}), .c ({new_AGEMA_signal_3268, KeyArray_S00reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_2_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_1989, keyStateIn[2]}), .a ({new_AGEMA_signal_3269, KeyArray_S00reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3377, KeyArray_S00reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3251, KeyArray_inS00ser[2]}), .a ({new_AGEMA_signal_2497, KeyArray_outS10ser[2]}), .c ({new_AGEMA_signal_3269, KeyArray_S00reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_3_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_1992, keyStateIn[3]}), .a ({new_AGEMA_signal_3270, KeyArray_S00reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3378, KeyArray_S00reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3253, KeyArray_inS00ser[3]}), .a ({new_AGEMA_signal_2500, KeyArray_outS10ser[3]}), .c ({new_AGEMA_signal_3270, KeyArray_S00reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_4_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_1995, keyStateIn[4]}), .a ({new_AGEMA_signal_3271, KeyArray_S00reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3379, KeyArray_S00reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3255, KeyArray_inS00ser[4]}), .a ({new_AGEMA_signal_2503, KeyArray_outS10ser[4]}), .c ({new_AGEMA_signal_3271, KeyArray_S00reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_5_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_1998, keyStateIn[5]}), .a ({new_AGEMA_signal_3272, KeyArray_S00reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3380, KeyArray_S00reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3257, KeyArray_inS00ser[5]}), .a ({new_AGEMA_signal_2506, KeyArray_outS10ser[5]}), .c ({new_AGEMA_signal_3272, KeyArray_S00reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_6_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2001, keyStateIn[6]}), .a ({new_AGEMA_signal_3273, KeyArray_S00reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3381, KeyArray_S00reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3259, KeyArray_inS00ser[6]}), .a ({new_AGEMA_signal_2509, KeyArray_outS10ser[6]}), .c ({new_AGEMA_signal_3273, KeyArray_S00reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_7_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2004, keyStateIn[7]}), .a ({new_AGEMA_signal_3274, KeyArray_S00reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3382, KeyArray_S00reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_3261, KeyArray_inS00ser[7]}), .a ({new_AGEMA_signal_2512, KeyArray_outS10ser[7]}), .c ({new_AGEMA_signal_3274, KeyArray_S00reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_0_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2020, KeyArray_outS01ser_0_}), .a ({new_AGEMA_signal_2888, KeyArray_S01reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3275, KeyArray_S01reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_2444, KeyArray_inS01ser[0]}), .a ({new_AGEMA_signal_2515, KeyArray_outS11ser[0]}), .c ({new_AGEMA_signal_2888, KeyArray_S01reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_1_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2018, KeyArray_outS01ser_1_}), .a ({new_AGEMA_signal_2889, KeyArray_S01reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3276, KeyArray_S01reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_2447, KeyArray_inS01ser[1]}), .a ({new_AGEMA_signal_2518, KeyArray_outS11ser[1]}), .c ({new_AGEMA_signal_2889, KeyArray_S01reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_2_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2016, KeyArray_outS01ser_2_}), .a ({new_AGEMA_signal_2890, KeyArray_S01reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3277, KeyArray_S01reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_2450, KeyArray_inS01ser[2]}), .a ({new_AGEMA_signal_2521, KeyArray_outS11ser[2]}), .c ({new_AGEMA_signal_2890, KeyArray_S01reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_3_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2014, KeyArray_outS01ser_3_}), .a ({new_AGEMA_signal_2891, KeyArray_S01reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3278, KeyArray_S01reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_2453, KeyArray_inS01ser[3]}), .a ({new_AGEMA_signal_2524, KeyArray_outS11ser[3]}), .c ({new_AGEMA_signal_2891, KeyArray_S01reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_4_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2012, KeyArray_outS01ser_4_}), .a ({new_AGEMA_signal_2892, KeyArray_S01reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3279, KeyArray_S01reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_2456, KeyArray_inS01ser[4]}), .a ({new_AGEMA_signal_2527, KeyArray_outS11ser[4]}), .c ({new_AGEMA_signal_2892, KeyArray_S01reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_5_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2010, KeyArray_outS01ser_5_}), .a ({new_AGEMA_signal_2893, KeyArray_S01reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3280, KeyArray_S01reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_2459, KeyArray_inS01ser[5]}), .a ({new_AGEMA_signal_2530, KeyArray_outS11ser[5]}), .c ({new_AGEMA_signal_2893, KeyArray_S01reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_6_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2008, KeyArray_outS01ser_6_}), .a ({new_AGEMA_signal_2894, KeyArray_S01reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3281, KeyArray_S01reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_2462, KeyArray_inS01ser[6]}), .a ({new_AGEMA_signal_2533, KeyArray_outS11ser[6]}), .c ({new_AGEMA_signal_2894, KeyArray_S01reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_7_U1 ( .s (KeyArray_n28), .b ({new_AGEMA_signal_2006, KeyArray_outS01ser_7_}), .a ({new_AGEMA_signal_2895, KeyArray_S01reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3282, KeyArray_S01reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n37), .b ({new_AGEMA_signal_2465, KeyArray_inS01ser[7]}), .a ({new_AGEMA_signal_2536, KeyArray_outS11ser[7]}), .c ({new_AGEMA_signal_2895, KeyArray_S01reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_0_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2443, KeyArray_outS02ser[0]}), .a ({new_AGEMA_signal_2896, KeyArray_S02reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3283, KeyArray_S02reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2468, KeyArray_inS02ser[0]}), .a ({new_AGEMA_signal_2539, KeyArray_outS12ser[0]}), .c ({new_AGEMA_signal_2896, KeyArray_S02reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_1_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2446, KeyArray_outS02ser[1]}), .a ({new_AGEMA_signal_2897, KeyArray_S02reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3284, KeyArray_S02reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2471, KeyArray_inS02ser[1]}), .a ({new_AGEMA_signal_2542, KeyArray_outS12ser[1]}), .c ({new_AGEMA_signal_2897, KeyArray_S02reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_2_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2449, KeyArray_outS02ser[2]}), .a ({new_AGEMA_signal_2898, KeyArray_S02reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3285, KeyArray_S02reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2474, KeyArray_inS02ser[2]}), .a ({new_AGEMA_signal_2545, KeyArray_outS12ser[2]}), .c ({new_AGEMA_signal_2898, KeyArray_S02reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_3_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2452, KeyArray_outS02ser[3]}), .a ({new_AGEMA_signal_2899, KeyArray_S02reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3286, KeyArray_S02reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2477, KeyArray_inS02ser[3]}), .a ({new_AGEMA_signal_2548, KeyArray_outS12ser[3]}), .c ({new_AGEMA_signal_2899, KeyArray_S02reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_4_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2455, KeyArray_outS02ser[4]}), .a ({new_AGEMA_signal_2900, KeyArray_S02reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3287, KeyArray_S02reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2480, KeyArray_inS02ser[4]}), .a ({new_AGEMA_signal_2551, KeyArray_outS12ser[4]}), .c ({new_AGEMA_signal_2900, KeyArray_S02reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_5_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2458, KeyArray_outS02ser[5]}), .a ({new_AGEMA_signal_2901, KeyArray_S02reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3288, KeyArray_S02reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2483, KeyArray_inS02ser[5]}), .a ({new_AGEMA_signal_2554, KeyArray_outS12ser[5]}), .c ({new_AGEMA_signal_2901, KeyArray_S02reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_6_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2461, KeyArray_outS02ser[6]}), .a ({new_AGEMA_signal_2902, KeyArray_S02reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3289, KeyArray_S02reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2486, KeyArray_inS02ser[6]}), .a ({new_AGEMA_signal_2557, KeyArray_outS12ser[6]}), .c ({new_AGEMA_signal_2902, KeyArray_S02reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_7_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2464, KeyArray_outS02ser[7]}), .a ({new_AGEMA_signal_2903, KeyArray_S02reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3290, KeyArray_S02reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2489, KeyArray_inS02ser[7]}), .a ({new_AGEMA_signal_2560, KeyArray_outS12ser[7]}), .c ({new_AGEMA_signal_2903, KeyArray_S02reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_0_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2467, KeyArray_outS03ser[0]}), .a ({new_AGEMA_signal_2904, KeyArray_S03reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3291, KeyArray_S03reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2492, KeyArray_inS03ser[0]}), .a ({new_AGEMA_signal_2563, keySBIn[0]}), .c ({new_AGEMA_signal_2904, KeyArray_S03reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_1_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2470, KeyArray_outS03ser[1]}), .a ({new_AGEMA_signal_2905, KeyArray_S03reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3292, KeyArray_S03reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2495, KeyArray_inS03ser[1]}), .a ({new_AGEMA_signal_2566, keySBIn[1]}), .c ({new_AGEMA_signal_2905, KeyArray_S03reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_2_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2473, KeyArray_outS03ser[2]}), .a ({new_AGEMA_signal_2906, KeyArray_S03reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3293, KeyArray_S03reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2498, KeyArray_inS03ser[2]}), .a ({new_AGEMA_signal_2569, keySBIn[2]}), .c ({new_AGEMA_signal_2906, KeyArray_S03reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_3_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2476, KeyArray_outS03ser[3]}), .a ({new_AGEMA_signal_2907, KeyArray_S03reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3294, KeyArray_S03reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2501, KeyArray_inS03ser[3]}), .a ({new_AGEMA_signal_2572, keySBIn[3]}), .c ({new_AGEMA_signal_2907, KeyArray_S03reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_4_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2479, KeyArray_outS03ser[4]}), .a ({new_AGEMA_signal_2908, KeyArray_S03reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3295, KeyArray_S03reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2504, KeyArray_inS03ser[4]}), .a ({new_AGEMA_signal_2575, keySBIn[4]}), .c ({new_AGEMA_signal_2908, KeyArray_S03reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_5_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2482, KeyArray_outS03ser[5]}), .a ({new_AGEMA_signal_2909, KeyArray_S03reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3296, KeyArray_S03reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2507, KeyArray_inS03ser[5]}), .a ({new_AGEMA_signal_2578, keySBIn[5]}), .c ({new_AGEMA_signal_2909, KeyArray_S03reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_6_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2485, KeyArray_outS03ser[6]}), .a ({new_AGEMA_signal_2910, KeyArray_S03reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3297, KeyArray_S03reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2510, KeyArray_inS03ser[6]}), .a ({new_AGEMA_signal_2581, keySBIn[6]}), .c ({new_AGEMA_signal_2910, KeyArray_S03reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_7_U1 ( .s (KeyArray_n27), .b ({new_AGEMA_signal_2488, KeyArray_outS03ser[7]}), .a ({new_AGEMA_signal_2911, KeyArray_S03reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3298, KeyArray_S03reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n36), .b ({new_AGEMA_signal_2513, KeyArray_inS03ser[7]}), .a ({new_AGEMA_signal_2584, keySBIn[7]}), .c ({new_AGEMA_signal_2911, KeyArray_S03reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_0_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2491, KeyArray_outS10ser[0]}), .a ({new_AGEMA_signal_2912, KeyArray_S10reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3299, KeyArray_S10reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2516, KeyArray_inS10ser[0]}), .a ({new_AGEMA_signal_2587, KeyArray_outS20ser[0]}), .c ({new_AGEMA_signal_2912, KeyArray_S10reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_1_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2494, KeyArray_outS10ser[1]}), .a ({new_AGEMA_signal_2913, KeyArray_S10reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3300, KeyArray_S10reg_gff_1_SFF_1_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2519, KeyArray_inS10ser[1]}), .a ({new_AGEMA_signal_2590, KeyArray_outS20ser[1]}), .c ({new_AGEMA_signal_2913, KeyArray_S10reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_2_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2497, KeyArray_outS10ser[2]}), .a ({new_AGEMA_signal_2914, KeyArray_S10reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3301, KeyArray_S10reg_gff_1_SFF_2_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2522, KeyArray_inS10ser[2]}), .a ({new_AGEMA_signal_2593, KeyArray_outS20ser[2]}), .c ({new_AGEMA_signal_2914, KeyArray_S10reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_3_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2500, KeyArray_outS10ser[3]}), .a ({new_AGEMA_signal_2915, KeyArray_S10reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3302, KeyArray_S10reg_gff_1_SFF_3_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2525, KeyArray_inS10ser[3]}), .a ({new_AGEMA_signal_2596, KeyArray_outS20ser[3]}), .c ({new_AGEMA_signal_2915, KeyArray_S10reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_4_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2503, KeyArray_outS10ser[4]}), .a ({new_AGEMA_signal_2916, KeyArray_S10reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3303, KeyArray_S10reg_gff_1_SFF_4_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2528, KeyArray_inS10ser[4]}), .a ({new_AGEMA_signal_2599, KeyArray_outS20ser[4]}), .c ({new_AGEMA_signal_2916, KeyArray_S10reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_5_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2506, KeyArray_outS10ser[5]}), .a ({new_AGEMA_signal_2917, KeyArray_S10reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3304, KeyArray_S10reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2531, KeyArray_inS10ser[5]}), .a ({new_AGEMA_signal_2602, KeyArray_outS20ser[5]}), .c ({new_AGEMA_signal_2917, KeyArray_S10reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_6_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2509, KeyArray_outS10ser[6]}), .a ({new_AGEMA_signal_2918, KeyArray_S10reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3305, KeyArray_S10reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2534, KeyArray_inS10ser[6]}), .a ({new_AGEMA_signal_2605, KeyArray_outS20ser[6]}), .c ({new_AGEMA_signal_2918, KeyArray_S10reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_7_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2512, KeyArray_outS10ser[7]}), .a ({new_AGEMA_signal_2919, KeyArray_S10reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3306, KeyArray_S10reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2537, KeyArray_inS10ser[7]}), .a ({new_AGEMA_signal_2608, KeyArray_outS20ser[7]}), .c ({new_AGEMA_signal_2919, KeyArray_S10reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_0_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2515, KeyArray_outS11ser[0]}), .a ({new_AGEMA_signal_2920, KeyArray_S11reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3307, KeyArray_S11reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2540, KeyArray_inS11ser[0]}), .a ({new_AGEMA_signal_2611, KeyArray_outS21ser[0]}), .c ({new_AGEMA_signal_2920, KeyArray_S11reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_1_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2518, KeyArray_outS11ser[1]}), .a ({new_AGEMA_signal_2921, KeyArray_S11reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3308, KeyArray_S11reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2543, KeyArray_inS11ser[1]}), .a ({new_AGEMA_signal_2614, KeyArray_outS21ser[1]}), .c ({new_AGEMA_signal_2921, KeyArray_S11reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_2_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2521, KeyArray_outS11ser[2]}), .a ({new_AGEMA_signal_2922, KeyArray_S11reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3309, KeyArray_S11reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2546, KeyArray_inS11ser[2]}), .a ({new_AGEMA_signal_2617, KeyArray_outS21ser[2]}), .c ({new_AGEMA_signal_2922, KeyArray_S11reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_3_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2524, KeyArray_outS11ser[3]}), .a ({new_AGEMA_signal_2923, KeyArray_S11reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3310, KeyArray_S11reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2549, KeyArray_inS11ser[3]}), .a ({new_AGEMA_signal_2620, KeyArray_outS21ser[3]}), .c ({new_AGEMA_signal_2923, KeyArray_S11reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_4_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2527, KeyArray_outS11ser[4]}), .a ({new_AGEMA_signal_2924, KeyArray_S11reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3311, KeyArray_S11reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2552, KeyArray_inS11ser[4]}), .a ({new_AGEMA_signal_2623, KeyArray_outS21ser[4]}), .c ({new_AGEMA_signal_2924, KeyArray_S11reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_5_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2530, KeyArray_outS11ser[5]}), .a ({new_AGEMA_signal_2925, KeyArray_S11reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3312, KeyArray_S11reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2555, KeyArray_inS11ser[5]}), .a ({new_AGEMA_signal_2626, KeyArray_outS21ser[5]}), .c ({new_AGEMA_signal_2925, KeyArray_S11reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_6_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2533, KeyArray_outS11ser[6]}), .a ({new_AGEMA_signal_2926, KeyArray_S11reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3313, KeyArray_S11reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2558, KeyArray_inS11ser[6]}), .a ({new_AGEMA_signal_2629, KeyArray_outS21ser[6]}), .c ({new_AGEMA_signal_2926, KeyArray_S11reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_7_U1 ( .s (KeyArray_n26), .b ({new_AGEMA_signal_2536, KeyArray_outS11ser[7]}), .a ({new_AGEMA_signal_2927, KeyArray_S11reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3314, KeyArray_S11reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n35), .b ({new_AGEMA_signal_2561, KeyArray_inS11ser[7]}), .a ({new_AGEMA_signal_2632, KeyArray_outS21ser[7]}), .c ({new_AGEMA_signal_2927, KeyArray_S11reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_0_U1 ( .s (n12), .b ({new_AGEMA_signal_2539, KeyArray_outS12ser[0]}), .a ({new_AGEMA_signal_2928, KeyArray_S12reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3093, KeyArray_S12reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2564, KeyArray_inS12ser[0]}), .a ({new_AGEMA_signal_2635, KeyArray_outS22ser[0]}), .c ({new_AGEMA_signal_2928, KeyArray_S12reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_1_U1 ( .s (n12), .b ({new_AGEMA_signal_2542, KeyArray_outS12ser[1]}), .a ({new_AGEMA_signal_2929, KeyArray_S12reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3094, KeyArray_S12reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2567, KeyArray_inS12ser[1]}), .a ({new_AGEMA_signal_2638, KeyArray_outS22ser[1]}), .c ({new_AGEMA_signal_2929, KeyArray_S12reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_2_U1 ( .s (n12), .b ({new_AGEMA_signal_2545, KeyArray_outS12ser[2]}), .a ({new_AGEMA_signal_2930, KeyArray_S12reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3095, KeyArray_S12reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2570, KeyArray_inS12ser[2]}), .a ({new_AGEMA_signal_2641, KeyArray_outS22ser[2]}), .c ({new_AGEMA_signal_2930, KeyArray_S12reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_3_U1 ( .s (n12), .b ({new_AGEMA_signal_2548, KeyArray_outS12ser[3]}), .a ({new_AGEMA_signal_2931, KeyArray_S12reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3096, KeyArray_S12reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2573, KeyArray_inS12ser[3]}), .a ({new_AGEMA_signal_2644, KeyArray_outS22ser[3]}), .c ({new_AGEMA_signal_2931, KeyArray_S12reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_4_U1 ( .s (n12), .b ({new_AGEMA_signal_2551, KeyArray_outS12ser[4]}), .a ({new_AGEMA_signal_2932, KeyArray_S12reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3097, KeyArray_S12reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2576, KeyArray_inS12ser[4]}), .a ({new_AGEMA_signal_2647, KeyArray_outS22ser[4]}), .c ({new_AGEMA_signal_2932, KeyArray_S12reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_5_U1 ( .s (n12), .b ({new_AGEMA_signal_2554, KeyArray_outS12ser[5]}), .a ({new_AGEMA_signal_2933, KeyArray_S12reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3098, KeyArray_S12reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2579, KeyArray_inS12ser[5]}), .a ({new_AGEMA_signal_2650, KeyArray_outS22ser[5]}), .c ({new_AGEMA_signal_2933, KeyArray_S12reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_6_U1 ( .s (n12), .b ({new_AGEMA_signal_2557, KeyArray_outS12ser[6]}), .a ({new_AGEMA_signal_2934, KeyArray_S12reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3099, KeyArray_S12reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2582, KeyArray_inS12ser[6]}), .a ({new_AGEMA_signal_2653, KeyArray_outS22ser[6]}), .c ({new_AGEMA_signal_2934, KeyArray_S12reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_7_U1 ( .s (n12), .b ({new_AGEMA_signal_2560, KeyArray_outS12ser[7]}), .a ({new_AGEMA_signal_2935, KeyArray_S12reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3100, KeyArray_S12reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2585, KeyArray_inS12ser[7]}), .a ({new_AGEMA_signal_2656, KeyArray_outS22ser[7]}), .c ({new_AGEMA_signal_2935, KeyArray_S12reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_0_U1 ( .s (n12), .b ({new_AGEMA_signal_2563, keySBIn[0]}), .a ({new_AGEMA_signal_2936, KeyArray_S13reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3101, KeyArray_S13reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2588, KeyArray_inS13ser[0]}), .a ({new_AGEMA_signal_2659, KeyArray_outS23ser[0]}), .c ({new_AGEMA_signal_2936, KeyArray_S13reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_1_U1 ( .s (n12), .b ({new_AGEMA_signal_2566, keySBIn[1]}), .a ({new_AGEMA_signal_2937, KeyArray_S13reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3102, KeyArray_S13reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2591, KeyArray_inS13ser[1]}), .a ({new_AGEMA_signal_2662, KeyArray_outS23ser[1]}), .c ({new_AGEMA_signal_2937, KeyArray_S13reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_2_U1 ( .s (n12), .b ({new_AGEMA_signal_2569, keySBIn[2]}), .a ({new_AGEMA_signal_2938, KeyArray_S13reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3103, KeyArray_S13reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2594, KeyArray_inS13ser[2]}), .a ({new_AGEMA_signal_2665, KeyArray_outS23ser[2]}), .c ({new_AGEMA_signal_2938, KeyArray_S13reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_3_U1 ( .s (n12), .b ({new_AGEMA_signal_2572, keySBIn[3]}), .a ({new_AGEMA_signal_2939, KeyArray_S13reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3104, KeyArray_S13reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2597, KeyArray_inS13ser[3]}), .a ({new_AGEMA_signal_2668, KeyArray_outS23ser[3]}), .c ({new_AGEMA_signal_2939, KeyArray_S13reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_4_U1 ( .s (n12), .b ({new_AGEMA_signal_2575, keySBIn[4]}), .a ({new_AGEMA_signal_2940, KeyArray_S13reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3105, KeyArray_S13reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2600, KeyArray_inS13ser[4]}), .a ({new_AGEMA_signal_2671, KeyArray_outS23ser[4]}), .c ({new_AGEMA_signal_2940, KeyArray_S13reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_5_U1 ( .s (n12), .b ({new_AGEMA_signal_2578, keySBIn[5]}), .a ({new_AGEMA_signal_2941, KeyArray_S13reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3106, KeyArray_S13reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2603, KeyArray_inS13ser[5]}), .a ({new_AGEMA_signal_2674, KeyArray_outS23ser[5]}), .c ({new_AGEMA_signal_2941, KeyArray_S13reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_6_U1 ( .s (n12), .b ({new_AGEMA_signal_2581, keySBIn[6]}), .a ({new_AGEMA_signal_2942, KeyArray_S13reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3107, KeyArray_S13reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2606, KeyArray_inS13ser[6]}), .a ({new_AGEMA_signal_2677, KeyArray_outS23ser[6]}), .c ({new_AGEMA_signal_2942, KeyArray_S13reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_7_U1 ( .s (n12), .b ({new_AGEMA_signal_2584, keySBIn[7]}), .a ({new_AGEMA_signal_2943, KeyArray_S13reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3108, KeyArray_S13reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n34), .b ({new_AGEMA_signal_2609, KeyArray_inS13ser[7]}), .a ({new_AGEMA_signal_2680, KeyArray_outS23ser[7]}), .c ({new_AGEMA_signal_2943, KeyArray_S13reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_0_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2587, KeyArray_outS20ser[0]}), .a ({new_AGEMA_signal_2944, KeyArray_S20reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3315, KeyArray_S20reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2612, KeyArray_inS20ser[0]}), .a ({new_AGEMA_signal_2683, KeyArray_outS30ser[0]}), .c ({new_AGEMA_signal_2944, KeyArray_S20reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_1_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2590, KeyArray_outS20ser[1]}), .a ({new_AGEMA_signal_2945, KeyArray_S20reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3316, KeyArray_S20reg_gff_1_SFF_1_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2615, KeyArray_inS20ser[1]}), .a ({new_AGEMA_signal_2686, KeyArray_outS30ser[1]}), .c ({new_AGEMA_signal_2945, KeyArray_S20reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_2_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2593, KeyArray_outS20ser[2]}), .a ({new_AGEMA_signal_2946, KeyArray_S20reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3317, KeyArray_S20reg_gff_1_SFF_2_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2618, KeyArray_inS20ser[2]}), .a ({new_AGEMA_signal_2689, KeyArray_outS30ser[2]}), .c ({new_AGEMA_signal_2946, KeyArray_S20reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_3_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2596, KeyArray_outS20ser[3]}), .a ({new_AGEMA_signal_2947, KeyArray_S20reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3318, KeyArray_S20reg_gff_1_SFF_3_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2621, KeyArray_inS20ser[3]}), .a ({new_AGEMA_signal_2692, KeyArray_outS30ser[3]}), .c ({new_AGEMA_signal_2947, KeyArray_S20reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_4_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2599, KeyArray_outS20ser[4]}), .a ({new_AGEMA_signal_2948, KeyArray_S20reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3319, KeyArray_S20reg_gff_1_SFF_4_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2624, KeyArray_inS20ser[4]}), .a ({new_AGEMA_signal_2695, KeyArray_outS30ser[4]}), .c ({new_AGEMA_signal_2948, KeyArray_S20reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_5_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2602, KeyArray_outS20ser[5]}), .a ({new_AGEMA_signal_2949, KeyArray_S20reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3320, KeyArray_S20reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2627, KeyArray_inS20ser[5]}), .a ({new_AGEMA_signal_2698, KeyArray_outS30ser[5]}), .c ({new_AGEMA_signal_2949, KeyArray_S20reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_6_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2605, KeyArray_outS20ser[6]}), .a ({new_AGEMA_signal_2950, KeyArray_S20reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3321, KeyArray_S20reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2630, KeyArray_inS20ser[6]}), .a ({new_AGEMA_signal_2701, KeyArray_outS30ser[6]}), .c ({new_AGEMA_signal_2950, KeyArray_S20reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_7_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2608, KeyArray_outS20ser[7]}), .a ({new_AGEMA_signal_2951, KeyArray_S20reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3322, KeyArray_S20reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2633, KeyArray_inS20ser[7]}), .a ({new_AGEMA_signal_2704, KeyArray_outS30ser[7]}), .c ({new_AGEMA_signal_2951, KeyArray_S20reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_0_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2611, KeyArray_outS21ser[0]}), .a ({new_AGEMA_signal_2952, KeyArray_S21reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3323, KeyArray_S21reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2636, KeyArray_inS21ser[0]}), .a ({new_AGEMA_signal_2707, KeyArray_outS31ser[0]}), .c ({new_AGEMA_signal_2952, KeyArray_S21reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_1_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2614, KeyArray_outS21ser[1]}), .a ({new_AGEMA_signal_2953, KeyArray_S21reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3324, KeyArray_S21reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2639, KeyArray_inS21ser[1]}), .a ({new_AGEMA_signal_2710, KeyArray_outS31ser[1]}), .c ({new_AGEMA_signal_2953, KeyArray_S21reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_2_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2617, KeyArray_outS21ser[2]}), .a ({new_AGEMA_signal_2954, KeyArray_S21reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3325, KeyArray_S21reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2642, KeyArray_inS21ser[2]}), .a ({new_AGEMA_signal_2713, KeyArray_outS31ser[2]}), .c ({new_AGEMA_signal_2954, KeyArray_S21reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_3_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2620, KeyArray_outS21ser[3]}), .a ({new_AGEMA_signal_2955, KeyArray_S21reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3326, KeyArray_S21reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2645, KeyArray_inS21ser[3]}), .a ({new_AGEMA_signal_2716, KeyArray_outS31ser[3]}), .c ({new_AGEMA_signal_2955, KeyArray_S21reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_4_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2623, KeyArray_outS21ser[4]}), .a ({new_AGEMA_signal_2956, KeyArray_S21reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3327, KeyArray_S21reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2648, KeyArray_inS21ser[4]}), .a ({new_AGEMA_signal_2719, KeyArray_outS31ser[4]}), .c ({new_AGEMA_signal_2956, KeyArray_S21reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_5_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2626, KeyArray_outS21ser[5]}), .a ({new_AGEMA_signal_2957, KeyArray_S21reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3328, KeyArray_S21reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2651, KeyArray_inS21ser[5]}), .a ({new_AGEMA_signal_2722, KeyArray_outS31ser[5]}), .c ({new_AGEMA_signal_2957, KeyArray_S21reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_6_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2629, KeyArray_outS21ser[6]}), .a ({new_AGEMA_signal_2958, KeyArray_S21reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3329, KeyArray_S21reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2654, KeyArray_inS21ser[6]}), .a ({new_AGEMA_signal_2725, KeyArray_outS31ser[6]}), .c ({new_AGEMA_signal_2958, KeyArray_S21reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_7_U1 ( .s (KeyArray_n25), .b ({new_AGEMA_signal_2632, KeyArray_outS21ser[7]}), .a ({new_AGEMA_signal_2959, KeyArray_S21reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3330, KeyArray_S21reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n33), .b ({new_AGEMA_signal_2657, KeyArray_inS21ser[7]}), .a ({new_AGEMA_signal_2728, KeyArray_outS31ser[7]}), .c ({new_AGEMA_signal_2959, KeyArray_S21reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_0_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2635, KeyArray_outS22ser[0]}), .a ({new_AGEMA_signal_2960, KeyArray_S22reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3331, KeyArray_S22reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2660, KeyArray_inS22ser[0]}), .a ({new_AGEMA_signal_2731, KeyArray_outS32ser[0]}), .c ({new_AGEMA_signal_2960, KeyArray_S22reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_1_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2638, KeyArray_outS22ser[1]}), .a ({new_AGEMA_signal_2961, KeyArray_S22reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3332, KeyArray_S22reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2663, KeyArray_inS22ser[1]}), .a ({new_AGEMA_signal_2734, KeyArray_outS32ser[1]}), .c ({new_AGEMA_signal_2961, KeyArray_S22reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_2_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2641, KeyArray_outS22ser[2]}), .a ({new_AGEMA_signal_2962, KeyArray_S22reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3333, KeyArray_S22reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2666, KeyArray_inS22ser[2]}), .a ({new_AGEMA_signal_2737, KeyArray_outS32ser[2]}), .c ({new_AGEMA_signal_2962, KeyArray_S22reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_3_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2644, KeyArray_outS22ser[3]}), .a ({new_AGEMA_signal_2963, KeyArray_S22reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3334, KeyArray_S22reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2669, KeyArray_inS22ser[3]}), .a ({new_AGEMA_signal_2740, KeyArray_outS32ser[3]}), .c ({new_AGEMA_signal_2963, KeyArray_S22reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_4_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2647, KeyArray_outS22ser[4]}), .a ({new_AGEMA_signal_2964, KeyArray_S22reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3335, KeyArray_S22reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2672, KeyArray_inS22ser[4]}), .a ({new_AGEMA_signal_2743, KeyArray_outS32ser[4]}), .c ({new_AGEMA_signal_2964, KeyArray_S22reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_5_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2650, KeyArray_outS22ser[5]}), .a ({new_AGEMA_signal_2965, KeyArray_S22reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3336, KeyArray_S22reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2675, KeyArray_inS22ser[5]}), .a ({new_AGEMA_signal_2746, KeyArray_outS32ser[5]}), .c ({new_AGEMA_signal_2965, KeyArray_S22reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_6_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2653, KeyArray_outS22ser[6]}), .a ({new_AGEMA_signal_2966, KeyArray_S22reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3337, KeyArray_S22reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2678, KeyArray_inS22ser[6]}), .a ({new_AGEMA_signal_2749, KeyArray_outS32ser[6]}), .c ({new_AGEMA_signal_2966, KeyArray_S22reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_7_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2656, KeyArray_outS22ser[7]}), .a ({new_AGEMA_signal_2967, KeyArray_S22reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3338, KeyArray_S22reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2681, KeyArray_inS22ser[7]}), .a ({new_AGEMA_signal_2752, KeyArray_outS32ser[7]}), .c ({new_AGEMA_signal_2967, KeyArray_S22reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_0_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2659, KeyArray_outS23ser[0]}), .a ({new_AGEMA_signal_2968, KeyArray_S23reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3339, KeyArray_S23reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2684, KeyArray_inS23ser[0]}), .a ({new_AGEMA_signal_2755, KeyArray_outS33ser[0]}), .c ({new_AGEMA_signal_2968, KeyArray_S23reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_1_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2662, KeyArray_outS23ser[1]}), .a ({new_AGEMA_signal_2969, KeyArray_S23reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3340, KeyArray_S23reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2687, KeyArray_inS23ser[1]}), .a ({new_AGEMA_signal_2758, KeyArray_outS33ser[1]}), .c ({new_AGEMA_signal_2969, KeyArray_S23reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_2_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2665, KeyArray_outS23ser[2]}), .a ({new_AGEMA_signal_2970, KeyArray_S23reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3341, KeyArray_S23reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2690, KeyArray_inS23ser[2]}), .a ({new_AGEMA_signal_2761, KeyArray_outS33ser[2]}), .c ({new_AGEMA_signal_2970, KeyArray_S23reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_3_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2668, KeyArray_outS23ser[3]}), .a ({new_AGEMA_signal_2971, KeyArray_S23reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3342, KeyArray_S23reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2693, KeyArray_inS23ser[3]}), .a ({new_AGEMA_signal_2764, KeyArray_outS33ser[3]}), .c ({new_AGEMA_signal_2971, KeyArray_S23reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_4_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2671, KeyArray_outS23ser[4]}), .a ({new_AGEMA_signal_2972, KeyArray_S23reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3343, KeyArray_S23reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2696, KeyArray_inS23ser[4]}), .a ({new_AGEMA_signal_2767, KeyArray_outS33ser[4]}), .c ({new_AGEMA_signal_2972, KeyArray_S23reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_5_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2674, KeyArray_outS23ser[5]}), .a ({new_AGEMA_signal_2973, KeyArray_S23reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3344, KeyArray_S23reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2699, KeyArray_inS23ser[5]}), .a ({new_AGEMA_signal_2770, KeyArray_outS33ser[5]}), .c ({new_AGEMA_signal_2973, KeyArray_S23reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_6_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2677, KeyArray_outS23ser[6]}), .a ({new_AGEMA_signal_2974, KeyArray_S23reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3345, KeyArray_S23reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2702, KeyArray_inS23ser[6]}), .a ({new_AGEMA_signal_2773, KeyArray_outS33ser[6]}), .c ({new_AGEMA_signal_2974, KeyArray_S23reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_7_U1 ( .s (KeyArray_n24), .b ({new_AGEMA_signal_2680, KeyArray_outS23ser[7]}), .a ({new_AGEMA_signal_2975, KeyArray_S23reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3346, KeyArray_S23reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n32), .b ({new_AGEMA_signal_2705, KeyArray_inS23ser[7]}), .a ({new_AGEMA_signal_2776, KeyArray_outS33ser[7]}), .c ({new_AGEMA_signal_2975, KeyArray_S23reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_0_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2707, KeyArray_outS31ser[0]}), .a ({new_AGEMA_signal_2976, KeyArray_S31reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3347, KeyArray_S31reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2732, KeyArray_inS31ser[0]}), .a ({new_AGEMA_signal_2020, KeyArray_outS01ser_0_}), .c ({new_AGEMA_signal_2976, KeyArray_S31reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_1_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2710, KeyArray_outS31ser[1]}), .a ({new_AGEMA_signal_2977, KeyArray_S31reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3348, KeyArray_S31reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2735, KeyArray_inS31ser[1]}), .a ({new_AGEMA_signal_2018, KeyArray_outS01ser_1_}), .c ({new_AGEMA_signal_2977, KeyArray_S31reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_2_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2713, KeyArray_outS31ser[2]}), .a ({new_AGEMA_signal_2978, KeyArray_S31reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3349, KeyArray_S31reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2738, KeyArray_inS31ser[2]}), .a ({new_AGEMA_signal_2016, KeyArray_outS01ser_2_}), .c ({new_AGEMA_signal_2978, KeyArray_S31reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_3_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2716, KeyArray_outS31ser[3]}), .a ({new_AGEMA_signal_2979, KeyArray_S31reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3350, KeyArray_S31reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2741, KeyArray_inS31ser[3]}), .a ({new_AGEMA_signal_2014, KeyArray_outS01ser_3_}), .c ({new_AGEMA_signal_2979, KeyArray_S31reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_4_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2719, KeyArray_outS31ser[4]}), .a ({new_AGEMA_signal_2980, KeyArray_S31reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3351, KeyArray_S31reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2744, KeyArray_inS31ser[4]}), .a ({new_AGEMA_signal_2012, KeyArray_outS01ser_4_}), .c ({new_AGEMA_signal_2980, KeyArray_S31reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_5_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2722, KeyArray_outS31ser[5]}), .a ({new_AGEMA_signal_2981, KeyArray_S31reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3352, KeyArray_S31reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2747, KeyArray_inS31ser[5]}), .a ({new_AGEMA_signal_2010, KeyArray_outS01ser_5_}), .c ({new_AGEMA_signal_2981, KeyArray_S31reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_6_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2725, KeyArray_outS31ser[6]}), .a ({new_AGEMA_signal_2982, KeyArray_S31reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3353, KeyArray_S31reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2750, KeyArray_inS31ser[6]}), .a ({new_AGEMA_signal_2008, KeyArray_outS01ser_6_}), .c ({new_AGEMA_signal_2982, KeyArray_S31reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_7_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2728, KeyArray_outS31ser[7]}), .a ({new_AGEMA_signal_2983, KeyArray_S31reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3354, KeyArray_S31reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2753, KeyArray_inS31ser[7]}), .a ({new_AGEMA_signal_2006, KeyArray_outS01ser_7_}), .c ({new_AGEMA_signal_2983, KeyArray_S31reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_0_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2731, KeyArray_outS32ser[0]}), .a ({new_AGEMA_signal_2984, KeyArray_S32reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3355, KeyArray_S32reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2756, KeyArray_inS32ser[0]}), .a ({new_AGEMA_signal_2443, KeyArray_outS02ser[0]}), .c ({new_AGEMA_signal_2984, KeyArray_S32reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_1_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2734, KeyArray_outS32ser[1]}), .a ({new_AGEMA_signal_2985, KeyArray_S32reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3356, KeyArray_S32reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2759, KeyArray_inS32ser[1]}), .a ({new_AGEMA_signal_2446, KeyArray_outS02ser[1]}), .c ({new_AGEMA_signal_2985, KeyArray_S32reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_2_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2737, KeyArray_outS32ser[2]}), .a ({new_AGEMA_signal_2986, KeyArray_S32reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3357, KeyArray_S32reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2762, KeyArray_inS32ser[2]}), .a ({new_AGEMA_signal_2449, KeyArray_outS02ser[2]}), .c ({new_AGEMA_signal_2986, KeyArray_S32reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_3_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2740, KeyArray_outS32ser[3]}), .a ({new_AGEMA_signal_2987, KeyArray_S32reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3358, KeyArray_S32reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2765, KeyArray_inS32ser[3]}), .a ({new_AGEMA_signal_2452, KeyArray_outS02ser[3]}), .c ({new_AGEMA_signal_2987, KeyArray_S32reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_4_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2743, KeyArray_outS32ser[4]}), .a ({new_AGEMA_signal_2988, KeyArray_S32reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3359, KeyArray_S32reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2768, KeyArray_inS32ser[4]}), .a ({new_AGEMA_signal_2455, KeyArray_outS02ser[4]}), .c ({new_AGEMA_signal_2988, KeyArray_S32reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_5_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2746, KeyArray_outS32ser[5]}), .a ({new_AGEMA_signal_2989, KeyArray_S32reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3360, KeyArray_S32reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2771, KeyArray_inS32ser[5]}), .a ({new_AGEMA_signal_2458, KeyArray_outS02ser[5]}), .c ({new_AGEMA_signal_2989, KeyArray_S32reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_6_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2749, KeyArray_outS32ser[6]}), .a ({new_AGEMA_signal_2990, KeyArray_S32reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3361, KeyArray_S32reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2774, KeyArray_inS32ser[6]}), .a ({new_AGEMA_signal_2461, KeyArray_outS02ser[6]}), .c ({new_AGEMA_signal_2990, KeyArray_S32reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_7_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2752, KeyArray_outS32ser[7]}), .a ({new_AGEMA_signal_2991, KeyArray_S32reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3362, KeyArray_S32reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2777, KeyArray_inS32ser[7]}), .a ({new_AGEMA_signal_2464, KeyArray_outS02ser[7]}), .c ({new_AGEMA_signal_2991, KeyArray_S32reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_0_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2755, KeyArray_outS33ser[0]}), .a ({new_AGEMA_signal_2992, KeyArray_S33reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3363, KeyArray_S33reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2779, KeyArray_inS33ser[0]}), .a ({new_AGEMA_signal_2467, KeyArray_outS03ser[0]}), .c ({new_AGEMA_signal_2992, KeyArray_S33reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_1_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2758, KeyArray_outS33ser[1]}), .a ({new_AGEMA_signal_2993, KeyArray_S33reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3364, KeyArray_S33reg_gff_1_SFF_1_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2781, KeyArray_inS33ser[1]}), .a ({new_AGEMA_signal_2470, KeyArray_outS03ser[1]}), .c ({new_AGEMA_signal_2993, KeyArray_S33reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_2_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2761, KeyArray_outS33ser[2]}), .a ({new_AGEMA_signal_2994, KeyArray_S33reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3365, KeyArray_S33reg_gff_1_SFF_2_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2783, KeyArray_inS33ser[2]}), .a ({new_AGEMA_signal_2473, KeyArray_outS03ser[2]}), .c ({new_AGEMA_signal_2994, KeyArray_S33reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_3_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2764, KeyArray_outS33ser[3]}), .a ({new_AGEMA_signal_2995, KeyArray_S33reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3366, KeyArray_S33reg_gff_1_SFF_3_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2785, KeyArray_inS33ser[3]}), .a ({new_AGEMA_signal_2476, KeyArray_outS03ser[3]}), .c ({new_AGEMA_signal_2995, KeyArray_S33reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_4_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2767, KeyArray_outS33ser[4]}), .a ({new_AGEMA_signal_2996, KeyArray_S33reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3367, KeyArray_S33reg_gff_1_SFF_4_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2787, KeyArray_inS33ser[4]}), .a ({new_AGEMA_signal_2479, KeyArray_outS03ser[4]}), .c ({new_AGEMA_signal_2996, KeyArray_S33reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_5_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2770, KeyArray_outS33ser[5]}), .a ({new_AGEMA_signal_2997, KeyArray_S33reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3368, KeyArray_S33reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2789, KeyArray_inS33ser[5]}), .a ({new_AGEMA_signal_2482, KeyArray_outS03ser[5]}), .c ({new_AGEMA_signal_2997, KeyArray_S33reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_6_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2773, KeyArray_outS33ser[6]}), .a ({new_AGEMA_signal_2998, KeyArray_S33reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3369, KeyArray_S33reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2791, KeyArray_inS33ser[6]}), .a ({new_AGEMA_signal_2485, KeyArray_outS03ser[6]}), .c ({new_AGEMA_signal_2998, KeyArray_S33reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_7_U1 ( .s (KeyArray_n22), .b ({new_AGEMA_signal_2776, KeyArray_outS33ser[7]}), .a ({new_AGEMA_signal_2999, KeyArray_S33reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3370, KeyArray_S33reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n30), .b ({new_AGEMA_signal_2793, KeyArray_inS33ser[7]}), .a ({new_AGEMA_signal_2488, KeyArray_outS03ser[7]}), .c ({new_AGEMA_signal_2999, KeyArray_S33reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_selXOR_mux_inst_0_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2020, KeyArray_outS01ser_0_}), .a ({new_AGEMA_signal_2021, KeyArray_outS01ser_XOR_00[0]}), .c ({new_AGEMA_signal_3109, KeyArray_outS01ser_p[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_selXOR_mux_inst_1_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2018, KeyArray_outS01ser_1_}), .a ({new_AGEMA_signal_2019, KeyArray_outS01ser_XOR_00[1]}), .c ({new_AGEMA_signal_3110, KeyArray_outS01ser_p[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_selXOR_mux_inst_2_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2016, KeyArray_outS01ser_2_}), .a ({new_AGEMA_signal_2017, KeyArray_outS01ser_XOR_00[2]}), .c ({new_AGEMA_signal_3111, KeyArray_outS01ser_p[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_selXOR_mux_inst_3_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2014, KeyArray_outS01ser_3_}), .a ({new_AGEMA_signal_2015, KeyArray_outS01ser_XOR_00[3]}), .c ({new_AGEMA_signal_3112, KeyArray_outS01ser_p[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_selXOR_mux_inst_4_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2012, KeyArray_outS01ser_4_}), .a ({new_AGEMA_signal_2013, KeyArray_outS01ser_XOR_00[4]}), .c ({new_AGEMA_signal_3113, KeyArray_outS01ser_p[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_selXOR_mux_inst_5_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2010, KeyArray_outS01ser_5_}), .a ({new_AGEMA_signal_2011, KeyArray_outS01ser_XOR_00[5]}), .c ({new_AGEMA_signal_3114, KeyArray_outS01ser_p[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_selXOR_mux_inst_6_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2008, KeyArray_outS01ser_6_}), .a ({new_AGEMA_signal_2009, KeyArray_outS01ser_XOR_00[6]}), .c ({new_AGEMA_signal_3115, KeyArray_outS01ser_p[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_selXOR_mux_inst_7_U1 ( .s (intselXOR), .b ({new_AGEMA_signal_2006, KeyArray_outS01ser_7_}), .a ({new_AGEMA_signal_2007, KeyArray_outS01ser_XOR_00[7]}), .c ({new_AGEMA_signal_3116, KeyArray_outS01ser_p[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS00ser_mux_inst_0_U1 ( .s (KeyArray_n46), .b ({key_s1[120], key_s0[120]}), .a ({new_AGEMA_signal_3109, KeyArray_outS01ser_p[0]}), .c ({new_AGEMA_signal_3247, KeyArray_inS00ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS00ser_mux_inst_1_U1 ( .s (KeyArray_n46), .b ({key_s1[121], key_s0[121]}), .a ({new_AGEMA_signal_3110, KeyArray_outS01ser_p[1]}), .c ({new_AGEMA_signal_3249, KeyArray_inS00ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS00ser_mux_inst_2_U1 ( .s (KeyArray_n46), .b ({key_s1[122], key_s0[122]}), .a ({new_AGEMA_signal_3111, KeyArray_outS01ser_p[2]}), .c ({new_AGEMA_signal_3251, KeyArray_inS00ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS00ser_mux_inst_3_U1 ( .s (KeyArray_n46), .b ({key_s1[123], key_s0[123]}), .a ({new_AGEMA_signal_3112, KeyArray_outS01ser_p[3]}), .c ({new_AGEMA_signal_3253, KeyArray_inS00ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS00ser_mux_inst_4_U1 ( .s (KeyArray_n46), .b ({key_s1[124], key_s0[124]}), .a ({new_AGEMA_signal_3113, KeyArray_outS01ser_p[4]}), .c ({new_AGEMA_signal_3255, KeyArray_inS00ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS00ser_mux_inst_5_U1 ( .s (KeyArray_n46), .b ({key_s1[125], key_s0[125]}), .a ({new_AGEMA_signal_3114, KeyArray_outS01ser_p[5]}), .c ({new_AGEMA_signal_3257, KeyArray_inS00ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS00ser_mux_inst_6_U1 ( .s (KeyArray_n46), .b ({key_s1[126], key_s0[126]}), .a ({new_AGEMA_signal_3115, KeyArray_outS01ser_p[6]}), .c ({new_AGEMA_signal_3259, KeyArray_inS00ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS00ser_mux_inst_7_U1 ( .s (KeyArray_n46), .b ({key_s1[127], key_s0[127]}), .a ({new_AGEMA_signal_3116, KeyArray_outS01ser_p[7]}), .c ({new_AGEMA_signal_3261, KeyArray_inS00ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS01ser_mux_inst_0_U1 ( .s (KeyArray_n46), .b ({key_s1[112], key_s0[112]}), .a ({new_AGEMA_signal_2443, KeyArray_outS02ser[0]}), .c ({new_AGEMA_signal_2444, KeyArray_inS01ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS01ser_mux_inst_1_U1 ( .s (KeyArray_n46), .b ({key_s1[113], key_s0[113]}), .a ({new_AGEMA_signal_2446, KeyArray_outS02ser[1]}), .c ({new_AGEMA_signal_2447, KeyArray_inS01ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS01ser_mux_inst_2_U1 ( .s (KeyArray_n46), .b ({key_s1[114], key_s0[114]}), .a ({new_AGEMA_signal_2449, KeyArray_outS02ser[2]}), .c ({new_AGEMA_signal_2450, KeyArray_inS01ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS01ser_mux_inst_3_U1 ( .s (KeyArray_n46), .b ({key_s1[115], key_s0[115]}), .a ({new_AGEMA_signal_2452, KeyArray_outS02ser[3]}), .c ({new_AGEMA_signal_2453, KeyArray_inS01ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS01ser_mux_inst_4_U1 ( .s (KeyArray_n46), .b ({key_s1[116], key_s0[116]}), .a ({new_AGEMA_signal_2455, KeyArray_outS02ser[4]}), .c ({new_AGEMA_signal_2456, KeyArray_inS01ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS01ser_mux_inst_5_U1 ( .s (KeyArray_n46), .b ({key_s1[117], key_s0[117]}), .a ({new_AGEMA_signal_2458, KeyArray_outS02ser[5]}), .c ({new_AGEMA_signal_2459, KeyArray_inS01ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS01ser_mux_inst_6_U1 ( .s (KeyArray_n46), .b ({key_s1[118], key_s0[118]}), .a ({new_AGEMA_signal_2461, KeyArray_outS02ser[6]}), .c ({new_AGEMA_signal_2462, KeyArray_inS01ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS01ser_mux_inst_7_U1 ( .s (KeyArray_n46), .b ({key_s1[119], key_s0[119]}), .a ({new_AGEMA_signal_2464, KeyArray_outS02ser[7]}), .c ({new_AGEMA_signal_2465, KeyArray_inS01ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS02ser_mux_inst_0_U1 ( .s (KeyArray_n45), .b ({key_s1[104], key_s0[104]}), .a ({new_AGEMA_signal_2467, KeyArray_outS03ser[0]}), .c ({new_AGEMA_signal_2468, KeyArray_inS02ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS02ser_mux_inst_1_U1 ( .s (KeyArray_n45), .b ({key_s1[105], key_s0[105]}), .a ({new_AGEMA_signal_2470, KeyArray_outS03ser[1]}), .c ({new_AGEMA_signal_2471, KeyArray_inS02ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS02ser_mux_inst_2_U1 ( .s (KeyArray_n45), .b ({key_s1[106], key_s0[106]}), .a ({new_AGEMA_signal_2473, KeyArray_outS03ser[2]}), .c ({new_AGEMA_signal_2474, KeyArray_inS02ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS02ser_mux_inst_3_U1 ( .s (KeyArray_n45), .b ({key_s1[107], key_s0[107]}), .a ({new_AGEMA_signal_2476, KeyArray_outS03ser[3]}), .c ({new_AGEMA_signal_2477, KeyArray_inS02ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS02ser_mux_inst_4_U1 ( .s (KeyArray_n45), .b ({key_s1[108], key_s0[108]}), .a ({new_AGEMA_signal_2479, KeyArray_outS03ser[4]}), .c ({new_AGEMA_signal_2480, KeyArray_inS02ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS02ser_mux_inst_5_U1 ( .s (KeyArray_n45), .b ({key_s1[109], key_s0[109]}), .a ({new_AGEMA_signal_2482, KeyArray_outS03ser[5]}), .c ({new_AGEMA_signal_2483, KeyArray_inS02ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS02ser_mux_inst_6_U1 ( .s (KeyArray_n45), .b ({key_s1[110], key_s0[110]}), .a ({new_AGEMA_signal_2485, KeyArray_outS03ser[6]}), .c ({new_AGEMA_signal_2486, KeyArray_inS02ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS02ser_mux_inst_7_U1 ( .s (KeyArray_n45), .b ({key_s1[111], key_s0[111]}), .a ({new_AGEMA_signal_2488, KeyArray_outS03ser[7]}), .c ({new_AGEMA_signal_2489, KeyArray_inS02ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS03ser_mux_inst_0_U1 ( .s (KeyArray_n45), .b ({key_s1[96], key_s0[96]}), .a ({new_AGEMA_signal_2491, KeyArray_outS10ser[0]}), .c ({new_AGEMA_signal_2492, KeyArray_inS03ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS03ser_mux_inst_1_U1 ( .s (KeyArray_n45), .b ({key_s1[97], key_s0[97]}), .a ({new_AGEMA_signal_2494, KeyArray_outS10ser[1]}), .c ({new_AGEMA_signal_2495, KeyArray_inS03ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS03ser_mux_inst_2_U1 ( .s (KeyArray_n45), .b ({key_s1[98], key_s0[98]}), .a ({new_AGEMA_signal_2497, KeyArray_outS10ser[2]}), .c ({new_AGEMA_signal_2498, KeyArray_inS03ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS03ser_mux_inst_3_U1 ( .s (KeyArray_n45), .b ({key_s1[99], key_s0[99]}), .a ({new_AGEMA_signal_2500, KeyArray_outS10ser[3]}), .c ({new_AGEMA_signal_2501, KeyArray_inS03ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS03ser_mux_inst_4_U1 ( .s (KeyArray_n45), .b ({key_s1[100], key_s0[100]}), .a ({new_AGEMA_signal_2503, KeyArray_outS10ser[4]}), .c ({new_AGEMA_signal_2504, KeyArray_inS03ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS03ser_mux_inst_5_U1 ( .s (KeyArray_n45), .b ({key_s1[101], key_s0[101]}), .a ({new_AGEMA_signal_2506, KeyArray_outS10ser[5]}), .c ({new_AGEMA_signal_2507, KeyArray_inS03ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS03ser_mux_inst_6_U1 ( .s (KeyArray_n45), .b ({key_s1[102], key_s0[102]}), .a ({new_AGEMA_signal_2509, KeyArray_outS10ser[6]}), .c ({new_AGEMA_signal_2510, KeyArray_inS03ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS03ser_mux_inst_7_U1 ( .s (KeyArray_n45), .b ({key_s1[103], key_s0[103]}), .a ({new_AGEMA_signal_2512, KeyArray_outS10ser[7]}), .c ({new_AGEMA_signal_2513, KeyArray_inS03ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS10ser_mux_inst_0_U1 ( .s (KeyArray_n44), .b ({key_s1[88], key_s0[88]}), .a ({new_AGEMA_signal_2515, KeyArray_outS11ser[0]}), .c ({new_AGEMA_signal_2516, KeyArray_inS10ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS10ser_mux_inst_1_U1 ( .s (KeyArray_n44), .b ({key_s1[89], key_s0[89]}), .a ({new_AGEMA_signal_2518, KeyArray_outS11ser[1]}), .c ({new_AGEMA_signal_2519, KeyArray_inS10ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS10ser_mux_inst_2_U1 ( .s (KeyArray_n44), .b ({key_s1[90], key_s0[90]}), .a ({new_AGEMA_signal_2521, KeyArray_outS11ser[2]}), .c ({new_AGEMA_signal_2522, KeyArray_inS10ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS10ser_mux_inst_3_U1 ( .s (KeyArray_n44), .b ({key_s1[91], key_s0[91]}), .a ({new_AGEMA_signal_2524, KeyArray_outS11ser[3]}), .c ({new_AGEMA_signal_2525, KeyArray_inS10ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS10ser_mux_inst_4_U1 ( .s (KeyArray_n44), .b ({key_s1[92], key_s0[92]}), .a ({new_AGEMA_signal_2527, KeyArray_outS11ser[4]}), .c ({new_AGEMA_signal_2528, KeyArray_inS10ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS10ser_mux_inst_5_U1 ( .s (KeyArray_n44), .b ({key_s1[93], key_s0[93]}), .a ({new_AGEMA_signal_2530, KeyArray_outS11ser[5]}), .c ({new_AGEMA_signal_2531, KeyArray_inS10ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS10ser_mux_inst_6_U1 ( .s (KeyArray_n44), .b ({key_s1[94], key_s0[94]}), .a ({new_AGEMA_signal_2533, KeyArray_outS11ser[6]}), .c ({new_AGEMA_signal_2534, KeyArray_inS10ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS10ser_mux_inst_7_U1 ( .s (KeyArray_n44), .b ({key_s1[95], key_s0[95]}), .a ({new_AGEMA_signal_2536, KeyArray_outS11ser[7]}), .c ({new_AGEMA_signal_2537, KeyArray_inS10ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS11ser_mux_inst_0_U1 ( .s (KeyArray_n44), .b ({key_s1[80], key_s0[80]}), .a ({new_AGEMA_signal_2539, KeyArray_outS12ser[0]}), .c ({new_AGEMA_signal_2540, KeyArray_inS11ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS11ser_mux_inst_1_U1 ( .s (KeyArray_n44), .b ({key_s1[81], key_s0[81]}), .a ({new_AGEMA_signal_2542, KeyArray_outS12ser[1]}), .c ({new_AGEMA_signal_2543, KeyArray_inS11ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS11ser_mux_inst_2_U1 ( .s (KeyArray_n44), .b ({key_s1[82], key_s0[82]}), .a ({new_AGEMA_signal_2545, KeyArray_outS12ser[2]}), .c ({new_AGEMA_signal_2546, KeyArray_inS11ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS11ser_mux_inst_3_U1 ( .s (KeyArray_n44), .b ({key_s1[83], key_s0[83]}), .a ({new_AGEMA_signal_2548, KeyArray_outS12ser[3]}), .c ({new_AGEMA_signal_2549, KeyArray_inS11ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS11ser_mux_inst_4_U1 ( .s (KeyArray_n44), .b ({key_s1[84], key_s0[84]}), .a ({new_AGEMA_signal_2551, KeyArray_outS12ser[4]}), .c ({new_AGEMA_signal_2552, KeyArray_inS11ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS11ser_mux_inst_5_U1 ( .s (KeyArray_n44), .b ({key_s1[85], key_s0[85]}), .a ({new_AGEMA_signal_2554, KeyArray_outS12ser[5]}), .c ({new_AGEMA_signal_2555, KeyArray_inS11ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS11ser_mux_inst_6_U1 ( .s (KeyArray_n44), .b ({key_s1[86], key_s0[86]}), .a ({new_AGEMA_signal_2557, KeyArray_outS12ser[6]}), .c ({new_AGEMA_signal_2558, KeyArray_inS11ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS11ser_mux_inst_7_U1 ( .s (KeyArray_n44), .b ({key_s1[87], key_s0[87]}), .a ({new_AGEMA_signal_2560, KeyArray_outS12ser[7]}), .c ({new_AGEMA_signal_2561, KeyArray_inS11ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS12ser_mux_inst_0_U1 ( .s (KeyArray_n43), .b ({key_s1[72], key_s0[72]}), .a ({new_AGEMA_signal_2563, keySBIn[0]}), .c ({new_AGEMA_signal_2564, KeyArray_inS12ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS12ser_mux_inst_1_U1 ( .s (KeyArray_n43), .b ({key_s1[73], key_s0[73]}), .a ({new_AGEMA_signal_2566, keySBIn[1]}), .c ({new_AGEMA_signal_2567, KeyArray_inS12ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS12ser_mux_inst_2_U1 ( .s (KeyArray_n43), .b ({key_s1[74], key_s0[74]}), .a ({new_AGEMA_signal_2569, keySBIn[2]}), .c ({new_AGEMA_signal_2570, KeyArray_inS12ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS12ser_mux_inst_3_U1 ( .s (KeyArray_n43), .b ({key_s1[75], key_s0[75]}), .a ({new_AGEMA_signal_2572, keySBIn[3]}), .c ({new_AGEMA_signal_2573, KeyArray_inS12ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS12ser_mux_inst_4_U1 ( .s (KeyArray_n43), .b ({key_s1[76], key_s0[76]}), .a ({new_AGEMA_signal_2575, keySBIn[4]}), .c ({new_AGEMA_signal_2576, KeyArray_inS12ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS12ser_mux_inst_5_U1 ( .s (KeyArray_n43), .b ({key_s1[77], key_s0[77]}), .a ({new_AGEMA_signal_2578, keySBIn[5]}), .c ({new_AGEMA_signal_2579, KeyArray_inS12ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS12ser_mux_inst_6_U1 ( .s (KeyArray_n43), .b ({key_s1[78], key_s0[78]}), .a ({new_AGEMA_signal_2581, keySBIn[6]}), .c ({new_AGEMA_signal_2582, KeyArray_inS12ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS12ser_mux_inst_7_U1 ( .s (KeyArray_n43), .b ({key_s1[79], key_s0[79]}), .a ({new_AGEMA_signal_2584, keySBIn[7]}), .c ({new_AGEMA_signal_2585, KeyArray_inS12ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS13ser_mux_inst_0_U1 ( .s (KeyArray_n43), .b ({key_s1[64], key_s0[64]}), .a ({new_AGEMA_signal_2587, KeyArray_outS20ser[0]}), .c ({new_AGEMA_signal_2588, KeyArray_inS13ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS13ser_mux_inst_1_U1 ( .s (KeyArray_n43), .b ({key_s1[65], key_s0[65]}), .a ({new_AGEMA_signal_2590, KeyArray_outS20ser[1]}), .c ({new_AGEMA_signal_2591, KeyArray_inS13ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS13ser_mux_inst_2_U1 ( .s (KeyArray_n43), .b ({key_s1[66], key_s0[66]}), .a ({new_AGEMA_signal_2593, KeyArray_outS20ser[2]}), .c ({new_AGEMA_signal_2594, KeyArray_inS13ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS13ser_mux_inst_3_U1 ( .s (KeyArray_n43), .b ({key_s1[67], key_s0[67]}), .a ({new_AGEMA_signal_2596, KeyArray_outS20ser[3]}), .c ({new_AGEMA_signal_2597, KeyArray_inS13ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS13ser_mux_inst_4_U1 ( .s (KeyArray_n43), .b ({key_s1[68], key_s0[68]}), .a ({new_AGEMA_signal_2599, KeyArray_outS20ser[4]}), .c ({new_AGEMA_signal_2600, KeyArray_inS13ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS13ser_mux_inst_5_U1 ( .s (KeyArray_n43), .b ({key_s1[69], key_s0[69]}), .a ({new_AGEMA_signal_2602, KeyArray_outS20ser[5]}), .c ({new_AGEMA_signal_2603, KeyArray_inS13ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS13ser_mux_inst_6_U1 ( .s (KeyArray_n43), .b ({key_s1[70], key_s0[70]}), .a ({new_AGEMA_signal_2605, KeyArray_outS20ser[6]}), .c ({new_AGEMA_signal_2606, KeyArray_inS13ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS13ser_mux_inst_7_U1 ( .s (KeyArray_n43), .b ({key_s1[71], key_s0[71]}), .a ({new_AGEMA_signal_2608, KeyArray_outS20ser[7]}), .c ({new_AGEMA_signal_2609, KeyArray_inS13ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS20ser_mux_inst_0_U1 ( .s (KeyArray_n42), .b ({key_s1[56], key_s0[56]}), .a ({new_AGEMA_signal_2611, KeyArray_outS21ser[0]}), .c ({new_AGEMA_signal_2612, KeyArray_inS20ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS20ser_mux_inst_1_U1 ( .s (KeyArray_n42), .b ({key_s1[57], key_s0[57]}), .a ({new_AGEMA_signal_2614, KeyArray_outS21ser[1]}), .c ({new_AGEMA_signal_2615, KeyArray_inS20ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS20ser_mux_inst_2_U1 ( .s (KeyArray_n42), .b ({key_s1[58], key_s0[58]}), .a ({new_AGEMA_signal_2617, KeyArray_outS21ser[2]}), .c ({new_AGEMA_signal_2618, KeyArray_inS20ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS20ser_mux_inst_3_U1 ( .s (KeyArray_n42), .b ({key_s1[59], key_s0[59]}), .a ({new_AGEMA_signal_2620, KeyArray_outS21ser[3]}), .c ({new_AGEMA_signal_2621, KeyArray_inS20ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS20ser_mux_inst_4_U1 ( .s (KeyArray_n42), .b ({key_s1[60], key_s0[60]}), .a ({new_AGEMA_signal_2623, KeyArray_outS21ser[4]}), .c ({new_AGEMA_signal_2624, KeyArray_inS20ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS20ser_mux_inst_5_U1 ( .s (KeyArray_n42), .b ({key_s1[61], key_s0[61]}), .a ({new_AGEMA_signal_2626, KeyArray_outS21ser[5]}), .c ({new_AGEMA_signal_2627, KeyArray_inS20ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS20ser_mux_inst_6_U1 ( .s (KeyArray_n42), .b ({key_s1[62], key_s0[62]}), .a ({new_AGEMA_signal_2629, KeyArray_outS21ser[6]}), .c ({new_AGEMA_signal_2630, KeyArray_inS20ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS20ser_mux_inst_7_U1 ( .s (KeyArray_n42), .b ({key_s1[63], key_s0[63]}), .a ({new_AGEMA_signal_2632, KeyArray_outS21ser[7]}), .c ({new_AGEMA_signal_2633, KeyArray_inS20ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS21ser_mux_inst_0_U1 ( .s (KeyArray_n42), .b ({key_s1[48], key_s0[48]}), .a ({new_AGEMA_signal_2635, KeyArray_outS22ser[0]}), .c ({new_AGEMA_signal_2636, KeyArray_inS21ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS21ser_mux_inst_1_U1 ( .s (KeyArray_n42), .b ({key_s1[49], key_s0[49]}), .a ({new_AGEMA_signal_2638, KeyArray_outS22ser[1]}), .c ({new_AGEMA_signal_2639, KeyArray_inS21ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS21ser_mux_inst_2_U1 ( .s (KeyArray_n42), .b ({key_s1[50], key_s0[50]}), .a ({new_AGEMA_signal_2641, KeyArray_outS22ser[2]}), .c ({new_AGEMA_signal_2642, KeyArray_inS21ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS21ser_mux_inst_3_U1 ( .s (KeyArray_n42), .b ({key_s1[51], key_s0[51]}), .a ({new_AGEMA_signal_2644, KeyArray_outS22ser[3]}), .c ({new_AGEMA_signal_2645, KeyArray_inS21ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS21ser_mux_inst_4_U1 ( .s (KeyArray_n42), .b ({key_s1[52], key_s0[52]}), .a ({new_AGEMA_signal_2647, KeyArray_outS22ser[4]}), .c ({new_AGEMA_signal_2648, KeyArray_inS21ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS21ser_mux_inst_5_U1 ( .s (KeyArray_n42), .b ({key_s1[53], key_s0[53]}), .a ({new_AGEMA_signal_2650, KeyArray_outS22ser[5]}), .c ({new_AGEMA_signal_2651, KeyArray_inS21ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS21ser_mux_inst_6_U1 ( .s (KeyArray_n42), .b ({key_s1[54], key_s0[54]}), .a ({new_AGEMA_signal_2653, KeyArray_outS22ser[6]}), .c ({new_AGEMA_signal_2654, KeyArray_inS21ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS21ser_mux_inst_7_U1 ( .s (KeyArray_n42), .b ({key_s1[55], key_s0[55]}), .a ({new_AGEMA_signal_2656, KeyArray_outS22ser[7]}), .c ({new_AGEMA_signal_2657, KeyArray_inS21ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS22ser_mux_inst_0_U1 ( .s (KeyArray_n41), .b ({key_s1[40], key_s0[40]}), .a ({new_AGEMA_signal_2659, KeyArray_outS23ser[0]}), .c ({new_AGEMA_signal_2660, KeyArray_inS22ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS22ser_mux_inst_1_U1 ( .s (KeyArray_n41), .b ({key_s1[41], key_s0[41]}), .a ({new_AGEMA_signal_2662, KeyArray_outS23ser[1]}), .c ({new_AGEMA_signal_2663, KeyArray_inS22ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS22ser_mux_inst_2_U1 ( .s (KeyArray_n41), .b ({key_s1[42], key_s0[42]}), .a ({new_AGEMA_signal_2665, KeyArray_outS23ser[2]}), .c ({new_AGEMA_signal_2666, KeyArray_inS22ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS22ser_mux_inst_3_U1 ( .s (KeyArray_n41), .b ({key_s1[43], key_s0[43]}), .a ({new_AGEMA_signal_2668, KeyArray_outS23ser[3]}), .c ({new_AGEMA_signal_2669, KeyArray_inS22ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS22ser_mux_inst_4_U1 ( .s (KeyArray_n41), .b ({key_s1[44], key_s0[44]}), .a ({new_AGEMA_signal_2671, KeyArray_outS23ser[4]}), .c ({new_AGEMA_signal_2672, KeyArray_inS22ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS22ser_mux_inst_5_U1 ( .s (KeyArray_n41), .b ({key_s1[45], key_s0[45]}), .a ({new_AGEMA_signal_2674, KeyArray_outS23ser[5]}), .c ({new_AGEMA_signal_2675, KeyArray_inS22ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS22ser_mux_inst_6_U1 ( .s (KeyArray_n41), .b ({key_s1[46], key_s0[46]}), .a ({new_AGEMA_signal_2677, KeyArray_outS23ser[6]}), .c ({new_AGEMA_signal_2678, KeyArray_inS22ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS22ser_mux_inst_7_U1 ( .s (KeyArray_n41), .b ({key_s1[47], key_s0[47]}), .a ({new_AGEMA_signal_2680, KeyArray_outS23ser[7]}), .c ({new_AGEMA_signal_2681, KeyArray_inS22ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS23ser_mux_inst_0_U1 ( .s (KeyArray_n41), .b ({key_s1[32], key_s0[32]}), .a ({new_AGEMA_signal_2683, KeyArray_outS30ser[0]}), .c ({new_AGEMA_signal_2684, KeyArray_inS23ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS23ser_mux_inst_1_U1 ( .s (KeyArray_n41), .b ({key_s1[33], key_s0[33]}), .a ({new_AGEMA_signal_2686, KeyArray_outS30ser[1]}), .c ({new_AGEMA_signal_2687, KeyArray_inS23ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS23ser_mux_inst_2_U1 ( .s (KeyArray_n41), .b ({key_s1[34], key_s0[34]}), .a ({new_AGEMA_signal_2689, KeyArray_outS30ser[2]}), .c ({new_AGEMA_signal_2690, KeyArray_inS23ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS23ser_mux_inst_3_U1 ( .s (KeyArray_n41), .b ({key_s1[35], key_s0[35]}), .a ({new_AGEMA_signal_2692, KeyArray_outS30ser[3]}), .c ({new_AGEMA_signal_2693, KeyArray_inS23ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS23ser_mux_inst_4_U1 ( .s (KeyArray_n41), .b ({key_s1[36], key_s0[36]}), .a ({new_AGEMA_signal_2695, KeyArray_outS30ser[4]}), .c ({new_AGEMA_signal_2696, KeyArray_inS23ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS23ser_mux_inst_5_U1 ( .s (KeyArray_n41), .b ({key_s1[37], key_s0[37]}), .a ({new_AGEMA_signal_2698, KeyArray_outS30ser[5]}), .c ({new_AGEMA_signal_2699, KeyArray_inS23ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS23ser_mux_inst_6_U1 ( .s (KeyArray_n41), .b ({key_s1[38], key_s0[38]}), .a ({new_AGEMA_signal_2701, KeyArray_outS30ser[6]}), .c ({new_AGEMA_signal_2702, KeyArray_inS23ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS23ser_mux_inst_7_U1 ( .s (KeyArray_n41), .b ({key_s1[39], key_s0[39]}), .a ({new_AGEMA_signal_2704, KeyArray_outS30ser[7]}), .c ({new_AGEMA_signal_2705, KeyArray_inS23ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS30ser_mux_inst_0_U1 ( .s (KeyArray_n40), .b ({key_s1[24], key_s0[24]}), .a ({new_AGEMA_signal_2707, KeyArray_outS31ser[0]}), .c ({new_AGEMA_signal_2708, KeyArray_inS30ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS30ser_mux_inst_1_U1 ( .s (KeyArray_n40), .b ({key_s1[25], key_s0[25]}), .a ({new_AGEMA_signal_2710, KeyArray_outS31ser[1]}), .c ({new_AGEMA_signal_2711, KeyArray_inS30ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS30ser_mux_inst_2_U1 ( .s (KeyArray_n40), .b ({key_s1[26], key_s0[26]}), .a ({new_AGEMA_signal_2713, KeyArray_outS31ser[2]}), .c ({new_AGEMA_signal_2714, KeyArray_inS30ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS30ser_mux_inst_3_U1 ( .s (KeyArray_n40), .b ({key_s1[27], key_s0[27]}), .a ({new_AGEMA_signal_2716, KeyArray_outS31ser[3]}), .c ({new_AGEMA_signal_2717, KeyArray_inS30ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS30ser_mux_inst_4_U1 ( .s (KeyArray_n40), .b ({key_s1[28], key_s0[28]}), .a ({new_AGEMA_signal_2719, KeyArray_outS31ser[4]}), .c ({new_AGEMA_signal_2720, KeyArray_inS30ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS30ser_mux_inst_5_U1 ( .s (KeyArray_n40), .b ({key_s1[29], key_s0[29]}), .a ({new_AGEMA_signal_2722, KeyArray_outS31ser[5]}), .c ({new_AGEMA_signal_2723, KeyArray_inS30ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS30ser_mux_inst_6_U1 ( .s (KeyArray_n40), .b ({key_s1[30], key_s0[30]}), .a ({new_AGEMA_signal_2725, KeyArray_outS31ser[6]}), .c ({new_AGEMA_signal_2726, KeyArray_inS30ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS30ser_mux_inst_7_U1 ( .s (KeyArray_n40), .b ({key_s1[31], key_s0[31]}), .a ({new_AGEMA_signal_2728, KeyArray_outS31ser[7]}), .c ({new_AGEMA_signal_2729, KeyArray_inS30ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS31ser_mux_inst_0_U1 ( .s (KeyArray_n40), .b ({key_s1[16], key_s0[16]}), .a ({new_AGEMA_signal_2731, KeyArray_outS32ser[0]}), .c ({new_AGEMA_signal_2732, KeyArray_inS31ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS31ser_mux_inst_1_U1 ( .s (KeyArray_n40), .b ({key_s1[17], key_s0[17]}), .a ({new_AGEMA_signal_2734, KeyArray_outS32ser[1]}), .c ({new_AGEMA_signal_2735, KeyArray_inS31ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS31ser_mux_inst_2_U1 ( .s (KeyArray_n40), .b ({key_s1[18], key_s0[18]}), .a ({new_AGEMA_signal_2737, KeyArray_outS32ser[2]}), .c ({new_AGEMA_signal_2738, KeyArray_inS31ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS31ser_mux_inst_3_U1 ( .s (KeyArray_n40), .b ({key_s1[19], key_s0[19]}), .a ({new_AGEMA_signal_2740, KeyArray_outS32ser[3]}), .c ({new_AGEMA_signal_2741, KeyArray_inS31ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS31ser_mux_inst_4_U1 ( .s (KeyArray_n40), .b ({key_s1[20], key_s0[20]}), .a ({new_AGEMA_signal_2743, KeyArray_outS32ser[4]}), .c ({new_AGEMA_signal_2744, KeyArray_inS31ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS31ser_mux_inst_5_U1 ( .s (KeyArray_n40), .b ({key_s1[21], key_s0[21]}), .a ({new_AGEMA_signal_2746, KeyArray_outS32ser[5]}), .c ({new_AGEMA_signal_2747, KeyArray_inS31ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS31ser_mux_inst_6_U1 ( .s (KeyArray_n40), .b ({key_s1[22], key_s0[22]}), .a ({new_AGEMA_signal_2749, KeyArray_outS32ser[6]}), .c ({new_AGEMA_signal_2750, KeyArray_inS31ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS31ser_mux_inst_7_U1 ( .s (KeyArray_n40), .b ({key_s1[23], key_s0[23]}), .a ({new_AGEMA_signal_2752, KeyArray_outS32ser[7]}), .c ({new_AGEMA_signal_2753, KeyArray_inS31ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS32ser_mux_inst_0_U1 ( .s (KeyArray_n39), .b ({key_s1[8], key_s0[8]}), .a ({new_AGEMA_signal_2755, KeyArray_outS33ser[0]}), .c ({new_AGEMA_signal_2756, KeyArray_inS32ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS32ser_mux_inst_1_U1 ( .s (KeyArray_n39), .b ({key_s1[9], key_s0[9]}), .a ({new_AGEMA_signal_2758, KeyArray_outS33ser[1]}), .c ({new_AGEMA_signal_2759, KeyArray_inS32ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS32ser_mux_inst_2_U1 ( .s (KeyArray_n39), .b ({key_s1[10], key_s0[10]}), .a ({new_AGEMA_signal_2761, KeyArray_outS33ser[2]}), .c ({new_AGEMA_signal_2762, KeyArray_inS32ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS32ser_mux_inst_3_U1 ( .s (KeyArray_n39), .b ({key_s1[11], key_s0[11]}), .a ({new_AGEMA_signal_2764, KeyArray_outS33ser[3]}), .c ({new_AGEMA_signal_2765, KeyArray_inS32ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS32ser_mux_inst_4_U1 ( .s (KeyArray_n39), .b ({key_s1[12], key_s0[12]}), .a ({new_AGEMA_signal_2767, KeyArray_outS33ser[4]}), .c ({new_AGEMA_signal_2768, KeyArray_inS32ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS32ser_mux_inst_5_U1 ( .s (KeyArray_n39), .b ({key_s1[13], key_s0[13]}), .a ({new_AGEMA_signal_2770, KeyArray_outS33ser[5]}), .c ({new_AGEMA_signal_2771, KeyArray_inS32ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS32ser_mux_inst_6_U1 ( .s (KeyArray_n39), .b ({key_s1[14], key_s0[14]}), .a ({new_AGEMA_signal_2773, KeyArray_outS33ser[6]}), .c ({new_AGEMA_signal_2774, KeyArray_inS32ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS32ser_mux_inst_7_U1 ( .s (KeyArray_n39), .b ({key_s1[15], key_s0[15]}), .a ({new_AGEMA_signal_2776, KeyArray_outS33ser[7]}), .c ({new_AGEMA_signal_2777, KeyArray_inS32ser[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS33ser_mux_inst_0_U1 ( .s (KeyArray_n39), .b ({key_s1[0], key_s0[0]}), .a ({new_AGEMA_signal_1983, keyStateIn[0]}), .c ({new_AGEMA_signal_2779, KeyArray_inS33ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS33ser_mux_inst_1_U1 ( .s (KeyArray_n39), .b ({key_s1[1], key_s0[1]}), .a ({new_AGEMA_signal_1986, keyStateIn[1]}), .c ({new_AGEMA_signal_2781, KeyArray_inS33ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS33ser_mux_inst_2_U1 ( .s (KeyArray_n39), .b ({key_s1[2], key_s0[2]}), .a ({new_AGEMA_signal_1989, keyStateIn[2]}), .c ({new_AGEMA_signal_2783, KeyArray_inS33ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS33ser_mux_inst_3_U1 ( .s (KeyArray_n39), .b ({key_s1[3], key_s0[3]}), .a ({new_AGEMA_signal_1992, keyStateIn[3]}), .c ({new_AGEMA_signal_2785, KeyArray_inS33ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS33ser_mux_inst_4_U1 ( .s (KeyArray_n39), .b ({key_s1[4], key_s0[4]}), .a ({new_AGEMA_signal_1995, keyStateIn[4]}), .c ({new_AGEMA_signal_2787, KeyArray_inS33ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS33ser_mux_inst_5_U1 ( .s (KeyArray_n39), .b ({key_s1[5], key_s0[5]}), .a ({new_AGEMA_signal_1998, keyStateIn[5]}), .c ({new_AGEMA_signal_2789, KeyArray_inS33ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS33ser_mux_inst_6_U1 ( .s (KeyArray_n39), .b ({key_s1[6], key_s0[6]}), .a ({new_AGEMA_signal_2001, keyStateIn[6]}), .c ({new_AGEMA_signal_2791, KeyArray_inS33ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_MUX_inS33ser_mux_inst_7_U1 ( .s (KeyArray_n39), .b ({key_s1[7], key_s0[7]}), .a ({new_AGEMA_signal_2004, keyStateIn[7]}), .c ({new_AGEMA_signal_2793, KeyArray_inS33ser[7]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U24 ( .a ({new_AGEMA_signal_2122, MixColumns_line0_n16}), .b ({new_AGEMA_signal_2024, MixColumns_line0_n15}), .c ({new_AGEMA_signal_2794, MCout[31]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U23 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({new_AGEMA_signal_2024, MixColumns_line0_n15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U22 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({new_AGEMA_signal_2051, MixColumns_line0_S13[7]}), .c ({new_AGEMA_signal_2122, MixColumns_line0_n16}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U21 ( .a ({new_AGEMA_signal_2123, MixColumns_line0_n14}), .b ({new_AGEMA_signal_2027, MixColumns_line0_n13}), .c ({new_AGEMA_signal_2795, MCout[30]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U20 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({new_AGEMA_signal_2027, MixColumns_line0_n13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U19 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({new_AGEMA_signal_2053, MixColumns_line0_S13[6]}), .c ({new_AGEMA_signal_2123, MixColumns_line0_n14}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U18 ( .a ({new_AGEMA_signal_2124, MixColumns_line0_n12}), .b ({new_AGEMA_signal_2030, MixColumns_line0_n11}), .c ({new_AGEMA_signal_2796, MCout[29]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U17 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_2030, MixColumns_line0_n11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U16 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_2055, MixColumns_line0_S13[5]}), .c ({new_AGEMA_signal_2124, MixColumns_line0_n12}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U15 ( .a ({new_AGEMA_signal_2797, MixColumns_line0_n10}), .b ({new_AGEMA_signal_2033, MixColumns_line0_n9}), .c ({new_AGEMA_signal_2838, MCout[28]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U14 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_2033, MixColumns_line0_n9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U13 ( .a ({new_AGEMA_signal_2046, MixColumns_line0_S02[4]}), .b ({new_AGEMA_signal_2127, MixColumns_line0_S13[4]}), .c ({new_AGEMA_signal_2797, MixColumns_line0_n10}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U12 ( .a ({new_AGEMA_signal_2798, MixColumns_line0_n8}), .b ({new_AGEMA_signal_2036, MixColumns_line0_n7}), .c ({new_AGEMA_signal_2839, MCout[27]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U11 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_2036, MixColumns_line0_n7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U10 ( .a ({new_AGEMA_signal_2047, MixColumns_line0_S02[3]}), .b ({new_AGEMA_signal_2128, MixColumns_line0_S13[3]}), .c ({new_AGEMA_signal_2798, MixColumns_line0_n8}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U9 ( .a ({new_AGEMA_signal_2125, MixColumns_line0_n6}), .b ({new_AGEMA_signal_2039, MixColumns_line0_n5}), .c ({new_AGEMA_signal_2799, MCout[26]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U8 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_2039, MixColumns_line0_n5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U7 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_2058, MixColumns_line0_S13[2]}), .c ({new_AGEMA_signal_2125, MixColumns_line0_n6}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U6 ( .a ({new_AGEMA_signal_2800, MixColumns_line0_n4}), .b ({new_AGEMA_signal_2042, MixColumns_line0_n3}), .c ({new_AGEMA_signal_2840, MCout[25]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U5 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_2042, MixColumns_line0_n3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U4 ( .a ({new_AGEMA_signal_2048, MixColumns_line0_S02[1]}), .b ({new_AGEMA_signal_2129, MixColumns_line0_S13[1]}), .c ({new_AGEMA_signal_2800, MixColumns_line0_n4}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U3 ( .a ({new_AGEMA_signal_2126, MixColumns_line0_n2}), .b ({new_AGEMA_signal_2045, MixColumns_line0_n1}), .c ({new_AGEMA_signal_2801, MCout[24]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U2 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_2045, MixColumns_line0_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_U1 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2060, MixColumns_line0_S13[0]}), .c ({new_AGEMA_signal_2126, MixColumns_line0_n2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_timesTWO_U3 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_2046, MixColumns_line0_S02[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_timesTWO_U2 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_2047, MixColumns_line0_S02[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_timesTWO_U1 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_2048, MixColumns_line0_S02[1]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_timesTHREE_U8 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({new_AGEMA_signal_2051, MixColumns_line0_S13[7]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_timesTHREE_U7 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_2053, MixColumns_line0_S13[6]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_timesTHREE_U6 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_2055, MixColumns_line0_S13[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_timesTHREE_U5 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({new_AGEMA_signal_2062, MixColumns_line0_timesTHREE_input2[4]}), .c ({new_AGEMA_signal_2127, MixColumns_line0_S13[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_timesTHREE_U4 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({new_AGEMA_signal_2063, MixColumns_line0_timesTHREE_input2[3]}), .c ({new_AGEMA_signal_2128, MixColumns_line0_S13[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_timesTHREE_U3 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_2058, MixColumns_line0_S13[2]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_timesTHREE_U2 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({new_AGEMA_signal_2064, MixColumns_line0_timesTHREE_input2[1]}), .c ({new_AGEMA_signal_2129, MixColumns_line0_S13[1]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_timesTHREE_U1 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({new_AGEMA_signal_2060, MixColumns_line0_S13[0]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_timesTHREE_timesTWO_U3 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_2062, MixColumns_line0_timesTHREE_input2[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_timesTHREE_timesTWO_U2 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_2063, MixColumns_line0_timesTHREE_input2[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line0_timesTHREE_timesTWO_U1 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_2064, MixColumns_line0_timesTHREE_input2[1]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U24 ( .a ({new_AGEMA_signal_2130, MixColumns_line1_n16}), .b ({new_AGEMA_signal_2065, MixColumns_line1_n15}), .c ({new_AGEMA_signal_2802, MCout[23]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U23 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({new_AGEMA_signal_2065, MixColumns_line1_n15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U22 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({new_AGEMA_signal_2076, MixColumns_line1_S13[7]}), .c ({new_AGEMA_signal_2130, MixColumns_line1_n16}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U21 ( .a ({new_AGEMA_signal_2131, MixColumns_line1_n14}), .b ({new_AGEMA_signal_2066, MixColumns_line1_n13}), .c ({new_AGEMA_signal_2803, MCout[22]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U20 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({new_AGEMA_signal_2066, MixColumns_line1_n13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U19 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({new_AGEMA_signal_2077, MixColumns_line1_S13[6]}), .c ({new_AGEMA_signal_2131, MixColumns_line1_n14}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U18 ( .a ({new_AGEMA_signal_2132, MixColumns_line1_n12}), .b ({new_AGEMA_signal_2067, MixColumns_line1_n11}), .c ({new_AGEMA_signal_2804, MCout[21]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U17 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_2067, MixColumns_line1_n11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U16 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({new_AGEMA_signal_2078, MixColumns_line1_S13[5]}), .c ({new_AGEMA_signal_2132, MixColumns_line1_n12}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U15 ( .a ({new_AGEMA_signal_2805, MixColumns_line1_n10}), .b ({new_AGEMA_signal_2068, MixColumns_line1_n9}), .c ({new_AGEMA_signal_2841, MCout[20]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U14 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_2068, MixColumns_line1_n9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U13 ( .a ({new_AGEMA_signal_2073, MixColumns_line1_S02_4_}), .b ({new_AGEMA_signal_2135, MixColumns_line1_S13[4]}), .c ({new_AGEMA_signal_2805, MixColumns_line1_n10}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U12 ( .a ({new_AGEMA_signal_2806, MixColumns_line1_n8}), .b ({new_AGEMA_signal_2069, MixColumns_line1_n7}), .c ({new_AGEMA_signal_2842, MCout[19]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U11 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_2069, MixColumns_line1_n7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U10 ( .a ({new_AGEMA_signal_2074, MixColumns_line1_S02_3_}), .b ({new_AGEMA_signal_2136, MixColumns_line1_S13[3]}), .c ({new_AGEMA_signal_2806, MixColumns_line1_n8}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U9 ( .a ({new_AGEMA_signal_2133, MixColumns_line1_n6}), .b ({new_AGEMA_signal_2070, MixColumns_line1_n5}), .c ({new_AGEMA_signal_2807, MCout[18]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U8 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_2070, MixColumns_line1_n5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U7 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({new_AGEMA_signal_2079, MixColumns_line1_S13[2]}), .c ({new_AGEMA_signal_2133, MixColumns_line1_n6}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U6 ( .a ({new_AGEMA_signal_2808, MixColumns_line1_n4}), .b ({new_AGEMA_signal_2071, MixColumns_line1_n3}), .c ({new_AGEMA_signal_2843, MCout[17]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U5 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_2071, MixColumns_line1_n3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U4 ( .a ({new_AGEMA_signal_2075, MixColumns_line1_S02_1_}), .b ({new_AGEMA_signal_2137, MixColumns_line1_S13[1]}), .c ({new_AGEMA_signal_2808, MixColumns_line1_n4}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U3 ( .a ({new_AGEMA_signal_2134, MixColumns_line1_n2}), .b ({new_AGEMA_signal_2072, MixColumns_line1_n1}), .c ({new_AGEMA_signal_2809, MCout[16]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U2 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_2072, MixColumns_line1_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_U1 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_2080, MixColumns_line1_S13[0]}), .c ({new_AGEMA_signal_2134, MixColumns_line1_n2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_timesTWO_U3 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_2073, MixColumns_line1_S02_4_}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_timesTWO_U2 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_2074, MixColumns_line1_S02_3_}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_timesTWO_U1 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_2075, MixColumns_line1_S02_1_}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_timesTHREE_U8 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({new_AGEMA_signal_2076, MixColumns_line1_S13[7]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_timesTHREE_U7 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_2077, MixColumns_line1_S13[6]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_timesTHREE_U6 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_2078, MixColumns_line1_S13[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_timesTHREE_U5 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_2081, MixColumns_line1_timesTHREE_input2[4]}), .c ({new_AGEMA_signal_2135, MixColumns_line1_S13[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_timesTHREE_U4 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_2082, MixColumns_line1_timesTHREE_input2[3]}), .c ({new_AGEMA_signal_2136, MixColumns_line1_S13[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_timesTHREE_U3 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_2079, MixColumns_line1_S13[2]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_timesTHREE_U2 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_2083, MixColumns_line1_timesTHREE_input2[1]}), .c ({new_AGEMA_signal_2137, MixColumns_line1_S13[1]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_timesTHREE_U1 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({new_AGEMA_signal_2080, MixColumns_line1_S13[0]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_timesTHREE_timesTWO_U3 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_2081, MixColumns_line1_timesTHREE_input2[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_timesTHREE_timesTWO_U2 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_2082, MixColumns_line1_timesTHREE_input2[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line1_timesTHREE_timesTWO_U1 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_2083, MixColumns_line1_timesTHREE_input2[1]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U24 ( .a ({new_AGEMA_signal_2138, MixColumns_line2_n16}), .b ({new_AGEMA_signal_2084, MixColumns_line2_n15}), .c ({new_AGEMA_signal_2810, MCout[15]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U23 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({new_AGEMA_signal_2084, MixColumns_line2_n15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U22 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_2095, MixColumns_line2_S13[7]}), .c ({new_AGEMA_signal_2138, MixColumns_line2_n16}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U21 ( .a ({new_AGEMA_signal_2139, MixColumns_line2_n14}), .b ({new_AGEMA_signal_2085, MixColumns_line2_n13}), .c ({new_AGEMA_signal_2811, MCout[14]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U20 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({new_AGEMA_signal_2085, MixColumns_line2_n13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U19 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({new_AGEMA_signal_2096, MixColumns_line2_S13[6]}), .c ({new_AGEMA_signal_2139, MixColumns_line2_n14}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U18 ( .a ({new_AGEMA_signal_2140, MixColumns_line2_n12}), .b ({new_AGEMA_signal_2086, MixColumns_line2_n11}), .c ({new_AGEMA_signal_2812, MCout[13]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U17 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_2086, MixColumns_line2_n11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U16 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_2097, MixColumns_line2_S13[5]}), .c ({new_AGEMA_signal_2140, MixColumns_line2_n12}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U15 ( .a ({new_AGEMA_signal_2813, MixColumns_line2_n10}), .b ({new_AGEMA_signal_2087, MixColumns_line2_n9}), .c ({new_AGEMA_signal_2844, MCout[12]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U14 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_2087, MixColumns_line2_n9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U13 ( .a ({new_AGEMA_signal_2092, MixColumns_line2_S02_4_}), .b ({new_AGEMA_signal_2143, MixColumns_line2_S13[4]}), .c ({new_AGEMA_signal_2813, MixColumns_line2_n10}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U12 ( .a ({new_AGEMA_signal_2814, MixColumns_line2_n8}), .b ({new_AGEMA_signal_2088, MixColumns_line2_n7}), .c ({new_AGEMA_signal_2845, MCout[11]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U11 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_2088, MixColumns_line2_n7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U10 ( .a ({new_AGEMA_signal_2093, MixColumns_line2_S02_3_}), .b ({new_AGEMA_signal_2144, MixColumns_line2_S13[3]}), .c ({new_AGEMA_signal_2814, MixColumns_line2_n8}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U9 ( .a ({new_AGEMA_signal_2141, MixColumns_line2_n6}), .b ({new_AGEMA_signal_2089, MixColumns_line2_n5}), .c ({new_AGEMA_signal_2815, MCout[10]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U8 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_2089, MixColumns_line2_n5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U7 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_2098, MixColumns_line2_S13[2]}), .c ({new_AGEMA_signal_2141, MixColumns_line2_n6}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U6 ( .a ({new_AGEMA_signal_2816, MixColumns_line2_n4}), .b ({new_AGEMA_signal_2090, MixColumns_line2_n3}), .c ({new_AGEMA_signal_2846, MCout[9]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U5 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_2090, MixColumns_line2_n3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U4 ( .a ({new_AGEMA_signal_2094, MixColumns_line2_S02_1_}), .b ({new_AGEMA_signal_2145, MixColumns_line2_S13[1]}), .c ({new_AGEMA_signal_2816, MixColumns_line2_n4}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U3 ( .a ({new_AGEMA_signal_2142, MixColumns_line2_n2}), .b ({new_AGEMA_signal_2091, MixColumns_line2_n1}), .c ({new_AGEMA_signal_2817, MCout[8]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U2 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_2091, MixColumns_line2_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_U1 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_2099, MixColumns_line2_S13[0]}), .c ({new_AGEMA_signal_2142, MixColumns_line2_n2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_timesTWO_U3 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_2092, MixColumns_line2_S02_4_}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_timesTWO_U2 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_2093, MixColumns_line2_S02_3_}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_timesTWO_U1 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_2094, MixColumns_line2_S02_1_}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_timesTHREE_U8 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({new_AGEMA_signal_2095, MixColumns_line2_S13[7]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_timesTHREE_U7 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_2096, MixColumns_line2_S13[6]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_timesTHREE_U6 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_2097, MixColumns_line2_S13[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_timesTHREE_U5 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_2100, MixColumns_line2_timesTHREE_input2[4]}), .c ({new_AGEMA_signal_2143, MixColumns_line2_S13[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_timesTHREE_U4 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_2101, MixColumns_line2_timesTHREE_input2[3]}), .c ({new_AGEMA_signal_2144, MixColumns_line2_S13[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_timesTHREE_U3 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_2098, MixColumns_line2_S13[2]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_timesTHREE_U2 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_2102, MixColumns_line2_timesTHREE_input2[1]}), .c ({new_AGEMA_signal_2145, MixColumns_line2_S13[1]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_timesTHREE_U1 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({new_AGEMA_signal_2099, MixColumns_line2_S13[0]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_timesTHREE_timesTWO_U3 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_2100, MixColumns_line2_timesTHREE_input2[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_timesTHREE_timesTWO_U2 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_2101, MixColumns_line2_timesTHREE_input2[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line2_timesTHREE_timesTWO_U1 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_2102, MixColumns_line2_timesTHREE_input2[1]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U24 ( .a ({new_AGEMA_signal_2146, MixColumns_line3_n16}), .b ({new_AGEMA_signal_2103, MixColumns_line3_n15}), .c ({new_AGEMA_signal_2818, MCout[7]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U23 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({new_AGEMA_signal_2103, MixColumns_line3_n15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U22 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_2114, MixColumns_line3_S13[7]}), .c ({new_AGEMA_signal_2146, MixColumns_line3_n16}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U21 ( .a ({new_AGEMA_signal_2147, MixColumns_line3_n14}), .b ({new_AGEMA_signal_2104, MixColumns_line3_n13}), .c ({new_AGEMA_signal_2819, MCout[6]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U20 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({new_AGEMA_signal_2104, MixColumns_line3_n13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U19 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({new_AGEMA_signal_2115, MixColumns_line3_S13[6]}), .c ({new_AGEMA_signal_2147, MixColumns_line3_n14}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U18 ( .a ({new_AGEMA_signal_2148, MixColumns_line3_n12}), .b ({new_AGEMA_signal_2105, MixColumns_line3_n11}), .c ({new_AGEMA_signal_2820, MCout[5]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U17 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_2105, MixColumns_line3_n11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U16 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_2116, MixColumns_line3_S13[5]}), .c ({new_AGEMA_signal_2148, MixColumns_line3_n12}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U15 ( .a ({new_AGEMA_signal_2821, MixColumns_line3_n10}), .b ({new_AGEMA_signal_2106, MixColumns_line3_n9}), .c ({new_AGEMA_signal_2847, MCout[4]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U14 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_2106, MixColumns_line3_n9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U13 ( .a ({new_AGEMA_signal_2111, MixColumns_line3_S02_4_}), .b ({new_AGEMA_signal_2151, MixColumns_line3_S13[4]}), .c ({new_AGEMA_signal_2821, MixColumns_line3_n10}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U12 ( .a ({new_AGEMA_signal_2822, MixColumns_line3_n8}), .b ({new_AGEMA_signal_2107, MixColumns_line3_n7}), .c ({new_AGEMA_signal_2848, MCout[3]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U11 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_2107, MixColumns_line3_n7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U10 ( .a ({new_AGEMA_signal_2112, MixColumns_line3_S02_3_}), .b ({new_AGEMA_signal_2152, MixColumns_line3_S13[3]}), .c ({new_AGEMA_signal_2822, MixColumns_line3_n8}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U9 ( .a ({new_AGEMA_signal_2149, MixColumns_line3_n6}), .b ({new_AGEMA_signal_2108, MixColumns_line3_n5}), .c ({new_AGEMA_signal_2823, MCout[2]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U8 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_2108, MixColumns_line3_n5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U7 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_2117, MixColumns_line3_S13[2]}), .c ({new_AGEMA_signal_2149, MixColumns_line3_n6}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U6 ( .a ({new_AGEMA_signal_2824, MixColumns_line3_n4}), .b ({new_AGEMA_signal_2109, MixColumns_line3_n3}), .c ({new_AGEMA_signal_2849, MCout[1]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U5 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_2109, MixColumns_line3_n3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U4 ( .a ({new_AGEMA_signal_2113, MixColumns_line3_S02_1_}), .b ({new_AGEMA_signal_2153, MixColumns_line3_S13[1]}), .c ({new_AGEMA_signal_2824, MixColumns_line3_n4}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U3 ( .a ({new_AGEMA_signal_2150, MixColumns_line3_n2}), .b ({new_AGEMA_signal_2110, MixColumns_line3_n1}), .c ({new_AGEMA_signal_2825, MCout[0]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U2 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_2110, MixColumns_line3_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_U1 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2118, MixColumns_line3_S13[0]}), .c ({new_AGEMA_signal_2150, MixColumns_line3_n2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_timesTWO_U3 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_2111, MixColumns_line3_S02_4_}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_timesTWO_U2 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_2112, MixColumns_line3_S02_3_}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_timesTWO_U1 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_2113, MixColumns_line3_S02_1_}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_timesTHREE_U8 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({new_AGEMA_signal_2114, MixColumns_line3_S13[7]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_timesTHREE_U7 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_2115, MixColumns_line3_S13[6]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_timesTHREE_U6 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_2116, MixColumns_line3_S13[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_timesTHREE_U5 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_2119, MixColumns_line3_timesTHREE_input2_4_}), .c ({new_AGEMA_signal_2151, MixColumns_line3_S13[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_timesTHREE_U4 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({new_AGEMA_signal_2120, MixColumns_line3_timesTHREE_input2_3_}), .c ({new_AGEMA_signal_2152, MixColumns_line3_S13[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_timesTHREE_U3 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_2117, MixColumns_line3_S13[2]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_timesTHREE_U2 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_2121, MixColumns_line3_timesTHREE_input2_1_}), .c ({new_AGEMA_signal_2153, MixColumns_line3_S13[1]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_timesTHREE_U1 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({new_AGEMA_signal_2118, MixColumns_line3_S13[0]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_timesTHREE_timesTWO_U3 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_2119, MixColumns_line3_timesTHREE_input2_4_}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_timesTHREE_timesTWO_U2 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_2120, MixColumns_line3_timesTHREE_input2_3_}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) MixColumns_line3_timesTHREE_timesTWO_U1 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_2121, MixColumns_line3_timesTHREE_input2_1_}) ) ;
    NOR2_X1 calcRCon_U46 ( .A1 (calcRCon_n11), .A2 (calcRCon_n38), .ZN (roundConstant[7]) ) ;
    NOR2_X1 calcRCon_U45 ( .A1 (calcRCon_n16), .A2 (calcRCon_n38), .ZN (roundConstant[6]) ) ;
    AND2_X1 calcRCon_U44 ( .A1 (calcRCon_s_current_state_5_), .A2 (enRCon), .ZN (roundConstant[5]) ) ;
    AND2_X1 calcRCon_U43 ( .A1 (calcRCon_s_current_state_4_), .A2 (enRCon), .ZN (roundConstant[4]) ) ;
    NOR2_X1 calcRCon_U42 ( .A1 (calcRCon_n15), .A2 (calcRCon_n38), .ZN (roundConstant[3]) ) ;
    NOR2_X1 calcRCon_U41 ( .A1 (calcRCon_n12), .A2 (calcRCon_n38), .ZN (roundConstant[2]) ) ;
    NOR2_X1 calcRCon_U40 ( .A1 (calcRCon_n14), .A2 (calcRCon_n38), .ZN (roundConstant[1]) ) ;
    NOR2_X1 calcRCon_U39 ( .A1 (calcRCon_n13), .A2 (calcRCon_n38), .ZN (roundConstant[0]) ) ;
    INV_X1 calcRCon_U38 ( .A (enRCon), .ZN (calcRCon_n38) ) ;
    NAND2_X1 calcRCon_U37 ( .A1 (calcRCon_n37), .A2 (calcRCon_n36), .ZN (notFirst) ) ;
    NOR2_X1 calcRCon_U36 ( .A1 (calcRCon_n35), .A2 (calcRCon_n34), .ZN (calcRCon_n36) ) ;
    NAND2_X1 calcRCon_U35 ( .A1 (calcRCon_n33), .A2 (calcRCon_n32), .ZN (calcRCon_n34) ) ;
    NOR2_X1 calcRCon_U34 ( .A1 (calcRCon_s_current_state_1_), .A2 (calcRCon_n15), .ZN (calcRCon_n32) ) ;
    NOR2_X1 calcRCon_U33 ( .A1 (calcRCon_s_current_state_6_), .A2 (calcRCon_n13), .ZN (calcRCon_n33) ) ;
    NAND2_X1 calcRCon_U32 ( .A1 (calcRCon_s_current_state_2_), .A2 (calcRCon_n3), .ZN (calcRCon_n35) ) ;
    NOR2_X1 calcRCon_U31 ( .A1 (calcRCon_s_current_state_4_), .A2 (calcRCon_s_current_state_5_), .ZN (calcRCon_n37) ) ;
    NAND2_X1 calcRCon_U30 ( .A1 (nReset), .A2 (calcRCon_n31), .ZN (calcRCon_n51) ) ;
    MUX2_X1 calcRCon_U29 ( .S (calcRCon_n5), .A (calcRCon_n11), .B (calcRCon_n13), .Z (calcRCon_n31) ) ;
    NAND2_X1 calcRCon_U28 ( .A1 (calcRCon_n30), .A2 (calcRCon_n29), .ZN (calcRCon_n50) ) ;
    NAND2_X1 calcRCon_U27 ( .A1 (calcRCon_n28), .A2 (calcRCon_s_current_state_1_), .ZN (calcRCon_n29) ) ;
    NAND2_X1 calcRCon_U26 ( .A1 (calcRCon_n27), .A2 (calcRCon_n26), .ZN (calcRCon_n30) ) ;
    XOR2_X1 calcRCon_U25 ( .A (calcRCon_s_current_state_0_), .B (calcRCon_n3), .Z (calcRCon_n27) ) ;
    NAND2_X1 calcRCon_U24 ( .A1 (nReset), .A2 (calcRCon_n25), .ZN (calcRCon_n49) ) ;
    MUX2_X1 calcRCon_U23 ( .S (calcRCon_n5), .A (calcRCon_n14), .B (calcRCon_n12), .Z (calcRCon_n25) ) ;
    NAND2_X1 calcRCon_U22 ( .A1 (nReset), .A2 (calcRCon_n24), .ZN (calcRCon_n48) ) ;
    MUX2_X1 calcRCon_U21 ( .S (calcRCon_n5), .A (calcRCon_n23), .B (calcRCon_n15), .Z (calcRCon_n24) ) ;
    XNOR2_X1 calcRCon_U20 ( .A (calcRCon_n3), .B (calcRCon_s_current_state_2_), .ZN (calcRCon_n23) ) ;
    NAND2_X1 calcRCon_U19 ( .A1 (calcRCon_n22), .A2 (calcRCon_n21), .ZN (calcRCon_n47) ) ;
    NAND2_X1 calcRCon_U18 ( .A1 (calcRCon_s_current_state_4_), .A2 (calcRCon_n28), .ZN (calcRCon_n21) ) ;
    NAND2_X1 calcRCon_U17 ( .A1 (calcRCon_n20), .A2 (calcRCon_n26), .ZN (calcRCon_n22) ) ;
    XOR2_X1 calcRCon_U16 ( .A (calcRCon_n15), .B (calcRCon_n11), .Z (calcRCon_n20) ) ;
    NAND2_X1 calcRCon_U15 ( .A1 (calcRCon_n19), .A2 (calcRCon_n18), .ZN (calcRCon_n46) ) ;
    NAND2_X1 calcRCon_U14 ( .A1 (calcRCon_s_current_state_4_), .A2 (calcRCon_n26), .ZN (calcRCon_n18) ) ;
    NAND2_X1 calcRCon_U13 ( .A1 (calcRCon_s_current_state_5_), .A2 (calcRCon_n28), .ZN (calcRCon_n19) ) ;
    NAND2_X1 calcRCon_U12 ( .A1 (calcRCon_n17), .A2 (calcRCon_n10), .ZN (calcRCon_n45) ) ;
    NAND2_X1 calcRCon_U11 ( .A1 (calcRCon_s_current_state_5_), .A2 (calcRCon_n26), .ZN (calcRCon_n10) ) ;
    NOR2_X1 calcRCon_U10 ( .A1 (calcRCon_n5), .A2 (calcRCon_n6), .ZN (calcRCon_n26) ) ;
    NAND2_X1 calcRCon_U9 ( .A1 (calcRCon_s_current_state_6_), .A2 (calcRCon_n28), .ZN (calcRCon_n17) ) ;
    NOR2_X1 calcRCon_U8 ( .A1 (selSR), .A2 (calcRCon_n6), .ZN (calcRCon_n28) ) ;
    NAND2_X1 calcRCon_U7 ( .A1 (nReset), .A2 (calcRCon_n9), .ZN (calcRCon_n44) ) ;
    MUX2_X1 calcRCon_U6 ( .S (calcRCon_n5), .A (calcRCon_n16), .B (calcRCon_n11), .Z (calcRCon_n9) ) ;
    NAND2_X1 calcRCon_U5 ( .A1 (calcRCon_s_current_state_4_), .A2 (calcRCon_s_current_state_2_), .ZN (calcRCon_n7) ) ;
    NAND2_X1 calcRCon_U4 ( .A1 (calcRCon_s_current_state_1_), .A2 (calcRCon_s_current_state_5_), .ZN (calcRCon_n8) ) ;
    INV_X1 calcRCon_U3 ( .A (nReset), .ZN (calcRCon_n6) ) ;
    INV_X1 calcRCon_U2 ( .A (selSR), .ZN (calcRCon_n5) ) ;
    NOR2_X1 calcRCon_U1 ( .A1 (calcRCon_n8), .A2 (calcRCon_n7), .ZN (intFinal) ) ;
    INV_X1 calcRCon_s_current_state_reg_0__U1 ( .A (calcRCon_s_current_state_0_), .ZN (calcRCon_n13) ) ;
    INV_X1 calcRCon_s_current_state_reg_1__U1 ( .A (calcRCon_s_current_state_1_), .ZN (calcRCon_n14) ) ;
    INV_X1 calcRCon_s_current_state_reg_2__U1 ( .A (calcRCon_s_current_state_2_), .ZN (calcRCon_n12) ) ;
    INV_X1 calcRCon_s_current_state_reg_3__U1 ( .A (calcRCon_s_current_state_3_), .ZN (calcRCon_n15) ) ;
    INV_X1 calcRCon_s_current_state_reg_6__U1 ( .A (calcRCon_s_current_state_6_), .ZN (calcRCon_n16) ) ;
    INV_X1 calcRCon_s_current_state_reg_7__U1 ( .A (calcRCon_n3), .ZN (calcRCon_n11) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_SboxIn_mux_inst_0_U1 ( .s (selMC), .b ({new_AGEMA_signal_1984, StateOutXORroundKey[0]}), .a ({new_AGEMA_signal_2563, keySBIn[0]}), .c ({new_AGEMA_signal_2826, SboxIn[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_SboxIn_mux_inst_1_U1 ( .s (selMC), .b ({new_AGEMA_signal_1987, StateOutXORroundKey[1]}), .a ({new_AGEMA_signal_2566, keySBIn[1]}), .c ({new_AGEMA_signal_2827, SboxIn[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_SboxIn_mux_inst_2_U1 ( .s (selMC), .b ({new_AGEMA_signal_1990, StateOutXORroundKey[2]}), .a ({new_AGEMA_signal_2569, keySBIn[2]}), .c ({new_AGEMA_signal_2828, SboxIn[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_SboxIn_mux_inst_3_U1 ( .s (selMC), .b ({new_AGEMA_signal_1993, StateOutXORroundKey[3]}), .a ({new_AGEMA_signal_2572, keySBIn[3]}), .c ({new_AGEMA_signal_2829, SboxIn[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_SboxIn_mux_inst_4_U1 ( .s (selMC), .b ({new_AGEMA_signal_1996, StateOutXORroundKey[4]}), .a ({new_AGEMA_signal_2575, keySBIn[4]}), .c ({new_AGEMA_signal_2830, SboxIn[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_SboxIn_mux_inst_5_U1 ( .s (selMC), .b ({new_AGEMA_signal_1999, StateOutXORroundKey[5]}), .a ({new_AGEMA_signal_2578, keySBIn[5]}), .c ({new_AGEMA_signal_2831, SboxIn[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_SboxIn_mux_inst_6_U1 ( .s (selMC), .b ({new_AGEMA_signal_2002, StateOutXORroundKey[6]}), .a ({new_AGEMA_signal_2581, keySBIn[6]}), .c ({new_AGEMA_signal_2832, SboxIn[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_SboxIn_mux_inst_7_U1 ( .s (selMC), .b ({new_AGEMA_signal_2005, StateOutXORroundKey[7]}), .a ({new_AGEMA_signal_2584, keySBIn[7]}), .c ({new_AGEMA_signal_2833, SboxIn[7]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T1_U1 ( .a ({new_AGEMA_signal_2833, SboxIn[7]}), .b ({new_AGEMA_signal_2830, SboxIn[4]}), .c ({new_AGEMA_signal_2850, Inst_bSbox_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T2_U1 ( .a ({new_AGEMA_signal_2833, SboxIn[7]}), .b ({new_AGEMA_signal_2828, SboxIn[2]}), .c ({new_AGEMA_signal_2851, Inst_bSbox_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T3_U1 ( .a ({new_AGEMA_signal_2833, SboxIn[7]}), .b ({new_AGEMA_signal_2827, SboxIn[1]}), .c ({new_AGEMA_signal_2852, Inst_bSbox_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T4_U1 ( .a ({new_AGEMA_signal_2830, SboxIn[4]}), .b ({new_AGEMA_signal_2828, SboxIn[2]}), .c ({new_AGEMA_signal_2853, Inst_bSbox_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T5_U1 ( .a ({new_AGEMA_signal_2829, SboxIn[3]}), .b ({new_AGEMA_signal_2827, SboxIn[1]}), .c ({new_AGEMA_signal_2854, Inst_bSbox_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T6_U1 ( .a ({new_AGEMA_signal_2850, Inst_bSbox_T1}), .b ({new_AGEMA_signal_2854, Inst_bSbox_T5}), .c ({new_AGEMA_signal_3000, Inst_bSbox_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T7_U1 ( .a ({new_AGEMA_signal_2832, SboxIn[6]}), .b ({new_AGEMA_signal_2831, SboxIn[5]}), .c ({new_AGEMA_signal_2855, Inst_bSbox_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T8_U1 ( .a ({new_AGEMA_signal_2826, SboxIn[0]}), .b ({new_AGEMA_signal_3000, Inst_bSbox_T6}), .c ({new_AGEMA_signal_3032, Inst_bSbox_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T9_U1 ( .a ({new_AGEMA_signal_2826, SboxIn[0]}), .b ({new_AGEMA_signal_2855, Inst_bSbox_T7}), .c ({new_AGEMA_signal_3001, Inst_bSbox_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T10_U1 ( .a ({new_AGEMA_signal_3000, Inst_bSbox_T6}), .b ({new_AGEMA_signal_2855, Inst_bSbox_T7}), .c ({new_AGEMA_signal_3033, Inst_bSbox_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T11_U1 ( .a ({new_AGEMA_signal_2832, SboxIn[6]}), .b ({new_AGEMA_signal_2828, SboxIn[2]}), .c ({new_AGEMA_signal_2856, Inst_bSbox_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T12_U1 ( .a ({new_AGEMA_signal_2831, SboxIn[5]}), .b ({new_AGEMA_signal_2828, SboxIn[2]}), .c ({new_AGEMA_signal_2857, Inst_bSbox_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T13_U1 ( .a ({new_AGEMA_signal_2852, Inst_bSbox_T3}), .b ({new_AGEMA_signal_2853, Inst_bSbox_T4}), .c ({new_AGEMA_signal_3002, Inst_bSbox_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T14_U1 ( .a ({new_AGEMA_signal_3000, Inst_bSbox_T6}), .b ({new_AGEMA_signal_2856, Inst_bSbox_T11}), .c ({new_AGEMA_signal_3034, Inst_bSbox_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T15_U1 ( .a ({new_AGEMA_signal_2854, Inst_bSbox_T5}), .b ({new_AGEMA_signal_2856, Inst_bSbox_T11}), .c ({new_AGEMA_signal_3003, Inst_bSbox_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T16_U1 ( .a ({new_AGEMA_signal_2854, Inst_bSbox_T5}), .b ({new_AGEMA_signal_2857, Inst_bSbox_T12}), .c ({new_AGEMA_signal_3004, Inst_bSbox_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T17_U1 ( .a ({new_AGEMA_signal_3001, Inst_bSbox_T9}), .b ({new_AGEMA_signal_3004, Inst_bSbox_T16}), .c ({new_AGEMA_signal_3035, Inst_bSbox_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T18_U1 ( .a ({new_AGEMA_signal_2830, SboxIn[4]}), .b ({new_AGEMA_signal_2826, SboxIn[0]}), .c ({new_AGEMA_signal_2858, Inst_bSbox_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T19_U1 ( .a ({new_AGEMA_signal_2855, Inst_bSbox_T7}), .b ({new_AGEMA_signal_2858, Inst_bSbox_T18}), .c ({new_AGEMA_signal_3005, Inst_bSbox_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T20_U1 ( .a ({new_AGEMA_signal_2850, Inst_bSbox_T1}), .b ({new_AGEMA_signal_3005, Inst_bSbox_T19}), .c ({new_AGEMA_signal_3036, Inst_bSbox_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T21_U1 ( .a ({new_AGEMA_signal_2827, SboxIn[1]}), .b ({new_AGEMA_signal_2826, SboxIn[0]}), .c ({new_AGEMA_signal_2859, Inst_bSbox_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T22_U1 ( .a ({new_AGEMA_signal_2855, Inst_bSbox_T7}), .b ({new_AGEMA_signal_2859, Inst_bSbox_T21}), .c ({new_AGEMA_signal_3006, Inst_bSbox_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T23_U1 ( .a ({new_AGEMA_signal_2851, Inst_bSbox_T2}), .b ({new_AGEMA_signal_3006, Inst_bSbox_T22}), .c ({new_AGEMA_signal_3037, Inst_bSbox_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T24_U1 ( .a ({new_AGEMA_signal_2851, Inst_bSbox_T2}), .b ({new_AGEMA_signal_3033, Inst_bSbox_T10}), .c ({new_AGEMA_signal_3117, Inst_bSbox_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T25_U1 ( .a ({new_AGEMA_signal_3036, Inst_bSbox_T20}), .b ({new_AGEMA_signal_3035, Inst_bSbox_T17}), .c ({new_AGEMA_signal_3118, Inst_bSbox_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T26_U1 ( .a ({new_AGEMA_signal_2852, Inst_bSbox_T3}), .b ({new_AGEMA_signal_3004, Inst_bSbox_T16}), .c ({new_AGEMA_signal_3038, Inst_bSbox_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_T27_U1 ( .a ({new_AGEMA_signal_2850, Inst_bSbox_T1}), .b ({new_AGEMA_signal_2857, Inst_bSbox_T12}), .c ({new_AGEMA_signal_3007, Inst_bSbox_T27}) ) ;
    INV_X1 nReset_reg_U1 ( .A (nReset), .ZN (n10) ) ;
    ClockGatingController #(5) ClockGatingInst ( .clk (clk), .rst (start), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M1_U1 ( .a ({new_AGEMA_signal_3002, Inst_bSbox_T13}), .b ({new_AGEMA_signal_3000, Inst_bSbox_T6}), .clk (clk), .r ({Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_3039, Inst_bSbox_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M2_U1 ( .a ({new_AGEMA_signal_3037, Inst_bSbox_T23}), .b ({new_AGEMA_signal_3032, Inst_bSbox_T8}), .clk (clk), .r ({Fresh[3], Fresh[2]}), .c ({new_AGEMA_signal_3119, Inst_bSbox_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M3_U1 ( .a ({new_AGEMA_signal_3034, Inst_bSbox_T14}), .b ({new_AGEMA_signal_3039, Inst_bSbox_M1}), .c ({new_AGEMA_signal_3120, Inst_bSbox_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M4_U1 ( .a ({new_AGEMA_signal_3005, Inst_bSbox_T19}), .b ({new_AGEMA_signal_2826, SboxIn[0]}), .clk (clk), .r ({Fresh[5], Fresh[4]}), .c ({new_AGEMA_signal_3040, Inst_bSbox_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M5_U1 ( .a ({new_AGEMA_signal_3040, Inst_bSbox_M4}), .b ({new_AGEMA_signal_3039, Inst_bSbox_M1}), .c ({new_AGEMA_signal_3121, Inst_bSbox_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M6_U1 ( .a ({new_AGEMA_signal_2852, Inst_bSbox_T3}), .b ({new_AGEMA_signal_3004, Inst_bSbox_T16}), .clk (clk), .r ({Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_3041, Inst_bSbox_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M7_U1 ( .a ({new_AGEMA_signal_3006, Inst_bSbox_T22}), .b ({new_AGEMA_signal_3001, Inst_bSbox_T9}), .clk (clk), .r ({Fresh[9], Fresh[8]}), .c ({new_AGEMA_signal_3042, Inst_bSbox_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M8_U1 ( .a ({new_AGEMA_signal_3038, Inst_bSbox_T26}), .b ({new_AGEMA_signal_3041, Inst_bSbox_M6}), .c ({new_AGEMA_signal_3122, Inst_bSbox_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M9_U1 ( .a ({new_AGEMA_signal_3036, Inst_bSbox_T20}), .b ({new_AGEMA_signal_3035, Inst_bSbox_T17}), .clk (clk), .r ({Fresh[11], Fresh[10]}), .c ({new_AGEMA_signal_3123, Inst_bSbox_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M10_U1 ( .a ({new_AGEMA_signal_3123, Inst_bSbox_M9}), .b ({new_AGEMA_signal_3041, Inst_bSbox_M6}), .c ({new_AGEMA_signal_3262, Inst_bSbox_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M11_U1 ( .a ({new_AGEMA_signal_2850, Inst_bSbox_T1}), .b ({new_AGEMA_signal_3003, Inst_bSbox_T15}), .clk (clk), .r ({Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_3043, Inst_bSbox_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M12_U1 ( .a ({new_AGEMA_signal_2853, Inst_bSbox_T4}), .b ({new_AGEMA_signal_3007, Inst_bSbox_T27}), .clk (clk), .r ({Fresh[15], Fresh[14]}), .c ({new_AGEMA_signal_3044, Inst_bSbox_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M13_U1 ( .a ({new_AGEMA_signal_3044, Inst_bSbox_M12}), .b ({new_AGEMA_signal_3043, Inst_bSbox_M11}), .c ({new_AGEMA_signal_3124, Inst_bSbox_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M14_U1 ( .a ({new_AGEMA_signal_2851, Inst_bSbox_T2}), .b ({new_AGEMA_signal_3033, Inst_bSbox_T10}), .clk (clk), .r ({Fresh[17], Fresh[16]}), .c ({new_AGEMA_signal_3125, Inst_bSbox_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M15_U1 ( .a ({new_AGEMA_signal_3125, Inst_bSbox_M14}), .b ({new_AGEMA_signal_3043, Inst_bSbox_M11}), .c ({new_AGEMA_signal_3263, Inst_bSbox_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M16_U1 ( .a ({new_AGEMA_signal_3120, Inst_bSbox_M3}), .b ({new_AGEMA_signal_3119, Inst_bSbox_M2}), .c ({new_AGEMA_signal_3264, Inst_bSbox_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M17_U1 ( .a ({new_AGEMA_signal_3121, Inst_bSbox_M5}), .b ({new_AGEMA_signal_3117, Inst_bSbox_T24}), .c ({new_AGEMA_signal_3265, Inst_bSbox_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M18_U1 ( .a ({new_AGEMA_signal_3122, Inst_bSbox_M8}), .b ({new_AGEMA_signal_3042, Inst_bSbox_M7}), .c ({new_AGEMA_signal_3266, Inst_bSbox_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M19_U1 ( .a ({new_AGEMA_signal_3262, Inst_bSbox_M10}), .b ({new_AGEMA_signal_3263, Inst_bSbox_M15}), .c ({new_AGEMA_signal_3371, Inst_bSbox_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M20_U1 ( .a ({new_AGEMA_signal_3264, Inst_bSbox_M16}), .b ({new_AGEMA_signal_3124, Inst_bSbox_M13}), .c ({new_AGEMA_signal_3372, Inst_bSbox_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M21_U1 ( .a ({new_AGEMA_signal_3265, Inst_bSbox_M17}), .b ({new_AGEMA_signal_3263, Inst_bSbox_M15}), .c ({new_AGEMA_signal_3373, Inst_bSbox_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M22_U1 ( .a ({new_AGEMA_signal_3266, Inst_bSbox_M18}), .b ({new_AGEMA_signal_3124, Inst_bSbox_M13}), .c ({new_AGEMA_signal_3374, Inst_bSbox_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M23_U1 ( .a ({new_AGEMA_signal_3371, Inst_bSbox_M19}), .b ({new_AGEMA_signal_3118, Inst_bSbox_T25}), .c ({new_AGEMA_signal_3383, Inst_bSbox_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M24_U1 ( .a ({new_AGEMA_signal_3374, Inst_bSbox_M22}), .b ({new_AGEMA_signal_3383, Inst_bSbox_M23}), .c ({new_AGEMA_signal_3387, Inst_bSbox_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M27_U1 ( .a ({new_AGEMA_signal_3372, Inst_bSbox_M20}), .b ({new_AGEMA_signal_3373, Inst_bSbox_M21}), .c ({new_AGEMA_signal_3385, Inst_bSbox_M27}) ) ;

    /* cells in depth 2 */
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M25_U1 ( .a ({new_AGEMA_signal_3374, Inst_bSbox_M22}), .b ({new_AGEMA_signal_3372, Inst_bSbox_M20}), .clk (clk), .r ({Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_3384, Inst_bSbox_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M26_U1 ( .a ({new_AGEMA_signal_3373, Inst_bSbox_M21}), .b ({new_AGEMA_signal_3384, Inst_bSbox_M25}), .c ({new_AGEMA_signal_3388, Inst_bSbox_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M28_U1 ( .a ({new_AGEMA_signal_3383, Inst_bSbox_M23}), .b ({new_AGEMA_signal_3384, Inst_bSbox_M25}), .c ({new_AGEMA_signal_3389, Inst_bSbox_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M31_U1 ( .a ({new_AGEMA_signal_3372, Inst_bSbox_M20}), .b ({new_AGEMA_signal_3383, Inst_bSbox_M23}), .clk (clk), .r ({Fresh[21], Fresh[20]}), .c ({new_AGEMA_signal_3390, Inst_bSbox_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M33_U1 ( .a ({new_AGEMA_signal_3385, Inst_bSbox_M27}), .b ({new_AGEMA_signal_3384, Inst_bSbox_M25}), .c ({new_AGEMA_signal_3391, Inst_bSbox_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M34_U1 ( .a ({new_AGEMA_signal_3373, Inst_bSbox_M21}), .b ({new_AGEMA_signal_3374, Inst_bSbox_M22}), .clk (clk), .r ({Fresh[23], Fresh[22]}), .c ({new_AGEMA_signal_3386, Inst_bSbox_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M36_U1 ( .a ({new_AGEMA_signal_3387, Inst_bSbox_M24}), .b ({new_AGEMA_signal_3384, Inst_bSbox_M25}), .c ({new_AGEMA_signal_3396, Inst_bSbox_M36}) ) ;

    /* cells in depth 3 */
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M29_U1 ( .a ({new_AGEMA_signal_3389, Inst_bSbox_M28}), .b ({new_AGEMA_signal_3385, Inst_bSbox_M27}), .clk (clk), .r ({Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_3392, Inst_bSbox_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M30_U1 ( .a ({new_AGEMA_signal_3388, Inst_bSbox_M26}), .b ({new_AGEMA_signal_3387, Inst_bSbox_M24}), .clk (clk), .r ({Fresh[27], Fresh[26]}), .c ({new_AGEMA_signal_3393, Inst_bSbox_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M32_U1 ( .a ({new_AGEMA_signal_3385, Inst_bSbox_M27}), .b ({new_AGEMA_signal_3390, Inst_bSbox_M31}), .clk (clk), .r ({Fresh[29], Fresh[28]}), .c ({new_AGEMA_signal_3394, Inst_bSbox_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M35_U1 ( .a ({new_AGEMA_signal_3387, Inst_bSbox_M24}), .b ({new_AGEMA_signal_3386, Inst_bSbox_M34}), .clk (clk), .r ({Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_3395, Inst_bSbox_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M37_U1 ( .a ({new_AGEMA_signal_3373, Inst_bSbox_M21}), .b ({new_AGEMA_signal_3392, Inst_bSbox_M29}), .c ({new_AGEMA_signal_3397, Inst_bSbox_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M38_U1 ( .a ({new_AGEMA_signal_3394, Inst_bSbox_M32}), .b ({new_AGEMA_signal_3391, Inst_bSbox_M33}), .c ({new_AGEMA_signal_3398, Inst_bSbox_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M39_U1 ( .a ({new_AGEMA_signal_3383, Inst_bSbox_M23}), .b ({new_AGEMA_signal_3393, Inst_bSbox_M30}), .c ({new_AGEMA_signal_3399, Inst_bSbox_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M40_U1 ( .a ({new_AGEMA_signal_3395, Inst_bSbox_M35}), .b ({new_AGEMA_signal_3396, Inst_bSbox_M36}), .c ({new_AGEMA_signal_3400, Inst_bSbox_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M41_U1 ( .a ({new_AGEMA_signal_3398, Inst_bSbox_M38}), .b ({new_AGEMA_signal_3400, Inst_bSbox_M40}), .c ({new_AGEMA_signal_3401, Inst_bSbox_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M42_U1 ( .a ({new_AGEMA_signal_3397, Inst_bSbox_M37}), .b ({new_AGEMA_signal_3399, Inst_bSbox_M39}), .c ({new_AGEMA_signal_3402, Inst_bSbox_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M43_U1 ( .a ({new_AGEMA_signal_3397, Inst_bSbox_M37}), .b ({new_AGEMA_signal_3398, Inst_bSbox_M38}), .c ({new_AGEMA_signal_3403, Inst_bSbox_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M44_U1 ( .a ({new_AGEMA_signal_3399, Inst_bSbox_M39}), .b ({new_AGEMA_signal_3400, Inst_bSbox_M40}), .c ({new_AGEMA_signal_3404, Inst_bSbox_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_M45_U1 ( .a ({new_AGEMA_signal_3402, Inst_bSbox_M42}), .b ({new_AGEMA_signal_3401, Inst_bSbox_M41}), .c ({new_AGEMA_signal_3413, Inst_bSbox_M45}) ) ;

    /* cells in depth 4 */
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateIn_mux_inst_0_U1 ( .s (intFinal), .b ({new_AGEMA_signal_3454, SboxOut[0]}), .a ({new_AGEMA_signal_1984, StateOutXORroundKey[0]}), .c ({new_AGEMA_signal_3455, StateIn[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateIn_mux_inst_1_U1 ( .s (intFinal), .b ({new_AGEMA_signal_3463, SboxOut[1]}), .a ({new_AGEMA_signal_1987, StateOutXORroundKey[1]}), .c ({new_AGEMA_signal_3464, StateIn[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateIn_mux_inst_2_U1 ( .s (intFinal), .b ({new_AGEMA_signal_3462, SboxOut[2]}), .a ({new_AGEMA_signal_1990, StateOutXORroundKey[2]}), .c ({new_AGEMA_signal_3465, StateIn[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateIn_mux_inst_3_U1 ( .s (intFinal), .b ({new_AGEMA_signal_3461, SboxOut[3]}), .a ({new_AGEMA_signal_1993, StateOutXORroundKey[3]}), .c ({new_AGEMA_signal_3466, StateIn[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateIn_mux_inst_4_U1 ( .s (intFinal), .b ({new_AGEMA_signal_3460, SboxOut[4]}), .a ({new_AGEMA_signal_1996, StateOutXORroundKey[4]}), .c ({new_AGEMA_signal_3467, StateIn[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateIn_mux_inst_5_U1 ( .s (intFinal), .b ({new_AGEMA_signal_3459, SboxOut[5]}), .a ({new_AGEMA_signal_1999, StateOutXORroundKey[5]}), .c ({new_AGEMA_signal_3468, StateIn[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateIn_mux_inst_6_U1 ( .s (intFinal), .b ({new_AGEMA_signal_3458, SboxOut[6]}), .a ({new_AGEMA_signal_2002, StateOutXORroundKey[6]}), .c ({new_AGEMA_signal_3469, StateIn[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) MUX_StateIn_mux_inst_7_U1 ( .s (intFinal), .b ({new_AGEMA_signal_3457, SboxOut[7]}), .a ({new_AGEMA_signal_2005, StateOutXORroundKey[7]}), .c ({new_AGEMA_signal_3470, StateIn[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S33reg_gff_1_SFF_0_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_3488, stateArray_inS33ser[0]}), .a ({ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_3497, stateArray_S33reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S33reg_gff_1_SFF_1_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_3499, stateArray_inS33ser[1]}), .a ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_3520, stateArray_S33reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S33reg_gff_1_SFF_2_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_3501, stateArray_inS33ser[2]}), .a ({ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_3521, stateArray_S33reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S33reg_gff_1_SFF_3_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_3503, stateArray_inS33ser[3]}), .a ({ciphertext_s1[11], ciphertext_s0[11]}), .c ({new_AGEMA_signal_3522, stateArray_S33reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S33reg_gff_1_SFF_4_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_3505, stateArray_inS33ser[4]}), .a ({ciphertext_s1[12], ciphertext_s0[12]}), .c ({new_AGEMA_signal_3523, stateArray_S33reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S33reg_gff_1_SFF_5_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_3507, stateArray_inS33ser[5]}), .a ({ciphertext_s1[13], ciphertext_s0[13]}), .c ({new_AGEMA_signal_3524, stateArray_S33reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S33reg_gff_1_SFF_6_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_3509, stateArray_inS33ser[6]}), .a ({ciphertext_s1[14], ciphertext_s0[14]}), .c ({new_AGEMA_signal_3525, stateArray_S33reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_S33reg_gff_1_SFF_7_MUXInst_U1 ( .s (stateArray_n13), .b ({new_AGEMA_signal_3511, stateArray_inS33ser[7]}), .a ({ciphertext_s1[15], ciphertext_s0[15]}), .c ({new_AGEMA_signal_3526, stateArray_S33reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_input_MC_mux_inst_0_U1 ( .s (stateArray_n22), .b ({new_AGEMA_signal_3455, StateIn[0]}), .a ({new_AGEMA_signal_2860, StateInMC[0]}), .c ({new_AGEMA_signal_3471, stateArray_input_MC[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_input_MC_mux_inst_1_U1 ( .s (stateArray_n22), .b ({new_AGEMA_signal_3464, StateIn[1]}), .a ({new_AGEMA_signal_2861, StateInMC[1]}), .c ({new_AGEMA_signal_3480, stateArray_input_MC[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_input_MC_mux_inst_2_U1 ( .s (stateArray_n22), .b ({new_AGEMA_signal_3465, StateIn[2]}), .a ({new_AGEMA_signal_2834, StateInMC[2]}), .c ({new_AGEMA_signal_3481, stateArray_input_MC[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_input_MC_mux_inst_3_U1 ( .s (stateArray_n22), .b ({new_AGEMA_signal_3466, StateIn[3]}), .a ({new_AGEMA_signal_2862, StateInMC[3]}), .c ({new_AGEMA_signal_3482, stateArray_input_MC[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_input_MC_mux_inst_4_U1 ( .s (stateArray_n22), .b ({new_AGEMA_signal_3467, StateIn[4]}), .a ({new_AGEMA_signal_2863, StateInMC[4]}), .c ({new_AGEMA_signal_3483, stateArray_input_MC[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_input_MC_mux_inst_5_U1 ( .s (stateArray_n22), .b ({new_AGEMA_signal_3468, StateIn[5]}), .a ({new_AGEMA_signal_2835, StateInMC[5]}), .c ({new_AGEMA_signal_3484, stateArray_input_MC[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_input_MC_mux_inst_6_U1 ( .s (stateArray_n22), .b ({new_AGEMA_signal_3469, StateIn[6]}), .a ({new_AGEMA_signal_2836, StateInMC[6]}), .c ({new_AGEMA_signal_3485, stateArray_input_MC[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_input_MC_mux_inst_7_U1 ( .s (stateArray_n22), .b ({new_AGEMA_signal_3470, StateIn[7]}), .a ({new_AGEMA_signal_2837, StateInMC[7]}), .c ({new_AGEMA_signal_3486, stateArray_input_MC[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS33ser_mux_inst_0_U1 ( .s (stateArray_n25), .b ({plaintext_s1[0], plaintext_s0[0]}), .a ({new_AGEMA_signal_3471, stateArray_input_MC[0]}), .c ({new_AGEMA_signal_3488, stateArray_inS33ser[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS33ser_mux_inst_1_U1 ( .s (stateArray_n25), .b ({plaintext_s1[1], plaintext_s0[1]}), .a ({new_AGEMA_signal_3480, stateArray_input_MC[1]}), .c ({new_AGEMA_signal_3499, stateArray_inS33ser[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS33ser_mux_inst_2_U1 ( .s (stateArray_n25), .b ({plaintext_s1[2], plaintext_s0[2]}), .a ({new_AGEMA_signal_3481, stateArray_input_MC[2]}), .c ({new_AGEMA_signal_3501, stateArray_inS33ser[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS33ser_mux_inst_3_U1 ( .s (stateArray_n25), .b ({plaintext_s1[3], plaintext_s0[3]}), .a ({new_AGEMA_signal_3482, stateArray_input_MC[3]}), .c ({new_AGEMA_signal_3503, stateArray_inS33ser[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS33ser_mux_inst_4_U1 ( .s (stateArray_n25), .b ({plaintext_s1[4], plaintext_s0[4]}), .a ({new_AGEMA_signal_3483, stateArray_input_MC[4]}), .c ({new_AGEMA_signal_3505, stateArray_inS33ser[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS33ser_mux_inst_5_U1 ( .s (stateArray_n25), .b ({plaintext_s1[5], plaintext_s0[5]}), .a ({new_AGEMA_signal_3484, stateArray_input_MC[5]}), .c ({new_AGEMA_signal_3507, stateArray_inS33ser[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS33ser_mux_inst_6_U1 ( .s (stateArray_n25), .b ({plaintext_s1[6], plaintext_s0[6]}), .a ({new_AGEMA_signal_3485, stateArray_input_MC[6]}), .c ({new_AGEMA_signal_3509, stateArray_inS33ser[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) stateArray_MUX_inS33ser_mux_inst_7_U1 ( .s (stateArray_n25), .b ({plaintext_s1[7], plaintext_s0[7]}), .a ({new_AGEMA_signal_3486, stateArray_input_MC[7]}), .c ({new_AGEMA_signal_3511, stateArray_inS33ser[7]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U42 ( .a ({new_AGEMA_signal_3472, KeyArray_n55}), .b ({new_AGEMA_signal_2004, keyStateIn[7]}), .c ({new_AGEMA_signal_3489, KeyArray_inS30par[7]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U41 ( .a ({1'b0, roundConstant[7]}), .b ({new_AGEMA_signal_3457, SboxOut[7]}), .c ({new_AGEMA_signal_3472, KeyArray_n55}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U40 ( .a ({new_AGEMA_signal_3473, KeyArray_n54}), .b ({new_AGEMA_signal_2001, keyStateIn[6]}), .c ({new_AGEMA_signal_3490, KeyArray_inS30par[6]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U39 ( .a ({1'b0, roundConstant[6]}), .b ({new_AGEMA_signal_3458, SboxOut[6]}), .c ({new_AGEMA_signal_3473, KeyArray_n54}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U38 ( .a ({new_AGEMA_signal_3474, KeyArray_n53}), .b ({new_AGEMA_signal_1998, keyStateIn[5]}), .c ({new_AGEMA_signal_3491, KeyArray_inS30par[5]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U37 ( .a ({1'b0, roundConstant[5]}), .b ({new_AGEMA_signal_3459, SboxOut[5]}), .c ({new_AGEMA_signal_3474, KeyArray_n53}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U36 ( .a ({new_AGEMA_signal_3475, KeyArray_n52}), .b ({new_AGEMA_signal_1995, keyStateIn[4]}), .c ({new_AGEMA_signal_3492, KeyArray_inS30par[4]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U35 ( .a ({1'b0, roundConstant[4]}), .b ({new_AGEMA_signal_3460, SboxOut[4]}), .c ({new_AGEMA_signal_3475, KeyArray_n52}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U34 ( .a ({new_AGEMA_signal_3476, KeyArray_n51}), .b ({new_AGEMA_signal_1992, keyStateIn[3]}), .c ({new_AGEMA_signal_3493, KeyArray_inS30par[3]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U33 ( .a ({1'b0, roundConstant[3]}), .b ({new_AGEMA_signal_3461, SboxOut[3]}), .c ({new_AGEMA_signal_3476, KeyArray_n51}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U32 ( .a ({new_AGEMA_signal_3477, KeyArray_n50}), .b ({new_AGEMA_signal_1989, keyStateIn[2]}), .c ({new_AGEMA_signal_3494, KeyArray_inS30par[2]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U31 ( .a ({1'b0, roundConstant[2]}), .b ({new_AGEMA_signal_3462, SboxOut[2]}), .c ({new_AGEMA_signal_3477, KeyArray_n50}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U30 ( .a ({new_AGEMA_signal_3478, KeyArray_n49}), .b ({new_AGEMA_signal_1986, keyStateIn[1]}), .c ({new_AGEMA_signal_3495, KeyArray_inS30par[1]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U29 ( .a ({1'b0, roundConstant[1]}), .b ({new_AGEMA_signal_3463, SboxOut[1]}), .c ({new_AGEMA_signal_3478, KeyArray_n49}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U28 ( .a ({new_AGEMA_signal_3456, KeyArray_n48}), .b ({new_AGEMA_signal_1983, keyStateIn[0]}), .c ({new_AGEMA_signal_3479, KeyArray_inS30par[0]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) KeyArray_U27 ( .a ({1'b0, roundConstant[0]}), .b ({new_AGEMA_signal_3454, SboxOut[0]}), .c ({new_AGEMA_signal_3456, KeyArray_n48}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_0_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2683, KeyArray_outS30ser[0]}), .a ({new_AGEMA_signal_3496, KeyArray_S30reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_3512, KeyArray_S30reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2708, KeyArray_inS30ser[0]}), .a ({new_AGEMA_signal_3479, KeyArray_inS30par[0]}), .c ({new_AGEMA_signal_3496, KeyArray_S30reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_1_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2686, KeyArray_outS30ser[1]}), .a ({new_AGEMA_signal_3513, KeyArray_S30reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_3527, KeyArray_S30reg_gff_1_SFF_1_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2711, KeyArray_inS30ser[1]}), .a ({new_AGEMA_signal_3495, KeyArray_inS30par[1]}), .c ({new_AGEMA_signal_3513, KeyArray_S30reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_2_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2689, KeyArray_outS30ser[2]}), .a ({new_AGEMA_signal_3514, KeyArray_S30reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_3528, KeyArray_S30reg_gff_1_SFF_2_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2714, KeyArray_inS30ser[2]}), .a ({new_AGEMA_signal_3494, KeyArray_inS30par[2]}), .c ({new_AGEMA_signal_3514, KeyArray_S30reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_3_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2692, KeyArray_outS30ser[3]}), .a ({new_AGEMA_signal_3515, KeyArray_S30reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_3529, KeyArray_S30reg_gff_1_SFF_3_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2717, KeyArray_inS30ser[3]}), .a ({new_AGEMA_signal_3493, KeyArray_inS30par[3]}), .c ({new_AGEMA_signal_3515, KeyArray_S30reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_4_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2695, KeyArray_outS30ser[4]}), .a ({new_AGEMA_signal_3516, KeyArray_S30reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_3530, KeyArray_S30reg_gff_1_SFF_4_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2720, KeyArray_inS30ser[4]}), .a ({new_AGEMA_signal_3492, KeyArray_inS30par[4]}), .c ({new_AGEMA_signal_3516, KeyArray_S30reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_5_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2698, KeyArray_outS30ser[5]}), .a ({new_AGEMA_signal_3517, KeyArray_S30reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_3531, KeyArray_S30reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2723, KeyArray_inS30ser[5]}), .a ({new_AGEMA_signal_3491, KeyArray_inS30par[5]}), .c ({new_AGEMA_signal_3517, KeyArray_S30reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_6_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2701, KeyArray_outS30ser[6]}), .a ({new_AGEMA_signal_3518, KeyArray_S30reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_3532, KeyArray_S30reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2726, KeyArray_inS30ser[6]}), .a ({new_AGEMA_signal_3490, KeyArray_inS30par[6]}), .c ({new_AGEMA_signal_3518, KeyArray_S30reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_7_U1 ( .s (KeyArray_n23), .b ({new_AGEMA_signal_2704, KeyArray_outS30ser[7]}), .a ({new_AGEMA_signal_3519, KeyArray_S30reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_3533, KeyArray_S30reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1 ( .s (KeyArray_n31), .b ({new_AGEMA_signal_2729, KeyArray_inS30ser[7]}), .a ({new_AGEMA_signal_3489, KeyArray_inS30par[7]}), .c ({new_AGEMA_signal_3519, KeyArray_S30reg_gff_1_SFF_7_QD}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M46_U1 ( .a ({new_AGEMA_signal_3404, Inst_bSbox_M44}), .b ({new_AGEMA_signal_3000, Inst_bSbox_T6}), .clk (clk), .r ({Fresh[33], Fresh[32]}), .c ({new_AGEMA_signal_3414, Inst_bSbox_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M47_U1 ( .a ({new_AGEMA_signal_3400, Inst_bSbox_M40}), .b ({new_AGEMA_signal_3032, Inst_bSbox_T8}), .clk (clk), .r ({Fresh[35], Fresh[34]}), .c ({new_AGEMA_signal_3405, Inst_bSbox_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M48_U1 ( .a ({new_AGEMA_signal_3399, Inst_bSbox_M39}), .b ({new_AGEMA_signal_2826, SboxIn[0]}), .clk (clk), .r ({Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_3406, Inst_bSbox_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M49_U1 ( .a ({new_AGEMA_signal_3403, Inst_bSbox_M43}), .b ({new_AGEMA_signal_3004, Inst_bSbox_T16}), .clk (clk), .r ({Fresh[39], Fresh[38]}), .c ({new_AGEMA_signal_3415, Inst_bSbox_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M50_U1 ( .a ({new_AGEMA_signal_3398, Inst_bSbox_M38}), .b ({new_AGEMA_signal_3001, Inst_bSbox_T9}), .clk (clk), .r ({Fresh[41], Fresh[40]}), .c ({new_AGEMA_signal_3407, Inst_bSbox_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M51_U1 ( .a ({new_AGEMA_signal_3397, Inst_bSbox_M37}), .b ({new_AGEMA_signal_3035, Inst_bSbox_T17}), .clk (clk), .r ({Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_3408, Inst_bSbox_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M52_U1 ( .a ({new_AGEMA_signal_3402, Inst_bSbox_M42}), .b ({new_AGEMA_signal_3003, Inst_bSbox_T15}), .clk (clk), .r ({Fresh[45], Fresh[44]}), .c ({new_AGEMA_signal_3416, Inst_bSbox_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M53_U1 ( .a ({new_AGEMA_signal_3413, Inst_bSbox_M45}), .b ({new_AGEMA_signal_3007, Inst_bSbox_T27}), .clk (clk), .r ({Fresh[47], Fresh[46]}), .c ({new_AGEMA_signal_3425, Inst_bSbox_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M54_U1 ( .a ({new_AGEMA_signal_3401, Inst_bSbox_M41}), .b ({new_AGEMA_signal_3033, Inst_bSbox_T10}), .clk (clk), .r ({Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_3417, Inst_bSbox_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M55_U1 ( .a ({new_AGEMA_signal_3404, Inst_bSbox_M44}), .b ({new_AGEMA_signal_3002, Inst_bSbox_T13}), .clk (clk), .r ({Fresh[51], Fresh[50]}), .c ({new_AGEMA_signal_3418, Inst_bSbox_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M56_U1 ( .a ({new_AGEMA_signal_3400, Inst_bSbox_M40}), .b ({new_AGEMA_signal_3037, Inst_bSbox_T23}), .clk (clk), .r ({Fresh[53], Fresh[52]}), .c ({new_AGEMA_signal_3409, Inst_bSbox_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M57_U1 ( .a ({new_AGEMA_signal_3399, Inst_bSbox_M39}), .b ({new_AGEMA_signal_3005, Inst_bSbox_T19}), .clk (clk), .r ({Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_3410, Inst_bSbox_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M58_U1 ( .a ({new_AGEMA_signal_3403, Inst_bSbox_M43}), .b ({new_AGEMA_signal_2852, Inst_bSbox_T3}), .clk (clk), .r ({Fresh[57], Fresh[56]}), .c ({new_AGEMA_signal_3419, Inst_bSbox_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M59_U1 ( .a ({new_AGEMA_signal_3398, Inst_bSbox_M38}), .b ({new_AGEMA_signal_3006, Inst_bSbox_T22}), .clk (clk), .r ({Fresh[59], Fresh[58]}), .c ({new_AGEMA_signal_3411, Inst_bSbox_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M60_U1 ( .a ({new_AGEMA_signal_3397, Inst_bSbox_M37}), .b ({new_AGEMA_signal_3036, Inst_bSbox_T20}), .clk (clk), .r ({Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_3412, Inst_bSbox_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M61_U1 ( .a ({new_AGEMA_signal_3402, Inst_bSbox_M42}), .b ({new_AGEMA_signal_2850, Inst_bSbox_T1}), .clk (clk), .r ({Fresh[63], Fresh[62]}), .c ({new_AGEMA_signal_3420, Inst_bSbox_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M62_U1 ( .a ({new_AGEMA_signal_3413, Inst_bSbox_M45}), .b ({new_AGEMA_signal_2853, Inst_bSbox_T4}), .clk (clk), .r ({Fresh[65], Fresh[64]}), .c ({new_AGEMA_signal_3426, Inst_bSbox_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_AND_M63_U1 ( .a ({new_AGEMA_signal_3401, Inst_bSbox_M41}), .b ({new_AGEMA_signal_2851, Inst_bSbox_T2}), .clk (clk), .r ({Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_3421, Inst_bSbox_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L0_U1 ( .a ({new_AGEMA_signal_3420, Inst_bSbox_M61}), .b ({new_AGEMA_signal_3426, Inst_bSbox_M62}), .c ({new_AGEMA_signal_3435, Inst_bSbox_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L1_U1 ( .a ({new_AGEMA_signal_3407, Inst_bSbox_M50}), .b ({new_AGEMA_signal_3409, Inst_bSbox_M56}), .c ({new_AGEMA_signal_3422, Inst_bSbox_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L2_U1 ( .a ({new_AGEMA_signal_3414, Inst_bSbox_M46}), .b ({new_AGEMA_signal_3406, Inst_bSbox_M48}), .c ({new_AGEMA_signal_3427, Inst_bSbox_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L3_U1 ( .a ({new_AGEMA_signal_3405, Inst_bSbox_M47}), .b ({new_AGEMA_signal_3418, Inst_bSbox_M55}), .c ({new_AGEMA_signal_3428, Inst_bSbox_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L4_U1 ( .a ({new_AGEMA_signal_3417, Inst_bSbox_M54}), .b ({new_AGEMA_signal_3419, Inst_bSbox_M58}), .c ({new_AGEMA_signal_3429, Inst_bSbox_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L5_U1 ( .a ({new_AGEMA_signal_3415, Inst_bSbox_M49}), .b ({new_AGEMA_signal_3420, Inst_bSbox_M61}), .c ({new_AGEMA_signal_3430, Inst_bSbox_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L6_U1 ( .a ({new_AGEMA_signal_3426, Inst_bSbox_M62}), .b ({new_AGEMA_signal_3430, Inst_bSbox_L5}), .c ({new_AGEMA_signal_3436, Inst_bSbox_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L7_U1 ( .a ({new_AGEMA_signal_3414, Inst_bSbox_M46}), .b ({new_AGEMA_signal_3428, Inst_bSbox_L3}), .c ({new_AGEMA_signal_3437, Inst_bSbox_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L8_U1 ( .a ({new_AGEMA_signal_3408, Inst_bSbox_M51}), .b ({new_AGEMA_signal_3411, Inst_bSbox_M59}), .c ({new_AGEMA_signal_3423, Inst_bSbox_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L9_U1 ( .a ({new_AGEMA_signal_3416, Inst_bSbox_M52}), .b ({new_AGEMA_signal_3425, Inst_bSbox_M53}), .c ({new_AGEMA_signal_3438, Inst_bSbox_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L10_U1 ( .a ({new_AGEMA_signal_3425, Inst_bSbox_M53}), .b ({new_AGEMA_signal_3429, Inst_bSbox_L4}), .c ({new_AGEMA_signal_3439, Inst_bSbox_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L11_U1 ( .a ({new_AGEMA_signal_3412, Inst_bSbox_M60}), .b ({new_AGEMA_signal_3427, Inst_bSbox_L2}), .c ({new_AGEMA_signal_3440, Inst_bSbox_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L12_U1 ( .a ({new_AGEMA_signal_3406, Inst_bSbox_M48}), .b ({new_AGEMA_signal_3408, Inst_bSbox_M51}), .c ({new_AGEMA_signal_3424, Inst_bSbox_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L13_U1 ( .a ({new_AGEMA_signal_3407, Inst_bSbox_M50}), .b ({new_AGEMA_signal_3435, Inst_bSbox_L0}), .c ({new_AGEMA_signal_3444, Inst_bSbox_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L14_U1 ( .a ({new_AGEMA_signal_3416, Inst_bSbox_M52}), .b ({new_AGEMA_signal_3420, Inst_bSbox_M61}), .c ({new_AGEMA_signal_3431, Inst_bSbox_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L15_U1 ( .a ({new_AGEMA_signal_3418, Inst_bSbox_M55}), .b ({new_AGEMA_signal_3422, Inst_bSbox_L1}), .c ({new_AGEMA_signal_3432, Inst_bSbox_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L16_U1 ( .a ({new_AGEMA_signal_3409, Inst_bSbox_M56}), .b ({new_AGEMA_signal_3435, Inst_bSbox_L0}), .c ({new_AGEMA_signal_3445, Inst_bSbox_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L17_U1 ( .a ({new_AGEMA_signal_3410, Inst_bSbox_M57}), .b ({new_AGEMA_signal_3422, Inst_bSbox_L1}), .c ({new_AGEMA_signal_3433, Inst_bSbox_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L18_U1 ( .a ({new_AGEMA_signal_3419, Inst_bSbox_M58}), .b ({new_AGEMA_signal_3423, Inst_bSbox_L8}), .c ({new_AGEMA_signal_3434, Inst_bSbox_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L19_U1 ( .a ({new_AGEMA_signal_3421, Inst_bSbox_M63}), .b ({new_AGEMA_signal_3429, Inst_bSbox_L4}), .c ({new_AGEMA_signal_3441, Inst_bSbox_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L20_U1 ( .a ({new_AGEMA_signal_3435, Inst_bSbox_L0}), .b ({new_AGEMA_signal_3422, Inst_bSbox_L1}), .c ({new_AGEMA_signal_3446, Inst_bSbox_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L21_U1 ( .a ({new_AGEMA_signal_3422, Inst_bSbox_L1}), .b ({new_AGEMA_signal_3437, Inst_bSbox_L7}), .c ({new_AGEMA_signal_3447, Inst_bSbox_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L22_U1 ( .a ({new_AGEMA_signal_3428, Inst_bSbox_L3}), .b ({new_AGEMA_signal_3424, Inst_bSbox_L12}), .c ({new_AGEMA_signal_3442, Inst_bSbox_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L23_U1 ( .a ({new_AGEMA_signal_3434, Inst_bSbox_L18}), .b ({new_AGEMA_signal_3427, Inst_bSbox_L2}), .c ({new_AGEMA_signal_3443, Inst_bSbox_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L24_U1 ( .a ({new_AGEMA_signal_3432, Inst_bSbox_L15}), .b ({new_AGEMA_signal_3438, Inst_bSbox_L9}), .c ({new_AGEMA_signal_3448, Inst_bSbox_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L25_U1 ( .a ({new_AGEMA_signal_3436, Inst_bSbox_L6}), .b ({new_AGEMA_signal_3439, Inst_bSbox_L10}), .c ({new_AGEMA_signal_3449, Inst_bSbox_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L26_U1 ( .a ({new_AGEMA_signal_3437, Inst_bSbox_L7}), .b ({new_AGEMA_signal_3438, Inst_bSbox_L9}), .c ({new_AGEMA_signal_3450, Inst_bSbox_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L27_U1 ( .a ({new_AGEMA_signal_3423, Inst_bSbox_L8}), .b ({new_AGEMA_signal_3439, Inst_bSbox_L10}), .c ({new_AGEMA_signal_3451, Inst_bSbox_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L28_U1 ( .a ({new_AGEMA_signal_3440, Inst_bSbox_L11}), .b ({new_AGEMA_signal_3431, Inst_bSbox_L14}), .c ({new_AGEMA_signal_3452, Inst_bSbox_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_L29_U1 ( .a ({new_AGEMA_signal_3440, Inst_bSbox_L11}), .b ({new_AGEMA_signal_3433, Inst_bSbox_L17}), .c ({new_AGEMA_signal_3453, Inst_bSbox_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_S0_U1 ( .a ({new_AGEMA_signal_3436, Inst_bSbox_L6}), .b ({new_AGEMA_signal_3448, Inst_bSbox_L24}), .c ({new_AGEMA_signal_3457, SboxOut[7]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_S1_U1 ( .a ({new_AGEMA_signal_3445, Inst_bSbox_L16}), .b ({new_AGEMA_signal_3450, Inst_bSbox_L26}), .c ({new_AGEMA_signal_3458, SboxOut[6]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_S2_U1 ( .a ({new_AGEMA_signal_3441, Inst_bSbox_L19}), .b ({new_AGEMA_signal_3452, Inst_bSbox_L28}), .c ({new_AGEMA_signal_3459, SboxOut[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_S3_U1 ( .a ({new_AGEMA_signal_3436, Inst_bSbox_L6}), .b ({new_AGEMA_signal_3447, Inst_bSbox_L21}), .c ({new_AGEMA_signal_3460, SboxOut[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_S4_U1 ( .a ({new_AGEMA_signal_3446, Inst_bSbox_L20}), .b ({new_AGEMA_signal_3442, Inst_bSbox_L22}), .c ({new_AGEMA_signal_3461, SboxOut[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_S5_U1 ( .a ({new_AGEMA_signal_3449, Inst_bSbox_L25}), .b ({new_AGEMA_signal_3453, Inst_bSbox_L29}), .c ({new_AGEMA_signal_3462, SboxOut[2]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_S6_U1 ( .a ({new_AGEMA_signal_3444, Inst_bSbox_L13}), .b ({new_AGEMA_signal_3451, Inst_bSbox_L27}), .c ({new_AGEMA_signal_3463, SboxOut[1]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(0)) Inst_bSbox_XOR_S7_U1 ( .a ({new_AGEMA_signal_3436, Inst_bSbox_L6}), .b ({new_AGEMA_signal_3443, Inst_bSbox_L23}), .c ({new_AGEMA_signal_3454, SboxOut[0]}) ) ;

    /* register cells */
    DFF_X1 ctrl_seq6_SFF_0_Q_reg_FF_FF ( .CK (clk_gated), .D (ctrl_seq6_SFF_0_QD), .Q (ctrl_seq6In_1_), .QN () ) ;
    DFF_X1 ctrl_seq6_SFF_1_Q_reg_FF_FF ( .CK (clk_gated), .D (ctrl_seq6_SFF_1_QD), .Q (ctrl_seq6In_2_), .QN () ) ;
    DFF_X1 ctrl_seq6_SFF_2_Q_reg_FF_FF ( .CK (clk_gated), .D (ctrl_seq6_SFF_2_QD), .Q (ctrl_seq6In_3_), .QN () ) ;
    DFF_X1 ctrl_seq6_SFF_3_Q_reg_FF_FF ( .CK (clk_gated), .D (ctrl_seq6_SFF_3_QD), .Q (ctrl_seq6In_4_), .QN () ) ;
    DFF_X1 ctrl_seq6_SFF_4_Q_reg_FF_FF ( .CK (clk_gated), .D (ctrl_seq6_SFF_4_QD), .Q (ctrl_seq6Out_4_), .QN () ) ;
    DFF_X1 ctrl_seq4_SFF_0_Q_reg_FF_FF ( .CK (clk_gated), .D (ctrl_seq4_SFF_0_QD), .Q (ctrl_seq4In_1_), .QN () ) ;
    DFF_X1 ctrl_seq4_SFF_1_Q_reg_FF_FF ( .CK (clk_gated), .D (ctrl_seq4_SFF_1_QD), .Q (ctrl_seq4Out_1_), .QN () ) ;
    DFF_X1 ctrl_CSselMC_reg_FF_FF ( .CK (clk_gated), .D (ctrl_N14), .Q (ctrl_n6), .QN () ) ;
    DFF_X1 ctrl_CSenRC_reg_FF_FF ( .CK (clk_gated), .D (selSR), .Q (enRCon), .QN () ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3126, stateArray_S00reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3127, stateArray_S00reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3128, stateArray_S00reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3129, stateArray_S00reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3130, stateArray_S00reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3131, stateArray_S00reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3132, stateArray_S00reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3133, stateArray_S00reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3134, stateArray_S01reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3135, stateArray_S01reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3136, stateArray_S01reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3137, stateArray_S01reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3138, stateArray_S01reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3139, stateArray_S01reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3140, stateArray_S01reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3141, stateArray_S01reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3142, stateArray_S02reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3143, stateArray_S02reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3144, stateArray_S02reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3145, stateArray_S02reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3146, stateArray_S02reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3147, stateArray_S02reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3148, stateArray_S02reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3149, stateArray_S02reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3150, stateArray_S03reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3151, stateArray_S03reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3152, stateArray_S03reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3153, stateArray_S03reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3154, stateArray_S03reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3155, stateArray_S03reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3156, stateArray_S03reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3157, stateArray_S03reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3158, stateArray_S10reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3159, stateArray_S10reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3160, stateArray_S10reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3161, stateArray_S10reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3162, stateArray_S10reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3163, stateArray_S10reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3164, stateArray_S10reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3165, stateArray_S10reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3166, stateArray_S11reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3167, stateArray_S11reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3168, stateArray_S11reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3169, stateArray_S11reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3170, stateArray_S11reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3171, stateArray_S11reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3172, stateArray_S11reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3173, stateArray_S11reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3174, stateArray_S12reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3175, stateArray_S12reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3176, stateArray_S12reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3177, stateArray_S12reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3178, stateArray_S12reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3179, stateArray_S12reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3180, stateArray_S12reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3181, stateArray_S12reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3182, stateArray_S13reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3183, stateArray_S13reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3184, stateArray_S13reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3185, stateArray_S13reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3186, stateArray_S13reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3187, stateArray_S13reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3188, stateArray_S13reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3189, stateArray_S13reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3190, stateArray_S20reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3191, stateArray_S20reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3192, stateArray_S20reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3193, stateArray_S20reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3194, stateArray_S20reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3195, stateArray_S20reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3196, stateArray_S20reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3197, stateArray_S20reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3198, stateArray_S21reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3199, stateArray_S21reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3200, stateArray_S21reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3201, stateArray_S21reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3202, stateArray_S21reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3203, stateArray_S21reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3204, stateArray_S21reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3205, stateArray_S21reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3206, stateArray_S22reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3207, stateArray_S22reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3208, stateArray_S22reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3209, stateArray_S22reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3210, stateArray_S22reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3211, stateArray_S22reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3212, stateArray_S22reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3213, stateArray_S22reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3214, stateArray_S23reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3215, stateArray_S23reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3216, stateArray_S23reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3217, stateArray_S23reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3218, stateArray_S23reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3219, stateArray_S23reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3220, stateArray_S23reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3221, stateArray_S23reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3222, stateArray_S30reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3223, stateArray_S30reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3224, stateArray_S30reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3225, stateArray_S30reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3226, stateArray_S30reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3227, stateArray_S30reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3228, stateArray_S30reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3229, stateArray_S30reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3230, stateArray_S31reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3231, stateArray_S31reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3232, stateArray_S31reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3233, stateArray_S31reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3234, stateArray_S31reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3235, stateArray_S31reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3236, stateArray_S31reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3237, stateArray_S31reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3238, stateArray_S32reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3239, stateArray_S32reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3240, stateArray_S32reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3241, stateArray_S32reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3242, stateArray_S32reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3243, stateArray_S32reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3244, stateArray_S32reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3245, stateArray_S32reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3497, stateArray_S33reg_gff_1_SFF_0_QD}), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3520, stateArray_S33reg_gff_1_SFF_1_QD}), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3521, stateArray_S33reg_gff_1_SFF_2_QD}), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3522, stateArray_S33reg_gff_1_SFF_3_QD}), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3523, stateArray_S33reg_gff_1_SFF_4_QD}), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3524, stateArray_S33reg_gff_1_SFF_5_QD}), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3525, stateArray_S33reg_gff_1_SFF_6_QD}), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) stateArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3526, stateArray_S33reg_gff_1_SFF_7_QD}), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3375, KeyArray_S00reg_gff_1_SFF_0_n5}), .Q ({new_AGEMA_signal_1983, keyStateIn[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3376, KeyArray_S00reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_1986, keyStateIn[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3377, KeyArray_S00reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_1989, keyStateIn[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3378, KeyArray_S00reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_1992, keyStateIn[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3379, KeyArray_S00reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_1995, keyStateIn[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3380, KeyArray_S00reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_1998, keyStateIn[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3381, KeyArray_S00reg_gff_1_SFF_6_n6}), .Q ({new_AGEMA_signal_2001, keyStateIn[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3382, KeyArray_S00reg_gff_1_SFF_7_n6}), .Q ({new_AGEMA_signal_2004, keyStateIn[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3275, KeyArray_S01reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_2020, KeyArray_outS01ser_0_}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3276, KeyArray_S01reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_2018, KeyArray_outS01ser_1_}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3277, KeyArray_S01reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_2016, KeyArray_outS01ser_2_}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3278, KeyArray_S01reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_2014, KeyArray_outS01ser_3_}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3279, KeyArray_S01reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_2012, KeyArray_outS01ser_4_}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3280, KeyArray_S01reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_2010, KeyArray_outS01ser_5_}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3281, KeyArray_S01reg_gff_1_SFF_6_n6}), .Q ({new_AGEMA_signal_2008, KeyArray_outS01ser_6_}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3282, KeyArray_S01reg_gff_1_SFF_7_n6}), .Q ({new_AGEMA_signal_2006, KeyArray_outS01ser_7_}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3283, KeyArray_S02reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_2443, KeyArray_outS02ser[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3284, KeyArray_S02reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_2446, KeyArray_outS02ser[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3285, KeyArray_S02reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_2449, KeyArray_outS02ser[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3286, KeyArray_S02reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_2452, KeyArray_outS02ser[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3287, KeyArray_S02reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_2455, KeyArray_outS02ser[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3288, KeyArray_S02reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_2458, KeyArray_outS02ser[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3289, KeyArray_S02reg_gff_1_SFF_6_n6}), .Q ({new_AGEMA_signal_2461, KeyArray_outS02ser[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3290, KeyArray_S02reg_gff_1_SFF_7_n6}), .Q ({new_AGEMA_signal_2464, KeyArray_outS02ser[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3291, KeyArray_S03reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_2467, KeyArray_outS03ser[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3292, KeyArray_S03reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_2470, KeyArray_outS03ser[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3293, KeyArray_S03reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_2473, KeyArray_outS03ser[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3294, KeyArray_S03reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_2476, KeyArray_outS03ser[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3295, KeyArray_S03reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_2479, KeyArray_outS03ser[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3296, KeyArray_S03reg_gff_1_SFF_5_n5}), .Q ({new_AGEMA_signal_2482, KeyArray_outS03ser[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3297, KeyArray_S03reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_2485, KeyArray_outS03ser[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3298, KeyArray_S03reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_2488, KeyArray_outS03ser[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3299, KeyArray_S10reg_gff_1_SFF_0_n5}), .Q ({new_AGEMA_signal_2491, KeyArray_outS10ser[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3300, KeyArray_S10reg_gff_1_SFF_1_n5}), .Q ({new_AGEMA_signal_2494, KeyArray_outS10ser[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3301, KeyArray_S10reg_gff_1_SFF_2_n5}), .Q ({new_AGEMA_signal_2497, KeyArray_outS10ser[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3302, KeyArray_S10reg_gff_1_SFF_3_n5}), .Q ({new_AGEMA_signal_2500, KeyArray_outS10ser[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3303, KeyArray_S10reg_gff_1_SFF_4_n5}), .Q ({new_AGEMA_signal_2503, KeyArray_outS10ser[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3304, KeyArray_S10reg_gff_1_SFF_5_n5}), .Q ({new_AGEMA_signal_2506, KeyArray_outS10ser[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3305, KeyArray_S10reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_2509, KeyArray_outS10ser[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3306, KeyArray_S10reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_2512, KeyArray_outS10ser[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3307, KeyArray_S11reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_2515, KeyArray_outS11ser[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3308, KeyArray_S11reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_2518, KeyArray_outS11ser[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3309, KeyArray_S11reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_2521, KeyArray_outS11ser[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3310, KeyArray_S11reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_2524, KeyArray_outS11ser[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3311, KeyArray_S11reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_2527, KeyArray_outS11ser[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3312, KeyArray_S11reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_2530, KeyArray_outS11ser[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3313, KeyArray_S11reg_gff_1_SFF_6_n6}), .Q ({new_AGEMA_signal_2533, KeyArray_outS11ser[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3314, KeyArray_S11reg_gff_1_SFF_7_n6}), .Q ({new_AGEMA_signal_2536, KeyArray_outS11ser[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3093, KeyArray_S12reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_2539, KeyArray_outS12ser[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3094, KeyArray_S12reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_2542, KeyArray_outS12ser[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3095, KeyArray_S12reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_2545, KeyArray_outS12ser[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3096, KeyArray_S12reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_2548, KeyArray_outS12ser[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3097, KeyArray_S12reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_2551, KeyArray_outS12ser[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3098, KeyArray_S12reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_2554, KeyArray_outS12ser[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3099, KeyArray_S12reg_gff_1_SFF_6_n6}), .Q ({new_AGEMA_signal_2557, KeyArray_outS12ser[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3100, KeyArray_S12reg_gff_1_SFF_7_n6}), .Q ({new_AGEMA_signal_2560, KeyArray_outS12ser[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3101, KeyArray_S13reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_2563, keySBIn[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3102, KeyArray_S13reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_2566, keySBIn[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3103, KeyArray_S13reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_2569, keySBIn[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3104, KeyArray_S13reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_2572, keySBIn[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3105, KeyArray_S13reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_2575, keySBIn[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3106, KeyArray_S13reg_gff_1_SFF_5_n5}), .Q ({new_AGEMA_signal_2578, keySBIn[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3107, KeyArray_S13reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_2581, keySBIn[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3108, KeyArray_S13reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_2584, keySBIn[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3315, KeyArray_S20reg_gff_1_SFF_0_n5}), .Q ({new_AGEMA_signal_2587, KeyArray_outS20ser[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3316, KeyArray_S20reg_gff_1_SFF_1_n5}), .Q ({new_AGEMA_signal_2590, KeyArray_outS20ser[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3317, KeyArray_S20reg_gff_1_SFF_2_n5}), .Q ({new_AGEMA_signal_2593, KeyArray_outS20ser[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3318, KeyArray_S20reg_gff_1_SFF_3_n5}), .Q ({new_AGEMA_signal_2596, KeyArray_outS20ser[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3319, KeyArray_S20reg_gff_1_SFF_4_n5}), .Q ({new_AGEMA_signal_2599, KeyArray_outS20ser[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3320, KeyArray_S20reg_gff_1_SFF_5_n5}), .Q ({new_AGEMA_signal_2602, KeyArray_outS20ser[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3321, KeyArray_S20reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_2605, KeyArray_outS20ser[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3322, KeyArray_S20reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_2608, KeyArray_outS20ser[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3323, KeyArray_S21reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_2611, KeyArray_outS21ser[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3324, KeyArray_S21reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_2614, KeyArray_outS21ser[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3325, KeyArray_S21reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_2617, KeyArray_outS21ser[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3326, KeyArray_S21reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_2620, KeyArray_outS21ser[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3327, KeyArray_S21reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_2623, KeyArray_outS21ser[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3328, KeyArray_S21reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_2626, KeyArray_outS21ser[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3329, KeyArray_S21reg_gff_1_SFF_6_n6}), .Q ({new_AGEMA_signal_2629, KeyArray_outS21ser[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3330, KeyArray_S21reg_gff_1_SFF_7_n6}), .Q ({new_AGEMA_signal_2632, KeyArray_outS21ser[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3331, KeyArray_S22reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_2635, KeyArray_outS22ser[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3332, KeyArray_S22reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_2638, KeyArray_outS22ser[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3333, KeyArray_S22reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_2641, KeyArray_outS22ser[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3334, KeyArray_S22reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_2644, KeyArray_outS22ser[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3335, KeyArray_S22reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_2647, KeyArray_outS22ser[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3336, KeyArray_S22reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_2650, KeyArray_outS22ser[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3337, KeyArray_S22reg_gff_1_SFF_6_n6}), .Q ({new_AGEMA_signal_2653, KeyArray_outS22ser[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3338, KeyArray_S22reg_gff_1_SFF_7_n6}), .Q ({new_AGEMA_signal_2656, KeyArray_outS22ser[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3339, KeyArray_S23reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_2659, KeyArray_outS23ser[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3340, KeyArray_S23reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_2662, KeyArray_outS23ser[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3341, KeyArray_S23reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_2665, KeyArray_outS23ser[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3342, KeyArray_S23reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_2668, KeyArray_outS23ser[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3343, KeyArray_S23reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_2671, KeyArray_outS23ser[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3344, KeyArray_S23reg_gff_1_SFF_5_n5}), .Q ({new_AGEMA_signal_2674, KeyArray_outS23ser[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3345, KeyArray_S23reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_2677, KeyArray_outS23ser[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3346, KeyArray_S23reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_2680, KeyArray_outS23ser[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3512, KeyArray_S30reg_gff_1_SFF_0_n5}), .Q ({new_AGEMA_signal_2683, KeyArray_outS30ser[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3527, KeyArray_S30reg_gff_1_SFF_1_n5}), .Q ({new_AGEMA_signal_2686, KeyArray_outS30ser[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3528, KeyArray_S30reg_gff_1_SFF_2_n5}), .Q ({new_AGEMA_signal_2689, KeyArray_outS30ser[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3529, KeyArray_S30reg_gff_1_SFF_3_n5}), .Q ({new_AGEMA_signal_2692, KeyArray_outS30ser[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3530, KeyArray_S30reg_gff_1_SFF_4_n5}), .Q ({new_AGEMA_signal_2695, KeyArray_outS30ser[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3531, KeyArray_S30reg_gff_1_SFF_5_n5}), .Q ({new_AGEMA_signal_2698, KeyArray_outS30ser[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3532, KeyArray_S30reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_2701, KeyArray_outS30ser[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3533, KeyArray_S30reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_2704, KeyArray_outS30ser[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3347, KeyArray_S31reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_2707, KeyArray_outS31ser[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3348, KeyArray_S31reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_2710, KeyArray_outS31ser[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3349, KeyArray_S31reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_2713, KeyArray_outS31ser[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3350, KeyArray_S31reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_2716, KeyArray_outS31ser[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3351, KeyArray_S31reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_2719, KeyArray_outS31ser[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3352, KeyArray_S31reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_2722, KeyArray_outS31ser[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3353, KeyArray_S31reg_gff_1_SFF_6_n6}), .Q ({new_AGEMA_signal_2725, KeyArray_outS31ser[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3354, KeyArray_S31reg_gff_1_SFF_7_n6}), .Q ({new_AGEMA_signal_2728, KeyArray_outS31ser[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3355, KeyArray_S32reg_gff_1_SFF_0_n6}), .Q ({new_AGEMA_signal_2731, KeyArray_outS32ser[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3356, KeyArray_S32reg_gff_1_SFF_1_n6}), .Q ({new_AGEMA_signal_2734, KeyArray_outS32ser[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3357, KeyArray_S32reg_gff_1_SFF_2_n6}), .Q ({new_AGEMA_signal_2737, KeyArray_outS32ser[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3358, KeyArray_S32reg_gff_1_SFF_3_n6}), .Q ({new_AGEMA_signal_2740, KeyArray_outS32ser[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3359, KeyArray_S32reg_gff_1_SFF_4_n6}), .Q ({new_AGEMA_signal_2743, KeyArray_outS32ser[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3360, KeyArray_S32reg_gff_1_SFF_5_n6}), .Q ({new_AGEMA_signal_2746, KeyArray_outS32ser[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3361, KeyArray_S32reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_2749, KeyArray_outS32ser[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3362, KeyArray_S32reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_2752, KeyArray_outS32ser[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3363, KeyArray_S33reg_gff_1_SFF_0_n5}), .Q ({new_AGEMA_signal_2755, KeyArray_outS33ser[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3364, KeyArray_S33reg_gff_1_SFF_1_n5}), .Q ({new_AGEMA_signal_2758, KeyArray_outS33ser[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3365, KeyArray_S33reg_gff_1_SFF_2_n5}), .Q ({new_AGEMA_signal_2761, KeyArray_outS33ser[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3366, KeyArray_S33reg_gff_1_SFF_3_n5}), .Q ({new_AGEMA_signal_2764, KeyArray_outS33ser[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3367, KeyArray_S33reg_gff_1_SFF_4_n5}), .Q ({new_AGEMA_signal_2767, KeyArray_outS33ser[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3368, KeyArray_S33reg_gff_1_SFF_5_n5}), .Q ({new_AGEMA_signal_2770, KeyArray_outS33ser[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3369, KeyArray_S33reg_gff_1_SFF_6_n5}), .Q ({new_AGEMA_signal_2773, KeyArray_outS33ser[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) KeyArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3370, KeyArray_S33reg_gff_1_SFF_7_n5}), .Q ({new_AGEMA_signal_2776, KeyArray_outS33ser[7]}) ) ;
    DFF_X1 calcRCon_s_current_state_reg_0__FF_FF ( .CK (clk_gated), .D (calcRCon_n51), .Q (calcRCon_s_current_state_0_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_1__FF_FF ( .CK (clk_gated), .D (calcRCon_n50), .Q (calcRCon_s_current_state_1_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_2__FF_FF ( .CK (clk_gated), .D (calcRCon_n49), .Q (calcRCon_s_current_state_2_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_3__FF_FF ( .CK (clk_gated), .D (calcRCon_n48), .Q (calcRCon_s_current_state_3_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_4__FF_FF ( .CK (clk_gated), .D (calcRCon_n47), .Q (calcRCon_s_current_state_4_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_5__FF_FF ( .CK (clk_gated), .D (calcRCon_n46), .Q (calcRCon_s_current_state_5_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_6__FF_FF ( .CK (clk_gated), .D (calcRCon_n45), .Q (calcRCon_s_current_state_6_), .QN () ) ;
    DFF_X1 calcRCon_s_current_state_reg_7__FF_FF ( .CK (clk_gated), .D (calcRCon_n44), .Q (calcRCon_n3), .QN () ) ;
    DFF_X1 nReset_reg_FF_FF ( .CK (clk_gated), .D (n9), .Q (nReset), .QN () ) ;
endmodule
