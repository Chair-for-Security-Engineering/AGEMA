/* modified netlist. Source: module CRAFT in file Designs/CRAFT_round-based/AGEMA/CRAFT.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module CRAFT_HPC2_Pipeline_d1 (plaintext_s0, key_s0, clk, rst, key_s1, plaintext_s1, Fresh, ciphertext_s0, done, ciphertext_s1);
    input [63:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input rst ;
    input [127:0] key_s1 ;
    input [63:0] plaintext_s1 ;
    input [255:0] Fresh ;
    output [63:0] ciphertext_s0 ;
    output done ;
    output [63:0] ciphertext_s1 ;
    wire RoundConstant_4_ ;
    wire RoundConstant_0 ;
    wire done_internal ;
    wire MCInst_XOR_r0_Inst_0_n2 ;
    wire MCInst_XOR_r0_Inst_0_n1 ;
    wire MCInst_XOR_r1_Inst_0_n1 ;
    wire MCInst_XOR_r0_Inst_1_n2 ;
    wire MCInst_XOR_r0_Inst_1_n1 ;
    wire MCInst_XOR_r1_Inst_1_n1 ;
    wire MCInst_XOR_r0_Inst_2_n2 ;
    wire MCInst_XOR_r0_Inst_2_n1 ;
    wire MCInst_XOR_r1_Inst_2_n1 ;
    wire MCInst_XOR_r0_Inst_3_n2 ;
    wire MCInst_XOR_r0_Inst_3_n1 ;
    wire MCInst_XOR_r1_Inst_3_n1 ;
    wire MCInst_XOR_r0_Inst_4_n2 ;
    wire MCInst_XOR_r0_Inst_4_n1 ;
    wire MCInst_XOR_r1_Inst_4_n1 ;
    wire MCInst_XOR_r0_Inst_5_n2 ;
    wire MCInst_XOR_r0_Inst_5_n1 ;
    wire MCInst_XOR_r1_Inst_5_n1 ;
    wire MCInst_XOR_r0_Inst_6_n2 ;
    wire MCInst_XOR_r0_Inst_6_n1 ;
    wire MCInst_XOR_r1_Inst_6_n1 ;
    wire MCInst_XOR_r0_Inst_7_n2 ;
    wire MCInst_XOR_r0_Inst_7_n1 ;
    wire MCInst_XOR_r1_Inst_7_n1 ;
    wire MCInst_XOR_r0_Inst_8_n2 ;
    wire MCInst_XOR_r0_Inst_8_n1 ;
    wire MCInst_XOR_r1_Inst_8_n1 ;
    wire MCInst_XOR_r0_Inst_9_n2 ;
    wire MCInst_XOR_r0_Inst_9_n1 ;
    wire MCInst_XOR_r1_Inst_9_n1 ;
    wire MCInst_XOR_r0_Inst_10_n2 ;
    wire MCInst_XOR_r0_Inst_10_n1 ;
    wire MCInst_XOR_r1_Inst_10_n1 ;
    wire MCInst_XOR_r0_Inst_11_n2 ;
    wire MCInst_XOR_r0_Inst_11_n1 ;
    wire MCInst_XOR_r1_Inst_11_n1 ;
    wire MCInst_XOR_r0_Inst_12_n2 ;
    wire MCInst_XOR_r0_Inst_12_n1 ;
    wire MCInst_XOR_r1_Inst_12_n1 ;
    wire MCInst_XOR_r0_Inst_13_n2 ;
    wire MCInst_XOR_r0_Inst_13_n1 ;
    wire MCInst_XOR_r1_Inst_13_n1 ;
    wire MCInst_XOR_r0_Inst_14_n2 ;
    wire MCInst_XOR_r0_Inst_14_n1 ;
    wire MCInst_XOR_r1_Inst_14_n1 ;
    wire MCInst_XOR_r0_Inst_15_n2 ;
    wire MCInst_XOR_r0_Inst_15_n1 ;
    wire MCInst_XOR_r1_Inst_15_n1 ;
    wire AddKeyXOR1_XORInst_0_0_n1 ;
    wire AddKeyXOR1_XORInst_0_1_n1 ;
    wire AddKeyXOR1_XORInst_0_2_n1 ;
    wire AddKeyXOR1_XORInst_0_3_n1 ;
    wire AddKeyXOR1_XORInst_1_0_n1 ;
    wire AddKeyXOR1_XORInst_1_1_n1 ;
    wire AddKeyXOR1_XORInst_1_2_n1 ;
    wire AddKeyXOR1_XORInst_1_3_n1 ;
    wire AddKeyXOR1_XORInst_2_0_n1 ;
    wire AddKeyXOR1_XORInst_2_1_n1 ;
    wire AddKeyXOR1_XORInst_2_2_n1 ;
    wire AddKeyXOR1_XORInst_2_3_n1 ;
    wire AddKeyXOR1_XORInst_3_0_n1 ;
    wire AddKeyXOR1_XORInst_3_1_n1 ;
    wire AddKeyXOR1_XORInst_3_2_n1 ;
    wire AddKeyXOR1_XORInst_3_3_n1 ;
    wire AddKeyConstXOR_XORInst_0_0_n2 ;
    wire AddKeyConstXOR_XORInst_0_0_n1 ;
    wire AddKeyConstXOR_XORInst_0_1_n2 ;
    wire AddKeyConstXOR_XORInst_0_1_n1 ;
    wire AddKeyConstXOR_XORInst_0_2_n2 ;
    wire AddKeyConstXOR_XORInst_0_2_n1 ;
    wire AddKeyConstXOR_XORInst_0_3_n2 ;
    wire AddKeyConstXOR_XORInst_0_3_n1 ;
    wire AddKeyConstXOR_XORInst_1_0_n2 ;
    wire AddKeyConstXOR_XORInst_1_0_n1 ;
    wire AddKeyConstXOR_XORInst_1_1_n2 ;
    wire AddKeyConstXOR_XORInst_1_1_n1 ;
    wire AddKeyConstXOR_XORInst_1_2_n2 ;
    wire AddKeyConstXOR_XORInst_1_2_n1 ;
    wire AddKeyConstXOR_XORInst_1_3_n2 ;
    wire AddKeyConstXOR_XORInst_1_3_n1 ;
    wire AddKeyXOR2_XORInst_0_0_n1 ;
    wire AddKeyXOR2_XORInst_0_1_n1 ;
    wire AddKeyXOR2_XORInst_0_2_n1 ;
    wire AddKeyXOR2_XORInst_0_3_n1 ;
    wire AddKeyXOR2_XORInst_1_0_n1 ;
    wire AddKeyXOR2_XORInst_1_1_n1 ;
    wire AddKeyXOR2_XORInst_1_2_n1 ;
    wire AddKeyXOR2_XORInst_1_3_n1 ;
    wire AddKeyXOR2_XORInst_2_0_n1 ;
    wire AddKeyXOR2_XORInst_2_1_n1 ;
    wire AddKeyXOR2_XORInst_2_2_n1 ;
    wire AddKeyXOR2_XORInst_2_3_n1 ;
    wire AddKeyXOR2_XORInst_3_0_n1 ;
    wire AddKeyXOR2_XORInst_3_1_n1 ;
    wire AddKeyXOR2_XORInst_3_2_n1 ;
    wire AddKeyXOR2_XORInst_3_3_n1 ;
    wire AddKeyXOR2_XORInst_4_0_n1 ;
    wire AddKeyXOR2_XORInst_4_1_n1 ;
    wire AddKeyXOR2_XORInst_4_2_n1 ;
    wire AddKeyXOR2_XORInst_4_3_n1 ;
    wire AddKeyXOR2_XORInst_5_0_n1 ;
    wire AddKeyXOR2_XORInst_5_1_n1 ;
    wire AddKeyXOR2_XORInst_5_2_n1 ;
    wire AddKeyXOR2_XORInst_5_3_n1 ;
    wire AddKeyXOR2_XORInst_6_0_n1 ;
    wire AddKeyXOR2_XORInst_6_1_n1 ;
    wire AddKeyXOR2_XORInst_6_2_n1 ;
    wire AddKeyXOR2_XORInst_6_3_n1 ;
    wire AddKeyXOR2_XORInst_7_0_n1 ;
    wire AddKeyXOR2_XORInst_7_1_n1 ;
    wire AddKeyXOR2_XORInst_7_2_n1 ;
    wire AddKeyXOR2_XORInst_7_3_n1 ;
    wire AddKeyXOR2_XORInst_8_0_n1 ;
    wire AddKeyXOR2_XORInst_8_1_n1 ;
    wire AddKeyXOR2_XORInst_8_2_n1 ;
    wire AddKeyXOR2_XORInst_8_3_n1 ;
    wire AddKeyXOR2_XORInst_9_0_n1 ;
    wire AddKeyXOR2_XORInst_9_1_n1 ;
    wire AddKeyXOR2_XORInst_9_2_n1 ;
    wire AddKeyXOR2_XORInst_9_3_n1 ;
    wire SubCellInst_SboxInst_0_n15 ;
    wire SubCellInst_SboxInst_0_n14 ;
    wire SubCellInst_SboxInst_0_n13 ;
    wire SubCellInst_SboxInst_0_n12 ;
    wire SubCellInst_SboxInst_0_n11 ;
    wire SubCellInst_SboxInst_0_n10 ;
    wire SubCellInst_SboxInst_0_n9 ;
    wire SubCellInst_SboxInst_0_n8 ;
    wire SubCellInst_SboxInst_0_n7 ;
    wire SubCellInst_SboxInst_0_n6 ;
    wire SubCellInst_SboxInst_0_n5 ;
    wire SubCellInst_SboxInst_0_n4 ;
    wire SubCellInst_SboxInst_0_n3 ;
    wire SubCellInst_SboxInst_0_n2 ;
    wire SubCellInst_SboxInst_0_n1 ;
    wire SubCellInst_SboxInst_1_n15 ;
    wire SubCellInst_SboxInst_1_n14 ;
    wire SubCellInst_SboxInst_1_n13 ;
    wire SubCellInst_SboxInst_1_n12 ;
    wire SubCellInst_SboxInst_1_n11 ;
    wire SubCellInst_SboxInst_1_n10 ;
    wire SubCellInst_SboxInst_1_n9 ;
    wire SubCellInst_SboxInst_1_n8 ;
    wire SubCellInst_SboxInst_1_n7 ;
    wire SubCellInst_SboxInst_1_n6 ;
    wire SubCellInst_SboxInst_1_n5 ;
    wire SubCellInst_SboxInst_1_n4 ;
    wire SubCellInst_SboxInst_1_n3 ;
    wire SubCellInst_SboxInst_1_n2 ;
    wire SubCellInst_SboxInst_1_n1 ;
    wire SubCellInst_SboxInst_2_n15 ;
    wire SubCellInst_SboxInst_2_n14 ;
    wire SubCellInst_SboxInst_2_n13 ;
    wire SubCellInst_SboxInst_2_n12 ;
    wire SubCellInst_SboxInst_2_n11 ;
    wire SubCellInst_SboxInst_2_n10 ;
    wire SubCellInst_SboxInst_2_n9 ;
    wire SubCellInst_SboxInst_2_n8 ;
    wire SubCellInst_SboxInst_2_n7 ;
    wire SubCellInst_SboxInst_2_n6 ;
    wire SubCellInst_SboxInst_2_n5 ;
    wire SubCellInst_SboxInst_2_n4 ;
    wire SubCellInst_SboxInst_2_n3 ;
    wire SubCellInst_SboxInst_2_n2 ;
    wire SubCellInst_SboxInst_2_n1 ;
    wire SubCellInst_SboxInst_3_n15 ;
    wire SubCellInst_SboxInst_3_n14 ;
    wire SubCellInst_SboxInst_3_n13 ;
    wire SubCellInst_SboxInst_3_n12 ;
    wire SubCellInst_SboxInst_3_n11 ;
    wire SubCellInst_SboxInst_3_n10 ;
    wire SubCellInst_SboxInst_3_n9 ;
    wire SubCellInst_SboxInst_3_n8 ;
    wire SubCellInst_SboxInst_3_n7 ;
    wire SubCellInst_SboxInst_3_n6 ;
    wire SubCellInst_SboxInst_3_n5 ;
    wire SubCellInst_SboxInst_3_n4 ;
    wire SubCellInst_SboxInst_3_n3 ;
    wire SubCellInst_SboxInst_3_n2 ;
    wire SubCellInst_SboxInst_3_n1 ;
    wire SubCellInst_SboxInst_4_n15 ;
    wire SubCellInst_SboxInst_4_n14 ;
    wire SubCellInst_SboxInst_4_n13 ;
    wire SubCellInst_SboxInst_4_n12 ;
    wire SubCellInst_SboxInst_4_n11 ;
    wire SubCellInst_SboxInst_4_n10 ;
    wire SubCellInst_SboxInst_4_n9 ;
    wire SubCellInst_SboxInst_4_n8 ;
    wire SubCellInst_SboxInst_4_n7 ;
    wire SubCellInst_SboxInst_4_n6 ;
    wire SubCellInst_SboxInst_4_n5 ;
    wire SubCellInst_SboxInst_4_n4 ;
    wire SubCellInst_SboxInst_4_n3 ;
    wire SubCellInst_SboxInst_4_n2 ;
    wire SubCellInst_SboxInst_4_n1 ;
    wire SubCellInst_SboxInst_5_n15 ;
    wire SubCellInst_SboxInst_5_n14 ;
    wire SubCellInst_SboxInst_5_n13 ;
    wire SubCellInst_SboxInst_5_n12 ;
    wire SubCellInst_SboxInst_5_n11 ;
    wire SubCellInst_SboxInst_5_n10 ;
    wire SubCellInst_SboxInst_5_n9 ;
    wire SubCellInst_SboxInst_5_n8 ;
    wire SubCellInst_SboxInst_5_n7 ;
    wire SubCellInst_SboxInst_5_n6 ;
    wire SubCellInst_SboxInst_5_n5 ;
    wire SubCellInst_SboxInst_5_n4 ;
    wire SubCellInst_SboxInst_5_n3 ;
    wire SubCellInst_SboxInst_5_n2 ;
    wire SubCellInst_SboxInst_5_n1 ;
    wire SubCellInst_SboxInst_6_n15 ;
    wire SubCellInst_SboxInst_6_n14 ;
    wire SubCellInst_SboxInst_6_n13 ;
    wire SubCellInst_SboxInst_6_n12 ;
    wire SubCellInst_SboxInst_6_n11 ;
    wire SubCellInst_SboxInst_6_n10 ;
    wire SubCellInst_SboxInst_6_n9 ;
    wire SubCellInst_SboxInst_6_n8 ;
    wire SubCellInst_SboxInst_6_n7 ;
    wire SubCellInst_SboxInst_6_n6 ;
    wire SubCellInst_SboxInst_6_n5 ;
    wire SubCellInst_SboxInst_6_n4 ;
    wire SubCellInst_SboxInst_6_n3 ;
    wire SubCellInst_SboxInst_6_n2 ;
    wire SubCellInst_SboxInst_6_n1 ;
    wire SubCellInst_SboxInst_7_n15 ;
    wire SubCellInst_SboxInst_7_n14 ;
    wire SubCellInst_SboxInst_7_n13 ;
    wire SubCellInst_SboxInst_7_n12 ;
    wire SubCellInst_SboxInst_7_n11 ;
    wire SubCellInst_SboxInst_7_n10 ;
    wire SubCellInst_SboxInst_7_n9 ;
    wire SubCellInst_SboxInst_7_n8 ;
    wire SubCellInst_SboxInst_7_n7 ;
    wire SubCellInst_SboxInst_7_n6 ;
    wire SubCellInst_SboxInst_7_n5 ;
    wire SubCellInst_SboxInst_7_n4 ;
    wire SubCellInst_SboxInst_7_n3 ;
    wire SubCellInst_SboxInst_7_n2 ;
    wire SubCellInst_SboxInst_7_n1 ;
    wire SubCellInst_SboxInst_8_n15 ;
    wire SubCellInst_SboxInst_8_n14 ;
    wire SubCellInst_SboxInst_8_n13 ;
    wire SubCellInst_SboxInst_8_n12 ;
    wire SubCellInst_SboxInst_8_n11 ;
    wire SubCellInst_SboxInst_8_n10 ;
    wire SubCellInst_SboxInst_8_n9 ;
    wire SubCellInst_SboxInst_8_n8 ;
    wire SubCellInst_SboxInst_8_n7 ;
    wire SubCellInst_SboxInst_8_n6 ;
    wire SubCellInst_SboxInst_8_n5 ;
    wire SubCellInst_SboxInst_8_n4 ;
    wire SubCellInst_SboxInst_8_n3 ;
    wire SubCellInst_SboxInst_8_n2 ;
    wire SubCellInst_SboxInst_8_n1 ;
    wire SubCellInst_SboxInst_9_n15 ;
    wire SubCellInst_SboxInst_9_n14 ;
    wire SubCellInst_SboxInst_9_n13 ;
    wire SubCellInst_SboxInst_9_n12 ;
    wire SubCellInst_SboxInst_9_n11 ;
    wire SubCellInst_SboxInst_9_n10 ;
    wire SubCellInst_SboxInst_9_n9 ;
    wire SubCellInst_SboxInst_9_n8 ;
    wire SubCellInst_SboxInst_9_n7 ;
    wire SubCellInst_SboxInst_9_n6 ;
    wire SubCellInst_SboxInst_9_n5 ;
    wire SubCellInst_SboxInst_9_n4 ;
    wire SubCellInst_SboxInst_9_n3 ;
    wire SubCellInst_SboxInst_9_n2 ;
    wire SubCellInst_SboxInst_9_n1 ;
    wire SubCellInst_SboxInst_10_n15 ;
    wire SubCellInst_SboxInst_10_n14 ;
    wire SubCellInst_SboxInst_10_n13 ;
    wire SubCellInst_SboxInst_10_n12 ;
    wire SubCellInst_SboxInst_10_n11 ;
    wire SubCellInst_SboxInst_10_n10 ;
    wire SubCellInst_SboxInst_10_n9 ;
    wire SubCellInst_SboxInst_10_n8 ;
    wire SubCellInst_SboxInst_10_n7 ;
    wire SubCellInst_SboxInst_10_n6 ;
    wire SubCellInst_SboxInst_10_n5 ;
    wire SubCellInst_SboxInst_10_n4 ;
    wire SubCellInst_SboxInst_10_n3 ;
    wire SubCellInst_SboxInst_10_n2 ;
    wire SubCellInst_SboxInst_10_n1 ;
    wire SubCellInst_SboxInst_11_n15 ;
    wire SubCellInst_SboxInst_11_n14 ;
    wire SubCellInst_SboxInst_11_n13 ;
    wire SubCellInst_SboxInst_11_n12 ;
    wire SubCellInst_SboxInst_11_n11 ;
    wire SubCellInst_SboxInst_11_n10 ;
    wire SubCellInst_SboxInst_11_n9 ;
    wire SubCellInst_SboxInst_11_n8 ;
    wire SubCellInst_SboxInst_11_n7 ;
    wire SubCellInst_SboxInst_11_n6 ;
    wire SubCellInst_SboxInst_11_n5 ;
    wire SubCellInst_SboxInst_11_n4 ;
    wire SubCellInst_SboxInst_11_n3 ;
    wire SubCellInst_SboxInst_11_n2 ;
    wire SubCellInst_SboxInst_11_n1 ;
    wire SubCellInst_SboxInst_12_n15 ;
    wire SubCellInst_SboxInst_12_n14 ;
    wire SubCellInst_SboxInst_12_n13 ;
    wire SubCellInst_SboxInst_12_n12 ;
    wire SubCellInst_SboxInst_12_n11 ;
    wire SubCellInst_SboxInst_12_n10 ;
    wire SubCellInst_SboxInst_12_n9 ;
    wire SubCellInst_SboxInst_12_n8 ;
    wire SubCellInst_SboxInst_12_n7 ;
    wire SubCellInst_SboxInst_12_n6 ;
    wire SubCellInst_SboxInst_12_n5 ;
    wire SubCellInst_SboxInst_12_n4 ;
    wire SubCellInst_SboxInst_12_n3 ;
    wire SubCellInst_SboxInst_12_n2 ;
    wire SubCellInst_SboxInst_12_n1 ;
    wire SubCellInst_SboxInst_13_n15 ;
    wire SubCellInst_SboxInst_13_n14 ;
    wire SubCellInst_SboxInst_13_n13 ;
    wire SubCellInst_SboxInst_13_n12 ;
    wire SubCellInst_SboxInst_13_n11 ;
    wire SubCellInst_SboxInst_13_n10 ;
    wire SubCellInst_SboxInst_13_n9 ;
    wire SubCellInst_SboxInst_13_n8 ;
    wire SubCellInst_SboxInst_13_n7 ;
    wire SubCellInst_SboxInst_13_n6 ;
    wire SubCellInst_SboxInst_13_n5 ;
    wire SubCellInst_SboxInst_13_n4 ;
    wire SubCellInst_SboxInst_13_n3 ;
    wire SubCellInst_SboxInst_13_n2 ;
    wire SubCellInst_SboxInst_13_n1 ;
    wire SubCellInst_SboxInst_14_n15 ;
    wire SubCellInst_SboxInst_14_n14 ;
    wire SubCellInst_SboxInst_14_n13 ;
    wire SubCellInst_SboxInst_14_n12 ;
    wire SubCellInst_SboxInst_14_n11 ;
    wire SubCellInst_SboxInst_14_n10 ;
    wire SubCellInst_SboxInst_14_n9 ;
    wire SubCellInst_SboxInst_14_n8 ;
    wire SubCellInst_SboxInst_14_n7 ;
    wire SubCellInst_SboxInst_14_n6 ;
    wire SubCellInst_SboxInst_14_n5 ;
    wire SubCellInst_SboxInst_14_n4 ;
    wire SubCellInst_SboxInst_14_n3 ;
    wire SubCellInst_SboxInst_14_n2 ;
    wire SubCellInst_SboxInst_14_n1 ;
    wire SubCellInst_SboxInst_15_n15 ;
    wire SubCellInst_SboxInst_15_n14 ;
    wire SubCellInst_SboxInst_15_n13 ;
    wire SubCellInst_SboxInst_15_n12 ;
    wire SubCellInst_SboxInst_15_n11 ;
    wire SubCellInst_SboxInst_15_n10 ;
    wire SubCellInst_SboxInst_15_n9 ;
    wire SubCellInst_SboxInst_15_n8 ;
    wire SubCellInst_SboxInst_15_n7 ;
    wire SubCellInst_SboxInst_15_n6 ;
    wire SubCellInst_SboxInst_15_n5 ;
    wire SubCellInst_SboxInst_15_n4 ;
    wire SubCellInst_SboxInst_15_n3 ;
    wire SubCellInst_SboxInst_15_n2 ;
    wire SubCellInst_SboxInst_15_n1 ;
    wire KeyMUX_n9 ;
    wire KeyMUX_n8 ;
    wire KeyMUX_n7 ;
    wire FSMSignalsInst_n5 ;
    wire FSMSignalsInst_n4 ;
    wire FSMSignalsInst_n3 ;
    wire FSMSignalsInst_n2 ;
    wire FSMSignalsInst_n1 ;
    wire selectsUpdateInst_n3 ;
    wire [63:0] Feedback ;
    wire [63:32] MCInput ;
    wire [63:0] MCOutput ;
    wire [63:0] SelectedKey ;
    wire [63:0] AddRoundKeyOutput ;
    wire [1:0] selects ;
    wire [6:0] FSMReg ;
    wire [6:0] FSMUpdate ;
    wire [1:0] selectsReg ;
    wire [1:0] selectsNext ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;

    /* cells in depth 0 */
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_1524, SelectedKey[40]}), .b ({1'b0, RoundConstant_0}), .c ({new_AGEMA_signal_1707, AddKeyConstXOR_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_1527, SelectedKey[41]}), .b ({1'b0, FSMUpdate[0]}), .c ({new_AGEMA_signal_1708, AddKeyConstXOR_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_1530, SelectedKey[42]}), .b ({1'b0, FSMUpdate[1]}), .c ({new_AGEMA_signal_1709, AddKeyConstXOR_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_1533, SelectedKey[43]}), .b ({1'b0, 1'b0}), .c ({new_AGEMA_signal_1710, AddKeyConstXOR_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_1536, SelectedKey[44]}), .b ({1'b0, RoundConstant_4_}), .c ({new_AGEMA_signal_1711, AddKeyConstXOR_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_1539, SelectedKey[45]}), .b ({1'b0, FSMUpdate[3]}), .c ({new_AGEMA_signal_1712, AddKeyConstXOR_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_1542, SelectedKey[46]}), .b ({1'b0, FSMUpdate[4]}), .c ({new_AGEMA_signal_1713, AddKeyConstXOR_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_1545, SelectedKey[47]}), .b ({1'b0, FSMUpdate[5]}), .c ({new_AGEMA_signal_1714, AddKeyConstXOR_XORInst_1_3_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U4 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_1024, SubCellInst_SboxInst_0_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U2 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_1025, SubCellInst_SboxInst_0_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U1 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_1026, SubCellInst_SboxInst_0_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U4 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_1032, SubCellInst_SboxInst_1_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U2 ( .a ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({new_AGEMA_signal_1033, SubCellInst_SboxInst_1_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U1 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_1034, SubCellInst_SboxInst_1_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U4 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({new_AGEMA_signal_1040, SubCellInst_SboxInst_2_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U2 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({new_AGEMA_signal_1041, SubCellInst_SboxInst_2_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U1 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_1042, SubCellInst_SboxInst_2_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U4 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_1048, SubCellInst_SboxInst_3_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U2 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_1049, SubCellInst_SboxInst_3_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U1 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_1050, SubCellInst_SboxInst_3_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U4 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_1056, SubCellInst_SboxInst_4_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U2 ( .a ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({new_AGEMA_signal_1057, SubCellInst_SboxInst_4_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U1 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_1058, SubCellInst_SboxInst_4_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U4 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({new_AGEMA_signal_1064, SubCellInst_SboxInst_5_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U2 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({new_AGEMA_signal_1065, SubCellInst_SboxInst_5_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U1 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_1066, SubCellInst_SboxInst_5_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U4 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_1072, SubCellInst_SboxInst_6_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U2 ( .a ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({new_AGEMA_signal_1073, SubCellInst_SboxInst_6_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U1 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_1074, SubCellInst_SboxInst_6_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U4 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({new_AGEMA_signal_1080, SubCellInst_SboxInst_7_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U2 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({new_AGEMA_signal_1081, SubCellInst_SboxInst_7_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U1 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_1082, SubCellInst_SboxInst_7_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U4 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_1088, SubCellInst_SboxInst_8_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U2 ( .a ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({new_AGEMA_signal_1089, SubCellInst_SboxInst_8_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U1 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_1090, SubCellInst_SboxInst_8_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U4 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_1096, SubCellInst_SboxInst_9_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U2 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_1097, SubCellInst_SboxInst_9_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U1 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_1098, SubCellInst_SboxInst_9_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U4 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_1104, SubCellInst_SboxInst_10_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U2 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_1105, SubCellInst_SboxInst_10_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U1 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_1106, SubCellInst_SboxInst_10_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U4 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({new_AGEMA_signal_1112, SubCellInst_SboxInst_11_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U2 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({new_AGEMA_signal_1113, SubCellInst_SboxInst_11_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U1 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_1114, SubCellInst_SboxInst_11_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U4 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({new_AGEMA_signal_1120, SubCellInst_SboxInst_12_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U2 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({new_AGEMA_signal_1121, SubCellInst_SboxInst_12_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U1 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_1122, SubCellInst_SboxInst_12_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U4 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_1128, SubCellInst_SboxInst_13_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U2 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({new_AGEMA_signal_1129, SubCellInst_SboxInst_13_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U1 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_1130, SubCellInst_SboxInst_13_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U4 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({new_AGEMA_signal_1136, SubCellInst_SboxInst_14_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U2 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({new_AGEMA_signal_1137, SubCellInst_SboxInst_14_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U1 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_1138, SubCellInst_SboxInst_14_n9}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U4 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_1144, SubCellInst_SboxInst_15_n7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U2 ( .a ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({new_AGEMA_signal_1145, SubCellInst_SboxInst_15_n8}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U1 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_1146, SubCellInst_SboxInst_15_n9}) ) ;
    INV_X1 KeyMUX_U3 ( .A (selects[0]), .ZN (KeyMUX_n9) ) ;
    INV_X1 KeyMUX_U2 ( .A (KeyMUX_n9), .ZN (KeyMUX_n8) ) ;
    INV_X1 KeyMUX_U1 ( .A (KeyMUX_n9), .ZN (KeyMUX_n7) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_0_U1 ( .s (selects[0]), .b ({key_s1[64], key_s0[64]}), .a ({key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_1245, SelectedKey[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_1_U1 ( .s (KeyMUX_n8), .b ({key_s1[65], key_s0[65]}), .a ({key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_1437, SelectedKey[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_2_U1 ( .s (selects[0]), .b ({key_s1[66], key_s0[66]}), .a ({key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_1248, SelectedKey[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_3_U1 ( .s (KeyMUX_n8), .b ({key_s1[67], key_s0[67]}), .a ({key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_1440, SelectedKey[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_4_U1 ( .s (KeyMUX_n8), .b ({key_s1[68], key_s0[68]}), .a ({key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_1443, SelectedKey[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_5_U1 ( .s (KeyMUX_n8), .b ({key_s1[69], key_s0[69]}), .a ({key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_1446, SelectedKey[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_6_U1 ( .s (KeyMUX_n8), .b ({key_s1[70], key_s0[70]}), .a ({key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_1449, SelectedKey[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_7_U1 ( .s (KeyMUX_n8), .b ({key_s1[71], key_s0[71]}), .a ({key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_1452, SelectedKey[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_8_U1 ( .s (KeyMUX_n8), .b ({key_s1[72], key_s0[72]}), .a ({key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_1455, SelectedKey[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_9_U1 ( .s (KeyMUX_n8), .b ({key_s1[73], key_s0[73]}), .a ({key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_1458, SelectedKey[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_10_U1 ( .s (KeyMUX_n8), .b ({key_s1[74], key_s0[74]}), .a ({key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_1461, SelectedKey[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_11_U1 ( .s (KeyMUX_n8), .b ({key_s1[75], key_s0[75]}), .a ({key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_1464, SelectedKey[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_12_U1 ( .s (KeyMUX_n8), .b ({key_s1[76], key_s0[76]}), .a ({key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_1467, SelectedKey[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_13_U1 ( .s (KeyMUX_n8), .b ({key_s1[77], key_s0[77]}), .a ({key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_1470, SelectedKey[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_14_U1 ( .s (KeyMUX_n8), .b ({key_s1[78], key_s0[78]}), .a ({key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_1473, SelectedKey[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_15_U1 ( .s (KeyMUX_n8), .b ({key_s1[79], key_s0[79]}), .a ({key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_1476, SelectedKey[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_16_U1 ( .s (KeyMUX_n8), .b ({key_s1[80], key_s0[80]}), .a ({key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_1479, SelectedKey[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_17_U1 ( .s (KeyMUX_n8), .b ({key_s1[81], key_s0[81]}), .a ({key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_1482, SelectedKey[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_18_U1 ( .s (KeyMUX_n8), .b ({key_s1[82], key_s0[82]}), .a ({key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_1485, SelectedKey[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_19_U1 ( .s (KeyMUX_n8), .b ({key_s1[83], key_s0[83]}), .a ({key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_1488, SelectedKey[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_20_U1 ( .s (KeyMUX_n8), .b ({key_s1[84], key_s0[84]}), .a ({key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_1491, SelectedKey[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_21_U1 ( .s (KeyMUX_n8), .b ({key_s1[85], key_s0[85]}), .a ({key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_1494, SelectedKey[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_22_U1 ( .s (selects[0]), .b ({key_s1[86], key_s0[86]}), .a ({key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_1251, SelectedKey[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_23_U1 ( .s (selects[0]), .b ({key_s1[87], key_s0[87]}), .a ({key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_1254, SelectedKey[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_24_U1 ( .s (selects[0]), .b ({key_s1[88], key_s0[88]}), .a ({key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_1257, SelectedKey[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_25_U1 ( .s (selects[0]), .b ({key_s1[89], key_s0[89]}), .a ({key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_1260, SelectedKey[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_26_U1 ( .s (selects[0]), .b ({key_s1[90], key_s0[90]}), .a ({key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_1263, SelectedKey[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_27_U1 ( .s (selects[0]), .b ({key_s1[91], key_s0[91]}), .a ({key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_1266, SelectedKey[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_28_U1 ( .s (KeyMUX_n7), .b ({key_s1[92], key_s0[92]}), .a ({key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_1497, SelectedKey[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_29_U1 ( .s (KeyMUX_n7), .b ({key_s1[93], key_s0[93]}), .a ({key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_1500, SelectedKey[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_30_U1 ( .s (KeyMUX_n7), .b ({key_s1[94], key_s0[94]}), .a ({key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_1503, SelectedKey[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_31_U1 ( .s (KeyMUX_n7), .b ({key_s1[95], key_s0[95]}), .a ({key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_1506, SelectedKey[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_32_U1 ( .s (KeyMUX_n7), .b ({key_s1[96], key_s0[96]}), .a ({key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_1509, SelectedKey[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_33_U1 ( .s (selects[0]), .b ({key_s1[97], key_s0[97]}), .a ({key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_1269, SelectedKey[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_34_U1 ( .s (KeyMUX_n7), .b ({key_s1[98], key_s0[98]}), .a ({key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_1512, SelectedKey[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_35_U1 ( .s (KeyMUX_n7), .b ({key_s1[99], key_s0[99]}), .a ({key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_1515, SelectedKey[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_36_U1 ( .s (selects[0]), .b ({key_s1[100], key_s0[100]}), .a ({key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_1272, SelectedKey[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_37_U1 ( .s (KeyMUX_n7), .b ({key_s1[101], key_s0[101]}), .a ({key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_1518, SelectedKey[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_38_U1 ( .s (KeyMUX_n7), .b ({key_s1[102], key_s0[102]}), .a ({key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_1521, SelectedKey[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_39_U1 ( .s (selects[0]), .b ({key_s1[103], key_s0[103]}), .a ({key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_1275, SelectedKey[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_40_U1 ( .s (KeyMUX_n7), .b ({key_s1[104], key_s0[104]}), .a ({key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_1524, SelectedKey[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_41_U1 ( .s (KeyMUX_n7), .b ({key_s1[105], key_s0[105]}), .a ({key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_1527, SelectedKey[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_42_U1 ( .s (KeyMUX_n7), .b ({key_s1[106], key_s0[106]}), .a ({key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_1530, SelectedKey[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_43_U1 ( .s (KeyMUX_n7), .b ({key_s1[107], key_s0[107]}), .a ({key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_1533, SelectedKey[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_44_U1 ( .s (KeyMUX_n7), .b ({key_s1[108], key_s0[108]}), .a ({key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_1536, SelectedKey[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_45_U1 ( .s (KeyMUX_n7), .b ({key_s1[109], key_s0[109]}), .a ({key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_1539, SelectedKey[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_46_U1 ( .s (KeyMUX_n7), .b ({key_s1[110], key_s0[110]}), .a ({key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_1542, SelectedKey[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_47_U1 ( .s (KeyMUX_n7), .b ({key_s1[111], key_s0[111]}), .a ({key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_1545, SelectedKey[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_48_U1 ( .s (KeyMUX_n7), .b ({key_s1[112], key_s0[112]}), .a ({key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_1548, SelectedKey[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_49_U1 ( .s (KeyMUX_n7), .b ({key_s1[113], key_s0[113]}), .a ({key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_1551, SelectedKey[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_50_U1 ( .s (KeyMUX_n7), .b ({key_s1[114], key_s0[114]}), .a ({key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_1554, SelectedKey[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_51_U1 ( .s (KeyMUX_n7), .b ({key_s1[115], key_s0[115]}), .a ({key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_1557, SelectedKey[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_52_U1 ( .s (KeyMUX_n7), .b ({key_s1[116], key_s0[116]}), .a ({key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_1560, SelectedKey[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_53_U1 ( .s (selects[0]), .b ({key_s1[117], key_s0[117]}), .a ({key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_1278, SelectedKey[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_54_U1 ( .s (selects[0]), .b ({key_s1[118], key_s0[118]}), .a ({key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_1281, SelectedKey[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_55_U1 ( .s (KeyMUX_n7), .b ({key_s1[119], key_s0[119]}), .a ({key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_1563, SelectedKey[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_56_U1 ( .s (selects[0]), .b ({key_s1[120], key_s0[120]}), .a ({key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_1284, SelectedKey[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_57_U1 ( .s (KeyMUX_n7), .b ({key_s1[121], key_s0[121]}), .a ({key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_1566, SelectedKey[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_58_U1 ( .s (KeyMUX_n7), .b ({key_s1[122], key_s0[122]}), .a ({key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_1569, SelectedKey[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_59_U1 ( .s (selects[0]), .b ({key_s1[123], key_s0[123]}), .a ({key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_1287, SelectedKey[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_60_U1 ( .s (KeyMUX_n7), .b ({key_s1[124], key_s0[124]}), .a ({key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_1572, SelectedKey[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_61_U1 ( .s (KeyMUX_n7), .b ({key_s1[125], key_s0[125]}), .a ({key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_1575, SelectedKey[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_62_U1 ( .s (selects[0]), .b ({key_s1[126], key_s0[126]}), .a ({key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_1290, SelectedKey[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyMUX_MUXInst_63_U1 ( .s (KeyMUX_n7), .b ({key_s1[127], key_s0[127]}), .a ({key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_1578, SelectedKey[63]}) ) ;
    MUX2_X1 FSMMUX_MUXInst_0_U1 ( .S (rst), .A (FSMReg[0]), .B (1'b1), .Z (RoundConstant_0) ) ;
    MUX2_X1 FSMMUX_MUXInst_1_U1 ( .S (rst), .A (FSMReg[1]), .B (1'b0), .Z (FSMUpdate[0]) ) ;
    MUX2_X1 FSMMUX_MUXInst_2_U1 ( .S (rst), .A (FSMReg[2]), .B (1'b0), .Z (FSMUpdate[1]) ) ;
    MUX2_X1 FSMMUX_MUXInst_3_U1 ( .S (rst), .A (FSMReg[3]), .B (1'b1), .Z (RoundConstant_4_) ) ;
    MUX2_X1 FSMMUX_MUXInst_4_U1 ( .S (rst), .A (FSMReg[4]), .B (1'b0), .Z (FSMUpdate[3]) ) ;
    MUX2_X1 FSMMUX_MUXInst_5_U1 ( .S (rst), .A (FSMReg[5]), .B (1'b0), .Z (FSMUpdate[4]) ) ;
    MUX2_X1 FSMMUX_MUXInst_6_U1 ( .S (rst), .A (FSMReg[6]), .B (1'b0), .Z (FSMUpdate[5]) ) ;
    XOR2_X1 FSMUpdateInst_U2 ( .A (RoundConstant_4_), .B (FSMUpdate[3]), .Z (FSMUpdate[6]) ) ;
    XOR2_X1 FSMUpdateInst_U1 ( .A (FSMUpdate[0]), .B (RoundConstant_0), .Z (FSMUpdate[2]) ) ;
    AND2_X1 FSMSignalsInst_U6 ( .A1 (FSMUpdate[5]), .A2 (FSMSignalsInst_n5), .ZN (done_internal) ) ;
    NOR2_X1 FSMSignalsInst_U5 ( .A1 (FSMSignalsInst_n4), .A2 (FSMSignalsInst_n3), .ZN (FSMSignalsInst_n5) ) ;
    NAND2_X1 FSMSignalsInst_U4 ( .A1 (FSMSignalsInst_n2), .A2 (FSMSignalsInst_n1), .ZN (FSMSignalsInst_n3) ) ;
    NOR2_X1 FSMSignalsInst_U3 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdate[4]), .ZN (FSMSignalsInst_n1) ) ;
    NOR2_X1 FSMSignalsInst_U2 ( .A1 (FSMUpdate[0]), .A2 (RoundConstant_4_), .ZN (FSMSignalsInst_n2) ) ;
    NAND2_X1 FSMSignalsInst_U1 ( .A1 (RoundConstant_0), .A2 (FSMUpdate[1]), .ZN (FSMSignalsInst_n4) ) ;
    MUX2_X1 selectsMUX_MUXInst_0_U1 ( .S (rst), .A (selectsReg[0]), .B (1'b0), .Z (selects[0]) ) ;
    MUX2_X1 selectsMUX_MUXInst_1_U1 ( .S (rst), .A (selectsReg[1]), .B (1'b0), .Z (selects[1]) ) ;
    XNOR2_X1 selectsUpdateInst_U3 ( .A (selectsUpdateInst_n3), .B (selects[1]), .ZN (selectsNext[1]) ) ;
    XNOR2_X1 selectsUpdateInst_U2 ( .A (selects[0]), .B (1'b0), .ZN (selectsUpdateInst_n3) ) ;
    INV_X1 selectsUpdateInst_U1 ( .A (selects[0]), .ZN (selectsNext[0]) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_819 ( .C (clk), .D (ciphertext_s0[61]), .Q (new_AGEMA_signal_2179) ) ;
    buf_clk new_AGEMA_reg_buffer_821 ( .C (clk), .D (ciphertext_s1[61]), .Q (new_AGEMA_signal_2181) ) ;
    buf_clk new_AGEMA_reg_buffer_823 ( .C (clk), .D (SubCellInst_SboxInst_0_n9), .Q (new_AGEMA_signal_2183) ) ;
    buf_clk new_AGEMA_reg_buffer_825 ( .C (clk), .D (new_AGEMA_signal_1026), .Q (new_AGEMA_signal_2185) ) ;
    buf_clk new_AGEMA_reg_buffer_827 ( .C (clk), .D (ciphertext_s0[60]), .Q (new_AGEMA_signal_2187) ) ;
    buf_clk new_AGEMA_reg_buffer_829 ( .C (clk), .D (ciphertext_s1[60]), .Q (new_AGEMA_signal_2189) ) ;
    buf_clk new_AGEMA_reg_buffer_831 ( .C (clk), .D (SubCellInst_SboxInst_0_n7), .Q (new_AGEMA_signal_2191) ) ;
    buf_clk new_AGEMA_reg_buffer_833 ( .C (clk), .D (new_AGEMA_signal_1024), .Q (new_AGEMA_signal_2193) ) ;
    buf_clk new_AGEMA_reg_buffer_835 ( .C (clk), .D (ciphertext_s0[49]), .Q (new_AGEMA_signal_2195) ) ;
    buf_clk new_AGEMA_reg_buffer_837 ( .C (clk), .D (ciphertext_s1[49]), .Q (new_AGEMA_signal_2197) ) ;
    buf_clk new_AGEMA_reg_buffer_839 ( .C (clk), .D (SubCellInst_SboxInst_1_n9), .Q (new_AGEMA_signal_2199) ) ;
    buf_clk new_AGEMA_reg_buffer_841 ( .C (clk), .D (new_AGEMA_signal_1034), .Q (new_AGEMA_signal_2201) ) ;
    buf_clk new_AGEMA_reg_buffer_843 ( .C (clk), .D (ciphertext_s0[48]), .Q (new_AGEMA_signal_2203) ) ;
    buf_clk new_AGEMA_reg_buffer_845 ( .C (clk), .D (ciphertext_s1[48]), .Q (new_AGEMA_signal_2205) ) ;
    buf_clk new_AGEMA_reg_buffer_847 ( .C (clk), .D (SubCellInst_SboxInst_1_n7), .Q (new_AGEMA_signal_2207) ) ;
    buf_clk new_AGEMA_reg_buffer_849 ( .C (clk), .D (new_AGEMA_signal_1032), .Q (new_AGEMA_signal_2209) ) ;
    buf_clk new_AGEMA_reg_buffer_851 ( .C (clk), .D (ciphertext_s0[53]), .Q (new_AGEMA_signal_2211) ) ;
    buf_clk new_AGEMA_reg_buffer_853 ( .C (clk), .D (ciphertext_s1[53]), .Q (new_AGEMA_signal_2213) ) ;
    buf_clk new_AGEMA_reg_buffer_855 ( .C (clk), .D (SubCellInst_SboxInst_2_n9), .Q (new_AGEMA_signal_2215) ) ;
    buf_clk new_AGEMA_reg_buffer_857 ( .C (clk), .D (new_AGEMA_signal_1042), .Q (new_AGEMA_signal_2217) ) ;
    buf_clk new_AGEMA_reg_buffer_859 ( .C (clk), .D (ciphertext_s0[52]), .Q (new_AGEMA_signal_2219) ) ;
    buf_clk new_AGEMA_reg_buffer_861 ( .C (clk), .D (ciphertext_s1[52]), .Q (new_AGEMA_signal_2221) ) ;
    buf_clk new_AGEMA_reg_buffer_863 ( .C (clk), .D (SubCellInst_SboxInst_2_n7), .Q (new_AGEMA_signal_2223) ) ;
    buf_clk new_AGEMA_reg_buffer_865 ( .C (clk), .D (new_AGEMA_signal_1040), .Q (new_AGEMA_signal_2225) ) ;
    buf_clk new_AGEMA_reg_buffer_867 ( .C (clk), .D (ciphertext_s0[57]), .Q (new_AGEMA_signal_2227) ) ;
    buf_clk new_AGEMA_reg_buffer_869 ( .C (clk), .D (ciphertext_s1[57]), .Q (new_AGEMA_signal_2229) ) ;
    buf_clk new_AGEMA_reg_buffer_871 ( .C (clk), .D (SubCellInst_SboxInst_3_n9), .Q (new_AGEMA_signal_2231) ) ;
    buf_clk new_AGEMA_reg_buffer_873 ( .C (clk), .D (new_AGEMA_signal_1050), .Q (new_AGEMA_signal_2233) ) ;
    buf_clk new_AGEMA_reg_buffer_875 ( .C (clk), .D (ciphertext_s0[56]), .Q (new_AGEMA_signal_2235) ) ;
    buf_clk new_AGEMA_reg_buffer_877 ( .C (clk), .D (ciphertext_s1[56]), .Q (new_AGEMA_signal_2237) ) ;
    buf_clk new_AGEMA_reg_buffer_879 ( .C (clk), .D (SubCellInst_SboxInst_3_n7), .Q (new_AGEMA_signal_2239) ) ;
    buf_clk new_AGEMA_reg_buffer_881 ( .C (clk), .D (new_AGEMA_signal_1048), .Q (new_AGEMA_signal_2241) ) ;
    buf_clk new_AGEMA_reg_buffer_883 ( .C (clk), .D (ciphertext_s0[33]), .Q (new_AGEMA_signal_2243) ) ;
    buf_clk new_AGEMA_reg_buffer_885 ( .C (clk), .D (ciphertext_s1[33]), .Q (new_AGEMA_signal_2245) ) ;
    buf_clk new_AGEMA_reg_buffer_887 ( .C (clk), .D (SubCellInst_SboxInst_4_n9), .Q (new_AGEMA_signal_2247) ) ;
    buf_clk new_AGEMA_reg_buffer_889 ( .C (clk), .D (new_AGEMA_signal_1058), .Q (new_AGEMA_signal_2249) ) ;
    buf_clk new_AGEMA_reg_buffer_891 ( .C (clk), .D (ciphertext_s0[32]), .Q (new_AGEMA_signal_2251) ) ;
    buf_clk new_AGEMA_reg_buffer_893 ( .C (clk), .D (ciphertext_s1[32]), .Q (new_AGEMA_signal_2253) ) ;
    buf_clk new_AGEMA_reg_buffer_895 ( .C (clk), .D (SubCellInst_SboxInst_4_n7), .Q (new_AGEMA_signal_2255) ) ;
    buf_clk new_AGEMA_reg_buffer_897 ( .C (clk), .D (new_AGEMA_signal_1056), .Q (new_AGEMA_signal_2257) ) ;
    buf_clk new_AGEMA_reg_buffer_899 ( .C (clk), .D (ciphertext_s0[45]), .Q (new_AGEMA_signal_2259) ) ;
    buf_clk new_AGEMA_reg_buffer_901 ( .C (clk), .D (ciphertext_s1[45]), .Q (new_AGEMA_signal_2261) ) ;
    buf_clk new_AGEMA_reg_buffer_903 ( .C (clk), .D (SubCellInst_SboxInst_5_n9), .Q (new_AGEMA_signal_2263) ) ;
    buf_clk new_AGEMA_reg_buffer_905 ( .C (clk), .D (new_AGEMA_signal_1066), .Q (new_AGEMA_signal_2265) ) ;
    buf_clk new_AGEMA_reg_buffer_907 ( .C (clk), .D (ciphertext_s0[44]), .Q (new_AGEMA_signal_2267) ) ;
    buf_clk new_AGEMA_reg_buffer_909 ( .C (clk), .D (ciphertext_s1[44]), .Q (new_AGEMA_signal_2269) ) ;
    buf_clk new_AGEMA_reg_buffer_911 ( .C (clk), .D (SubCellInst_SboxInst_5_n7), .Q (new_AGEMA_signal_2271) ) ;
    buf_clk new_AGEMA_reg_buffer_913 ( .C (clk), .D (new_AGEMA_signal_1064), .Q (new_AGEMA_signal_2273) ) ;
    buf_clk new_AGEMA_reg_buffer_915 ( .C (clk), .D (ciphertext_s0[41]), .Q (new_AGEMA_signal_2275) ) ;
    buf_clk new_AGEMA_reg_buffer_917 ( .C (clk), .D (ciphertext_s1[41]), .Q (new_AGEMA_signal_2277) ) ;
    buf_clk new_AGEMA_reg_buffer_919 ( .C (clk), .D (SubCellInst_SboxInst_6_n9), .Q (new_AGEMA_signal_2279) ) ;
    buf_clk new_AGEMA_reg_buffer_921 ( .C (clk), .D (new_AGEMA_signal_1074), .Q (new_AGEMA_signal_2281) ) ;
    buf_clk new_AGEMA_reg_buffer_923 ( .C (clk), .D (ciphertext_s0[40]), .Q (new_AGEMA_signal_2283) ) ;
    buf_clk new_AGEMA_reg_buffer_925 ( .C (clk), .D (ciphertext_s1[40]), .Q (new_AGEMA_signal_2285) ) ;
    buf_clk new_AGEMA_reg_buffer_927 ( .C (clk), .D (SubCellInst_SboxInst_6_n7), .Q (new_AGEMA_signal_2287) ) ;
    buf_clk new_AGEMA_reg_buffer_929 ( .C (clk), .D (new_AGEMA_signal_1072), .Q (new_AGEMA_signal_2289) ) ;
    buf_clk new_AGEMA_reg_buffer_931 ( .C (clk), .D (ciphertext_s0[37]), .Q (new_AGEMA_signal_2291) ) ;
    buf_clk new_AGEMA_reg_buffer_933 ( .C (clk), .D (ciphertext_s1[37]), .Q (new_AGEMA_signal_2293) ) ;
    buf_clk new_AGEMA_reg_buffer_935 ( .C (clk), .D (SubCellInst_SboxInst_7_n9), .Q (new_AGEMA_signal_2295) ) ;
    buf_clk new_AGEMA_reg_buffer_937 ( .C (clk), .D (new_AGEMA_signal_1082), .Q (new_AGEMA_signal_2297) ) ;
    buf_clk new_AGEMA_reg_buffer_939 ( .C (clk), .D (ciphertext_s0[36]), .Q (new_AGEMA_signal_2299) ) ;
    buf_clk new_AGEMA_reg_buffer_941 ( .C (clk), .D (ciphertext_s1[36]), .Q (new_AGEMA_signal_2301) ) ;
    buf_clk new_AGEMA_reg_buffer_943 ( .C (clk), .D (SubCellInst_SboxInst_7_n7), .Q (new_AGEMA_signal_2303) ) ;
    buf_clk new_AGEMA_reg_buffer_945 ( .C (clk), .D (new_AGEMA_signal_1080), .Q (new_AGEMA_signal_2305) ) ;
    buf_clk new_AGEMA_reg_buffer_947 ( .C (clk), .D (ciphertext_s0[17]), .Q (new_AGEMA_signal_2307) ) ;
    buf_clk new_AGEMA_reg_buffer_949 ( .C (clk), .D (ciphertext_s1[17]), .Q (new_AGEMA_signal_2309) ) ;
    buf_clk new_AGEMA_reg_buffer_951 ( .C (clk), .D (SubCellInst_SboxInst_8_n9), .Q (new_AGEMA_signal_2311) ) ;
    buf_clk new_AGEMA_reg_buffer_953 ( .C (clk), .D (new_AGEMA_signal_1090), .Q (new_AGEMA_signal_2313) ) ;
    buf_clk new_AGEMA_reg_buffer_955 ( .C (clk), .D (ciphertext_s0[16]), .Q (new_AGEMA_signal_2315) ) ;
    buf_clk new_AGEMA_reg_buffer_957 ( .C (clk), .D (ciphertext_s1[16]), .Q (new_AGEMA_signal_2317) ) ;
    buf_clk new_AGEMA_reg_buffer_959 ( .C (clk), .D (SubCellInst_SboxInst_8_n7), .Q (new_AGEMA_signal_2319) ) ;
    buf_clk new_AGEMA_reg_buffer_961 ( .C (clk), .D (new_AGEMA_signal_1088), .Q (new_AGEMA_signal_2321) ) ;
    buf_clk new_AGEMA_reg_buffer_963 ( .C (clk), .D (ciphertext_s0[29]), .Q (new_AGEMA_signal_2323) ) ;
    buf_clk new_AGEMA_reg_buffer_965 ( .C (clk), .D (ciphertext_s1[29]), .Q (new_AGEMA_signal_2325) ) ;
    buf_clk new_AGEMA_reg_buffer_967 ( .C (clk), .D (SubCellInst_SboxInst_9_n9), .Q (new_AGEMA_signal_2327) ) ;
    buf_clk new_AGEMA_reg_buffer_969 ( .C (clk), .D (new_AGEMA_signal_1098), .Q (new_AGEMA_signal_2329) ) ;
    buf_clk new_AGEMA_reg_buffer_971 ( .C (clk), .D (ciphertext_s0[28]), .Q (new_AGEMA_signal_2331) ) ;
    buf_clk new_AGEMA_reg_buffer_973 ( .C (clk), .D (ciphertext_s1[28]), .Q (new_AGEMA_signal_2333) ) ;
    buf_clk new_AGEMA_reg_buffer_975 ( .C (clk), .D (SubCellInst_SboxInst_9_n7), .Q (new_AGEMA_signal_2335) ) ;
    buf_clk new_AGEMA_reg_buffer_977 ( .C (clk), .D (new_AGEMA_signal_1096), .Q (new_AGEMA_signal_2337) ) ;
    buf_clk new_AGEMA_reg_buffer_979 ( .C (clk), .D (ciphertext_s0[25]), .Q (new_AGEMA_signal_2339) ) ;
    buf_clk new_AGEMA_reg_buffer_981 ( .C (clk), .D (ciphertext_s1[25]), .Q (new_AGEMA_signal_2341) ) ;
    buf_clk new_AGEMA_reg_buffer_983 ( .C (clk), .D (SubCellInst_SboxInst_10_n9), .Q (new_AGEMA_signal_2343) ) ;
    buf_clk new_AGEMA_reg_buffer_985 ( .C (clk), .D (new_AGEMA_signal_1106), .Q (new_AGEMA_signal_2345) ) ;
    buf_clk new_AGEMA_reg_buffer_987 ( .C (clk), .D (ciphertext_s0[24]), .Q (new_AGEMA_signal_2347) ) ;
    buf_clk new_AGEMA_reg_buffer_989 ( .C (clk), .D (ciphertext_s1[24]), .Q (new_AGEMA_signal_2349) ) ;
    buf_clk new_AGEMA_reg_buffer_991 ( .C (clk), .D (SubCellInst_SboxInst_10_n7), .Q (new_AGEMA_signal_2351) ) ;
    buf_clk new_AGEMA_reg_buffer_993 ( .C (clk), .D (new_AGEMA_signal_1104), .Q (new_AGEMA_signal_2353) ) ;
    buf_clk new_AGEMA_reg_buffer_995 ( .C (clk), .D (ciphertext_s0[21]), .Q (new_AGEMA_signal_2355) ) ;
    buf_clk new_AGEMA_reg_buffer_997 ( .C (clk), .D (ciphertext_s1[21]), .Q (new_AGEMA_signal_2357) ) ;
    buf_clk new_AGEMA_reg_buffer_999 ( .C (clk), .D (SubCellInst_SboxInst_11_n9), .Q (new_AGEMA_signal_2359) ) ;
    buf_clk new_AGEMA_reg_buffer_1001 ( .C (clk), .D (new_AGEMA_signal_1114), .Q (new_AGEMA_signal_2361) ) ;
    buf_clk new_AGEMA_reg_buffer_1003 ( .C (clk), .D (ciphertext_s0[20]), .Q (new_AGEMA_signal_2363) ) ;
    buf_clk new_AGEMA_reg_buffer_1005 ( .C (clk), .D (ciphertext_s1[20]), .Q (new_AGEMA_signal_2365) ) ;
    buf_clk new_AGEMA_reg_buffer_1007 ( .C (clk), .D (SubCellInst_SboxInst_11_n7), .Q (new_AGEMA_signal_2367) ) ;
    buf_clk new_AGEMA_reg_buffer_1009 ( .C (clk), .D (new_AGEMA_signal_1112), .Q (new_AGEMA_signal_2369) ) ;
    buf_clk new_AGEMA_reg_buffer_1011 ( .C (clk), .D (ciphertext_s0[5]), .Q (new_AGEMA_signal_2371) ) ;
    buf_clk new_AGEMA_reg_buffer_1013 ( .C (clk), .D (ciphertext_s1[5]), .Q (new_AGEMA_signal_2373) ) ;
    buf_clk new_AGEMA_reg_buffer_1015 ( .C (clk), .D (SubCellInst_SboxInst_12_n9), .Q (new_AGEMA_signal_2375) ) ;
    buf_clk new_AGEMA_reg_buffer_1017 ( .C (clk), .D (new_AGEMA_signal_1122), .Q (new_AGEMA_signal_2377) ) ;
    buf_clk new_AGEMA_reg_buffer_1019 ( .C (clk), .D (ciphertext_s0[4]), .Q (new_AGEMA_signal_2379) ) ;
    buf_clk new_AGEMA_reg_buffer_1021 ( .C (clk), .D (ciphertext_s1[4]), .Q (new_AGEMA_signal_2381) ) ;
    buf_clk new_AGEMA_reg_buffer_1023 ( .C (clk), .D (SubCellInst_SboxInst_12_n7), .Q (new_AGEMA_signal_2383) ) ;
    buf_clk new_AGEMA_reg_buffer_1025 ( .C (clk), .D (new_AGEMA_signal_1120), .Q (new_AGEMA_signal_2385) ) ;
    buf_clk new_AGEMA_reg_buffer_1027 ( .C (clk), .D (ciphertext_s0[9]), .Q (new_AGEMA_signal_2387) ) ;
    buf_clk new_AGEMA_reg_buffer_1029 ( .C (clk), .D (ciphertext_s1[9]), .Q (new_AGEMA_signal_2389) ) ;
    buf_clk new_AGEMA_reg_buffer_1031 ( .C (clk), .D (SubCellInst_SboxInst_13_n9), .Q (new_AGEMA_signal_2391) ) ;
    buf_clk new_AGEMA_reg_buffer_1033 ( .C (clk), .D (new_AGEMA_signal_1130), .Q (new_AGEMA_signal_2393) ) ;
    buf_clk new_AGEMA_reg_buffer_1035 ( .C (clk), .D (ciphertext_s0[8]), .Q (new_AGEMA_signal_2395) ) ;
    buf_clk new_AGEMA_reg_buffer_1037 ( .C (clk), .D (ciphertext_s1[8]), .Q (new_AGEMA_signal_2397) ) ;
    buf_clk new_AGEMA_reg_buffer_1039 ( .C (clk), .D (SubCellInst_SboxInst_13_n7), .Q (new_AGEMA_signal_2399) ) ;
    buf_clk new_AGEMA_reg_buffer_1041 ( .C (clk), .D (new_AGEMA_signal_1128), .Q (new_AGEMA_signal_2401) ) ;
    buf_clk new_AGEMA_reg_buffer_1043 ( .C (clk), .D (ciphertext_s0[13]), .Q (new_AGEMA_signal_2403) ) ;
    buf_clk new_AGEMA_reg_buffer_1045 ( .C (clk), .D (ciphertext_s1[13]), .Q (new_AGEMA_signal_2405) ) ;
    buf_clk new_AGEMA_reg_buffer_1047 ( .C (clk), .D (SubCellInst_SboxInst_14_n9), .Q (new_AGEMA_signal_2407) ) ;
    buf_clk new_AGEMA_reg_buffer_1049 ( .C (clk), .D (new_AGEMA_signal_1138), .Q (new_AGEMA_signal_2409) ) ;
    buf_clk new_AGEMA_reg_buffer_1051 ( .C (clk), .D (ciphertext_s0[12]), .Q (new_AGEMA_signal_2411) ) ;
    buf_clk new_AGEMA_reg_buffer_1053 ( .C (clk), .D (ciphertext_s1[12]), .Q (new_AGEMA_signal_2413) ) ;
    buf_clk new_AGEMA_reg_buffer_1055 ( .C (clk), .D (SubCellInst_SboxInst_14_n7), .Q (new_AGEMA_signal_2415) ) ;
    buf_clk new_AGEMA_reg_buffer_1057 ( .C (clk), .D (new_AGEMA_signal_1136), .Q (new_AGEMA_signal_2417) ) ;
    buf_clk new_AGEMA_reg_buffer_1059 ( .C (clk), .D (ciphertext_s0[1]), .Q (new_AGEMA_signal_2419) ) ;
    buf_clk new_AGEMA_reg_buffer_1061 ( .C (clk), .D (ciphertext_s1[1]), .Q (new_AGEMA_signal_2421) ) ;
    buf_clk new_AGEMA_reg_buffer_1063 ( .C (clk), .D (SubCellInst_SboxInst_15_n9), .Q (new_AGEMA_signal_2423) ) ;
    buf_clk new_AGEMA_reg_buffer_1065 ( .C (clk), .D (new_AGEMA_signal_1146), .Q (new_AGEMA_signal_2425) ) ;
    buf_clk new_AGEMA_reg_buffer_1067 ( .C (clk), .D (ciphertext_s0[0]), .Q (new_AGEMA_signal_2427) ) ;
    buf_clk new_AGEMA_reg_buffer_1069 ( .C (clk), .D (ciphertext_s1[0]), .Q (new_AGEMA_signal_2429) ) ;
    buf_clk new_AGEMA_reg_buffer_1071 ( .C (clk), .D (SubCellInst_SboxInst_15_n7), .Q (new_AGEMA_signal_2431) ) ;
    buf_clk new_AGEMA_reg_buffer_1073 ( .C (clk), .D (new_AGEMA_signal_1144), .Q (new_AGEMA_signal_2433) ) ;
    buf_clk new_AGEMA_reg_buffer_1075 ( .C (clk), .D (rst), .Q (new_AGEMA_signal_2435) ) ;
    buf_clk new_AGEMA_reg_buffer_1081 ( .C (clk), .D (plaintext_s0[1]), .Q (new_AGEMA_signal_2441) ) ;
    buf_clk new_AGEMA_reg_buffer_1087 ( .C (clk), .D (plaintext_s1[1]), .Q (new_AGEMA_signal_2447) ) ;
    buf_clk new_AGEMA_reg_buffer_1093 ( .C (clk), .D (plaintext_s0[3]), .Q (new_AGEMA_signal_2453) ) ;
    buf_clk new_AGEMA_reg_buffer_1099 ( .C (clk), .D (plaintext_s1[3]), .Q (new_AGEMA_signal_2459) ) ;
    buf_clk new_AGEMA_reg_buffer_1105 ( .C (clk), .D (plaintext_s0[5]), .Q (new_AGEMA_signal_2465) ) ;
    buf_clk new_AGEMA_reg_buffer_1111 ( .C (clk), .D (plaintext_s1[5]), .Q (new_AGEMA_signal_2471) ) ;
    buf_clk new_AGEMA_reg_buffer_1117 ( .C (clk), .D (plaintext_s0[7]), .Q (new_AGEMA_signal_2477) ) ;
    buf_clk new_AGEMA_reg_buffer_1123 ( .C (clk), .D (plaintext_s1[7]), .Q (new_AGEMA_signal_2483) ) ;
    buf_clk new_AGEMA_reg_buffer_1129 ( .C (clk), .D (plaintext_s0[9]), .Q (new_AGEMA_signal_2489) ) ;
    buf_clk new_AGEMA_reg_buffer_1135 ( .C (clk), .D (plaintext_s1[9]), .Q (new_AGEMA_signal_2495) ) ;
    buf_clk new_AGEMA_reg_buffer_1141 ( .C (clk), .D (plaintext_s0[11]), .Q (new_AGEMA_signal_2501) ) ;
    buf_clk new_AGEMA_reg_buffer_1147 ( .C (clk), .D (plaintext_s1[11]), .Q (new_AGEMA_signal_2507) ) ;
    buf_clk new_AGEMA_reg_buffer_1153 ( .C (clk), .D (plaintext_s0[13]), .Q (new_AGEMA_signal_2513) ) ;
    buf_clk new_AGEMA_reg_buffer_1159 ( .C (clk), .D (plaintext_s1[13]), .Q (new_AGEMA_signal_2519) ) ;
    buf_clk new_AGEMA_reg_buffer_1165 ( .C (clk), .D (plaintext_s0[15]), .Q (new_AGEMA_signal_2525) ) ;
    buf_clk new_AGEMA_reg_buffer_1171 ( .C (clk), .D (plaintext_s1[15]), .Q (new_AGEMA_signal_2531) ) ;
    buf_clk new_AGEMA_reg_buffer_1177 ( .C (clk), .D (plaintext_s0[17]), .Q (new_AGEMA_signal_2537) ) ;
    buf_clk new_AGEMA_reg_buffer_1183 ( .C (clk), .D (plaintext_s1[17]), .Q (new_AGEMA_signal_2543) ) ;
    buf_clk new_AGEMA_reg_buffer_1189 ( .C (clk), .D (plaintext_s0[19]), .Q (new_AGEMA_signal_2549) ) ;
    buf_clk new_AGEMA_reg_buffer_1195 ( .C (clk), .D (plaintext_s1[19]), .Q (new_AGEMA_signal_2555) ) ;
    buf_clk new_AGEMA_reg_buffer_1201 ( .C (clk), .D (plaintext_s0[21]), .Q (new_AGEMA_signal_2561) ) ;
    buf_clk new_AGEMA_reg_buffer_1207 ( .C (clk), .D (plaintext_s1[21]), .Q (new_AGEMA_signal_2567) ) ;
    buf_clk new_AGEMA_reg_buffer_1213 ( .C (clk), .D (plaintext_s0[23]), .Q (new_AGEMA_signal_2573) ) ;
    buf_clk new_AGEMA_reg_buffer_1219 ( .C (clk), .D (plaintext_s1[23]), .Q (new_AGEMA_signal_2579) ) ;
    buf_clk new_AGEMA_reg_buffer_1225 ( .C (clk), .D (plaintext_s0[25]), .Q (new_AGEMA_signal_2585) ) ;
    buf_clk new_AGEMA_reg_buffer_1231 ( .C (clk), .D (plaintext_s1[25]), .Q (new_AGEMA_signal_2591) ) ;
    buf_clk new_AGEMA_reg_buffer_1237 ( .C (clk), .D (plaintext_s0[27]), .Q (new_AGEMA_signal_2597) ) ;
    buf_clk new_AGEMA_reg_buffer_1243 ( .C (clk), .D (plaintext_s1[27]), .Q (new_AGEMA_signal_2603) ) ;
    buf_clk new_AGEMA_reg_buffer_1249 ( .C (clk), .D (plaintext_s0[29]), .Q (new_AGEMA_signal_2609) ) ;
    buf_clk new_AGEMA_reg_buffer_1255 ( .C (clk), .D (plaintext_s1[29]), .Q (new_AGEMA_signal_2615) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C (clk), .D (plaintext_s0[31]), .Q (new_AGEMA_signal_2621) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C (clk), .D (plaintext_s1[31]), .Q (new_AGEMA_signal_2627) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C (clk), .D (plaintext_s0[33]), .Q (new_AGEMA_signal_2633) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C (clk), .D (plaintext_s1[33]), .Q (new_AGEMA_signal_2639) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C (clk), .D (plaintext_s0[35]), .Q (new_AGEMA_signal_2645) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C (clk), .D (plaintext_s1[35]), .Q (new_AGEMA_signal_2651) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C (clk), .D (plaintext_s0[37]), .Q (new_AGEMA_signal_2657) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C (clk), .D (plaintext_s1[37]), .Q (new_AGEMA_signal_2663) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C (clk), .D (plaintext_s0[39]), .Q (new_AGEMA_signal_2669) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C (clk), .D (plaintext_s1[39]), .Q (new_AGEMA_signal_2675) ) ;
    buf_clk new_AGEMA_reg_buffer_1321 ( .C (clk), .D (plaintext_s0[41]), .Q (new_AGEMA_signal_2681) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C (clk), .D (plaintext_s1[41]), .Q (new_AGEMA_signal_2687) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C (clk), .D (plaintext_s0[43]), .Q (new_AGEMA_signal_2693) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C (clk), .D (plaintext_s1[43]), .Q (new_AGEMA_signal_2699) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C (clk), .D (plaintext_s0[45]), .Q (new_AGEMA_signal_2705) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C (clk), .D (plaintext_s1[45]), .Q (new_AGEMA_signal_2711) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C (clk), .D (plaintext_s0[47]), .Q (new_AGEMA_signal_2717) ) ;
    buf_clk new_AGEMA_reg_buffer_1363 ( .C (clk), .D (plaintext_s1[47]), .Q (new_AGEMA_signal_2723) ) ;
    buf_clk new_AGEMA_reg_buffer_1369 ( .C (clk), .D (plaintext_s0[49]), .Q (new_AGEMA_signal_2729) ) ;
    buf_clk new_AGEMA_reg_buffer_1375 ( .C (clk), .D (plaintext_s1[49]), .Q (new_AGEMA_signal_2735) ) ;
    buf_clk new_AGEMA_reg_buffer_1381 ( .C (clk), .D (plaintext_s0[51]), .Q (new_AGEMA_signal_2741) ) ;
    buf_clk new_AGEMA_reg_buffer_1387 ( .C (clk), .D (plaintext_s1[51]), .Q (new_AGEMA_signal_2747) ) ;
    buf_clk new_AGEMA_reg_buffer_1393 ( .C (clk), .D (plaintext_s0[53]), .Q (new_AGEMA_signal_2753) ) ;
    buf_clk new_AGEMA_reg_buffer_1399 ( .C (clk), .D (plaintext_s1[53]), .Q (new_AGEMA_signal_2759) ) ;
    buf_clk new_AGEMA_reg_buffer_1405 ( .C (clk), .D (plaintext_s0[55]), .Q (new_AGEMA_signal_2765) ) ;
    buf_clk new_AGEMA_reg_buffer_1411 ( .C (clk), .D (plaintext_s1[55]), .Q (new_AGEMA_signal_2771) ) ;
    buf_clk new_AGEMA_reg_buffer_1417 ( .C (clk), .D (plaintext_s0[57]), .Q (new_AGEMA_signal_2777) ) ;
    buf_clk new_AGEMA_reg_buffer_1423 ( .C (clk), .D (plaintext_s1[57]), .Q (new_AGEMA_signal_2783) ) ;
    buf_clk new_AGEMA_reg_buffer_1429 ( .C (clk), .D (plaintext_s0[59]), .Q (new_AGEMA_signal_2789) ) ;
    buf_clk new_AGEMA_reg_buffer_1435 ( .C (clk), .D (plaintext_s1[59]), .Q (new_AGEMA_signal_2795) ) ;
    buf_clk new_AGEMA_reg_buffer_1441 ( .C (clk), .D (plaintext_s0[61]), .Q (new_AGEMA_signal_2801) ) ;
    buf_clk new_AGEMA_reg_buffer_1447 ( .C (clk), .D (plaintext_s1[61]), .Q (new_AGEMA_signal_2807) ) ;
    buf_clk new_AGEMA_reg_buffer_1453 ( .C (clk), .D (plaintext_s0[63]), .Q (new_AGEMA_signal_2813) ) ;
    buf_clk new_AGEMA_reg_buffer_1459 ( .C (clk), .D (plaintext_s1[63]), .Q (new_AGEMA_signal_2819) ) ;
    buf_clk new_AGEMA_reg_buffer_1465 ( .C (clk), .D (SelectedKey[49]), .Q (new_AGEMA_signal_2825) ) ;
    buf_clk new_AGEMA_reg_buffer_1471 ( .C (clk), .D (new_AGEMA_signal_1551), .Q (new_AGEMA_signal_2831) ) ;
    buf_clk new_AGEMA_reg_buffer_1477 ( .C (clk), .D (SelectedKey[51]), .Q (new_AGEMA_signal_2837) ) ;
    buf_clk new_AGEMA_reg_buffer_1483 ( .C (clk), .D (new_AGEMA_signal_1557), .Q (new_AGEMA_signal_2843) ) ;
    buf_clk new_AGEMA_reg_buffer_1489 ( .C (clk), .D (SelectedKey[53]), .Q (new_AGEMA_signal_2849) ) ;
    buf_clk new_AGEMA_reg_buffer_1495 ( .C (clk), .D (new_AGEMA_signal_1278), .Q (new_AGEMA_signal_2855) ) ;
    buf_clk new_AGEMA_reg_buffer_1501 ( .C (clk), .D (SelectedKey[55]), .Q (new_AGEMA_signal_2861) ) ;
    buf_clk new_AGEMA_reg_buffer_1507 ( .C (clk), .D (new_AGEMA_signal_1563), .Q (new_AGEMA_signal_2867) ) ;
    buf_clk new_AGEMA_reg_buffer_1513 ( .C (clk), .D (SelectedKey[57]), .Q (new_AGEMA_signal_2873) ) ;
    buf_clk new_AGEMA_reg_buffer_1519 ( .C (clk), .D (new_AGEMA_signal_1566), .Q (new_AGEMA_signal_2879) ) ;
    buf_clk new_AGEMA_reg_buffer_1525 ( .C (clk), .D (SelectedKey[59]), .Q (new_AGEMA_signal_2885) ) ;
    buf_clk new_AGEMA_reg_buffer_1531 ( .C (clk), .D (new_AGEMA_signal_1287), .Q (new_AGEMA_signal_2891) ) ;
    buf_clk new_AGEMA_reg_buffer_1537 ( .C (clk), .D (SelectedKey[61]), .Q (new_AGEMA_signal_2897) ) ;
    buf_clk new_AGEMA_reg_buffer_1543 ( .C (clk), .D (new_AGEMA_signal_1575), .Q (new_AGEMA_signal_2903) ) ;
    buf_clk new_AGEMA_reg_buffer_1549 ( .C (clk), .D (SelectedKey[63]), .Q (new_AGEMA_signal_2909) ) ;
    buf_clk new_AGEMA_reg_buffer_1555 ( .C (clk), .D (new_AGEMA_signal_1578), .Q (new_AGEMA_signal_2915) ) ;
    buf_clk new_AGEMA_reg_buffer_1561 ( .C (clk), .D (AddKeyConstXOR_XORInst_0_1_n1), .Q (new_AGEMA_signal_2921) ) ;
    buf_clk new_AGEMA_reg_buffer_1567 ( .C (clk), .D (new_AGEMA_signal_1708), .Q (new_AGEMA_signal_2927) ) ;
    buf_clk new_AGEMA_reg_buffer_1573 ( .C (clk), .D (AddKeyConstXOR_XORInst_0_3_n1), .Q (new_AGEMA_signal_2933) ) ;
    buf_clk new_AGEMA_reg_buffer_1579 ( .C (clk), .D (new_AGEMA_signal_1710), .Q (new_AGEMA_signal_2939) ) ;
    buf_clk new_AGEMA_reg_buffer_1585 ( .C (clk), .D (AddKeyConstXOR_XORInst_1_1_n1), .Q (new_AGEMA_signal_2945) ) ;
    buf_clk new_AGEMA_reg_buffer_1591 ( .C (clk), .D (new_AGEMA_signal_1712), .Q (new_AGEMA_signal_2951) ) ;
    buf_clk new_AGEMA_reg_buffer_1597 ( .C (clk), .D (AddKeyConstXOR_XORInst_1_3_n1), .Q (new_AGEMA_signal_2957) ) ;
    buf_clk new_AGEMA_reg_buffer_1603 ( .C (clk), .D (new_AGEMA_signal_1714), .Q (new_AGEMA_signal_2963) ) ;
    buf_clk new_AGEMA_reg_buffer_1609 ( .C (clk), .D (SelectedKey[1]), .Q (new_AGEMA_signal_2969) ) ;
    buf_clk new_AGEMA_reg_buffer_1615 ( .C (clk), .D (new_AGEMA_signal_1437), .Q (new_AGEMA_signal_2975) ) ;
    buf_clk new_AGEMA_reg_buffer_1621 ( .C (clk), .D (SelectedKey[3]), .Q (new_AGEMA_signal_2981) ) ;
    buf_clk new_AGEMA_reg_buffer_1627 ( .C (clk), .D (new_AGEMA_signal_1440), .Q (new_AGEMA_signal_2987) ) ;
    buf_clk new_AGEMA_reg_buffer_1633 ( .C (clk), .D (SelectedKey[5]), .Q (new_AGEMA_signal_2993) ) ;
    buf_clk new_AGEMA_reg_buffer_1639 ( .C (clk), .D (new_AGEMA_signal_1446), .Q (new_AGEMA_signal_2999) ) ;
    buf_clk new_AGEMA_reg_buffer_1645 ( .C (clk), .D (SelectedKey[7]), .Q (new_AGEMA_signal_3005) ) ;
    buf_clk new_AGEMA_reg_buffer_1651 ( .C (clk), .D (new_AGEMA_signal_1452), .Q (new_AGEMA_signal_3011) ) ;
    buf_clk new_AGEMA_reg_buffer_1657 ( .C (clk), .D (SelectedKey[9]), .Q (new_AGEMA_signal_3017) ) ;
    buf_clk new_AGEMA_reg_buffer_1663 ( .C (clk), .D (new_AGEMA_signal_1458), .Q (new_AGEMA_signal_3023) ) ;
    buf_clk new_AGEMA_reg_buffer_1669 ( .C (clk), .D (SelectedKey[11]), .Q (new_AGEMA_signal_3029) ) ;
    buf_clk new_AGEMA_reg_buffer_1675 ( .C (clk), .D (new_AGEMA_signal_1464), .Q (new_AGEMA_signal_3035) ) ;
    buf_clk new_AGEMA_reg_buffer_1681 ( .C (clk), .D (SelectedKey[13]), .Q (new_AGEMA_signal_3041) ) ;
    buf_clk new_AGEMA_reg_buffer_1687 ( .C (clk), .D (new_AGEMA_signal_1470), .Q (new_AGEMA_signal_3047) ) ;
    buf_clk new_AGEMA_reg_buffer_1693 ( .C (clk), .D (SelectedKey[15]), .Q (new_AGEMA_signal_3053) ) ;
    buf_clk new_AGEMA_reg_buffer_1699 ( .C (clk), .D (new_AGEMA_signal_1476), .Q (new_AGEMA_signal_3059) ) ;
    buf_clk new_AGEMA_reg_buffer_1705 ( .C (clk), .D (SelectedKey[17]), .Q (new_AGEMA_signal_3065) ) ;
    buf_clk new_AGEMA_reg_buffer_1711 ( .C (clk), .D (new_AGEMA_signal_1482), .Q (new_AGEMA_signal_3071) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C (clk), .D (SelectedKey[19]), .Q (new_AGEMA_signal_3077) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C (clk), .D (new_AGEMA_signal_1488), .Q (new_AGEMA_signal_3083) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C (clk), .D (SelectedKey[21]), .Q (new_AGEMA_signal_3089) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C (clk), .D (new_AGEMA_signal_1494), .Q (new_AGEMA_signal_3095) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C (clk), .D (SelectedKey[23]), .Q (new_AGEMA_signal_3101) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C (clk), .D (new_AGEMA_signal_1254), .Q (new_AGEMA_signal_3107) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C (clk), .D (SelectedKey[25]), .Q (new_AGEMA_signal_3113) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C (clk), .D (new_AGEMA_signal_1260), .Q (new_AGEMA_signal_3119) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C (clk), .D (SelectedKey[27]), .Q (new_AGEMA_signal_3125) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C (clk), .D (new_AGEMA_signal_1266), .Q (new_AGEMA_signal_3131) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C (clk), .D (SelectedKey[29]), .Q (new_AGEMA_signal_3137) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C (clk), .D (new_AGEMA_signal_1500), .Q (new_AGEMA_signal_3143) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C (clk), .D (SelectedKey[31]), .Q (new_AGEMA_signal_3149) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C (clk), .D (new_AGEMA_signal_1506), .Q (new_AGEMA_signal_3155) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C (clk), .D (SelectedKey[33]), .Q (new_AGEMA_signal_3161) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C (clk), .D (new_AGEMA_signal_1269), .Q (new_AGEMA_signal_3167) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C (clk), .D (SelectedKey[35]), .Q (new_AGEMA_signal_3173) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C (clk), .D (new_AGEMA_signal_1515), .Q (new_AGEMA_signal_3179) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C (clk), .D (SelectedKey[37]), .Q (new_AGEMA_signal_3185) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C (clk), .D (new_AGEMA_signal_1518), .Q (new_AGEMA_signal_3191) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C (clk), .D (SelectedKey[39]), .Q (new_AGEMA_signal_3197) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C (clk), .D (new_AGEMA_signal_1275), .Q (new_AGEMA_signal_3203) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C (clk), .D (plaintext_s0[0]), .Q (new_AGEMA_signal_3403) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C (clk), .D (plaintext_s1[0]), .Q (new_AGEMA_signal_3411) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C (clk), .D (plaintext_s0[2]), .Q (new_AGEMA_signal_3419) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C (clk), .D (plaintext_s1[2]), .Q (new_AGEMA_signal_3427) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C (clk), .D (plaintext_s0[4]), .Q (new_AGEMA_signal_3435) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C (clk), .D (plaintext_s1[4]), .Q (new_AGEMA_signal_3443) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C (clk), .D (plaintext_s0[6]), .Q (new_AGEMA_signal_3451) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C (clk), .D (plaintext_s1[6]), .Q (new_AGEMA_signal_3459) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C (clk), .D (plaintext_s0[8]), .Q (new_AGEMA_signal_3467) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C (clk), .D (plaintext_s1[8]), .Q (new_AGEMA_signal_3475) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C (clk), .D (plaintext_s0[10]), .Q (new_AGEMA_signal_3483) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C (clk), .D (plaintext_s1[10]), .Q (new_AGEMA_signal_3491) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C (clk), .D (plaintext_s0[12]), .Q (new_AGEMA_signal_3499) ) ;
    buf_clk new_AGEMA_reg_buffer_2147 ( .C (clk), .D (plaintext_s1[12]), .Q (new_AGEMA_signal_3507) ) ;
    buf_clk new_AGEMA_reg_buffer_2155 ( .C (clk), .D (plaintext_s0[14]), .Q (new_AGEMA_signal_3515) ) ;
    buf_clk new_AGEMA_reg_buffer_2163 ( .C (clk), .D (plaintext_s1[14]), .Q (new_AGEMA_signal_3523) ) ;
    buf_clk new_AGEMA_reg_buffer_2171 ( .C (clk), .D (plaintext_s0[16]), .Q (new_AGEMA_signal_3531) ) ;
    buf_clk new_AGEMA_reg_buffer_2179 ( .C (clk), .D (plaintext_s1[16]), .Q (new_AGEMA_signal_3539) ) ;
    buf_clk new_AGEMA_reg_buffer_2187 ( .C (clk), .D (plaintext_s0[18]), .Q (new_AGEMA_signal_3547) ) ;
    buf_clk new_AGEMA_reg_buffer_2195 ( .C (clk), .D (plaintext_s1[18]), .Q (new_AGEMA_signal_3555) ) ;
    buf_clk new_AGEMA_reg_buffer_2203 ( .C (clk), .D (plaintext_s0[20]), .Q (new_AGEMA_signal_3563) ) ;
    buf_clk new_AGEMA_reg_buffer_2211 ( .C (clk), .D (plaintext_s1[20]), .Q (new_AGEMA_signal_3571) ) ;
    buf_clk new_AGEMA_reg_buffer_2219 ( .C (clk), .D (plaintext_s0[22]), .Q (new_AGEMA_signal_3579) ) ;
    buf_clk new_AGEMA_reg_buffer_2227 ( .C (clk), .D (plaintext_s1[22]), .Q (new_AGEMA_signal_3587) ) ;
    buf_clk new_AGEMA_reg_buffer_2235 ( .C (clk), .D (plaintext_s0[24]), .Q (new_AGEMA_signal_3595) ) ;
    buf_clk new_AGEMA_reg_buffer_2243 ( .C (clk), .D (plaintext_s1[24]), .Q (new_AGEMA_signal_3603) ) ;
    buf_clk new_AGEMA_reg_buffer_2251 ( .C (clk), .D (plaintext_s0[26]), .Q (new_AGEMA_signal_3611) ) ;
    buf_clk new_AGEMA_reg_buffer_2259 ( .C (clk), .D (plaintext_s1[26]), .Q (new_AGEMA_signal_3619) ) ;
    buf_clk new_AGEMA_reg_buffer_2267 ( .C (clk), .D (plaintext_s0[28]), .Q (new_AGEMA_signal_3627) ) ;
    buf_clk new_AGEMA_reg_buffer_2275 ( .C (clk), .D (plaintext_s1[28]), .Q (new_AGEMA_signal_3635) ) ;
    buf_clk new_AGEMA_reg_buffer_2283 ( .C (clk), .D (plaintext_s0[30]), .Q (new_AGEMA_signal_3643) ) ;
    buf_clk new_AGEMA_reg_buffer_2291 ( .C (clk), .D (plaintext_s1[30]), .Q (new_AGEMA_signal_3651) ) ;
    buf_clk new_AGEMA_reg_buffer_2299 ( .C (clk), .D (plaintext_s0[32]), .Q (new_AGEMA_signal_3659) ) ;
    buf_clk new_AGEMA_reg_buffer_2307 ( .C (clk), .D (plaintext_s1[32]), .Q (new_AGEMA_signal_3667) ) ;
    buf_clk new_AGEMA_reg_buffer_2315 ( .C (clk), .D (plaintext_s0[34]), .Q (new_AGEMA_signal_3675) ) ;
    buf_clk new_AGEMA_reg_buffer_2323 ( .C (clk), .D (plaintext_s1[34]), .Q (new_AGEMA_signal_3683) ) ;
    buf_clk new_AGEMA_reg_buffer_2331 ( .C (clk), .D (plaintext_s0[36]), .Q (new_AGEMA_signal_3691) ) ;
    buf_clk new_AGEMA_reg_buffer_2339 ( .C (clk), .D (plaintext_s1[36]), .Q (new_AGEMA_signal_3699) ) ;
    buf_clk new_AGEMA_reg_buffer_2347 ( .C (clk), .D (plaintext_s0[38]), .Q (new_AGEMA_signal_3707) ) ;
    buf_clk new_AGEMA_reg_buffer_2355 ( .C (clk), .D (plaintext_s1[38]), .Q (new_AGEMA_signal_3715) ) ;
    buf_clk new_AGEMA_reg_buffer_2363 ( .C (clk), .D (plaintext_s0[40]), .Q (new_AGEMA_signal_3723) ) ;
    buf_clk new_AGEMA_reg_buffer_2371 ( .C (clk), .D (plaintext_s1[40]), .Q (new_AGEMA_signal_3731) ) ;
    buf_clk new_AGEMA_reg_buffer_2379 ( .C (clk), .D (plaintext_s0[42]), .Q (new_AGEMA_signal_3739) ) ;
    buf_clk new_AGEMA_reg_buffer_2387 ( .C (clk), .D (plaintext_s1[42]), .Q (new_AGEMA_signal_3747) ) ;
    buf_clk new_AGEMA_reg_buffer_2395 ( .C (clk), .D (plaintext_s0[44]), .Q (new_AGEMA_signal_3755) ) ;
    buf_clk new_AGEMA_reg_buffer_2403 ( .C (clk), .D (plaintext_s1[44]), .Q (new_AGEMA_signal_3763) ) ;
    buf_clk new_AGEMA_reg_buffer_2411 ( .C (clk), .D (plaintext_s0[46]), .Q (new_AGEMA_signal_3771) ) ;
    buf_clk new_AGEMA_reg_buffer_2419 ( .C (clk), .D (plaintext_s1[46]), .Q (new_AGEMA_signal_3779) ) ;
    buf_clk new_AGEMA_reg_buffer_2427 ( .C (clk), .D (plaintext_s0[48]), .Q (new_AGEMA_signal_3787) ) ;
    buf_clk new_AGEMA_reg_buffer_2435 ( .C (clk), .D (plaintext_s1[48]), .Q (new_AGEMA_signal_3795) ) ;
    buf_clk new_AGEMA_reg_buffer_2443 ( .C (clk), .D (plaintext_s0[50]), .Q (new_AGEMA_signal_3803) ) ;
    buf_clk new_AGEMA_reg_buffer_2451 ( .C (clk), .D (plaintext_s1[50]), .Q (new_AGEMA_signal_3811) ) ;
    buf_clk new_AGEMA_reg_buffer_2459 ( .C (clk), .D (plaintext_s0[52]), .Q (new_AGEMA_signal_3819) ) ;
    buf_clk new_AGEMA_reg_buffer_2467 ( .C (clk), .D (plaintext_s1[52]), .Q (new_AGEMA_signal_3827) ) ;
    buf_clk new_AGEMA_reg_buffer_2475 ( .C (clk), .D (plaintext_s0[54]), .Q (new_AGEMA_signal_3835) ) ;
    buf_clk new_AGEMA_reg_buffer_2483 ( .C (clk), .D (plaintext_s1[54]), .Q (new_AGEMA_signal_3843) ) ;
    buf_clk new_AGEMA_reg_buffer_2491 ( .C (clk), .D (plaintext_s0[56]), .Q (new_AGEMA_signal_3851) ) ;
    buf_clk new_AGEMA_reg_buffer_2499 ( .C (clk), .D (plaintext_s1[56]), .Q (new_AGEMA_signal_3859) ) ;
    buf_clk new_AGEMA_reg_buffer_2507 ( .C (clk), .D (plaintext_s0[58]), .Q (new_AGEMA_signal_3867) ) ;
    buf_clk new_AGEMA_reg_buffer_2515 ( .C (clk), .D (plaintext_s1[58]), .Q (new_AGEMA_signal_3875) ) ;
    buf_clk new_AGEMA_reg_buffer_2523 ( .C (clk), .D (plaintext_s0[60]), .Q (new_AGEMA_signal_3883) ) ;
    buf_clk new_AGEMA_reg_buffer_2531 ( .C (clk), .D (plaintext_s1[60]), .Q (new_AGEMA_signal_3891) ) ;
    buf_clk new_AGEMA_reg_buffer_2539 ( .C (clk), .D (plaintext_s0[62]), .Q (new_AGEMA_signal_3899) ) ;
    buf_clk new_AGEMA_reg_buffer_2547 ( .C (clk), .D (plaintext_s1[62]), .Q (new_AGEMA_signal_3907) ) ;
    buf_clk new_AGEMA_reg_buffer_2555 ( .C (clk), .D (SelectedKey[48]), .Q (new_AGEMA_signal_3915) ) ;
    buf_clk new_AGEMA_reg_buffer_2563 ( .C (clk), .D (new_AGEMA_signal_1548), .Q (new_AGEMA_signal_3923) ) ;
    buf_clk new_AGEMA_reg_buffer_2571 ( .C (clk), .D (SelectedKey[50]), .Q (new_AGEMA_signal_3931) ) ;
    buf_clk new_AGEMA_reg_buffer_2579 ( .C (clk), .D (new_AGEMA_signal_1554), .Q (new_AGEMA_signal_3939) ) ;
    buf_clk new_AGEMA_reg_buffer_2587 ( .C (clk), .D (SelectedKey[52]), .Q (new_AGEMA_signal_3947) ) ;
    buf_clk new_AGEMA_reg_buffer_2595 ( .C (clk), .D (new_AGEMA_signal_1560), .Q (new_AGEMA_signal_3955) ) ;
    buf_clk new_AGEMA_reg_buffer_2603 ( .C (clk), .D (SelectedKey[54]), .Q (new_AGEMA_signal_3963) ) ;
    buf_clk new_AGEMA_reg_buffer_2611 ( .C (clk), .D (new_AGEMA_signal_1281), .Q (new_AGEMA_signal_3971) ) ;
    buf_clk new_AGEMA_reg_buffer_2619 ( .C (clk), .D (SelectedKey[56]), .Q (new_AGEMA_signal_3979) ) ;
    buf_clk new_AGEMA_reg_buffer_2627 ( .C (clk), .D (new_AGEMA_signal_1284), .Q (new_AGEMA_signal_3987) ) ;
    buf_clk new_AGEMA_reg_buffer_2635 ( .C (clk), .D (SelectedKey[58]), .Q (new_AGEMA_signal_3995) ) ;
    buf_clk new_AGEMA_reg_buffer_2643 ( .C (clk), .D (new_AGEMA_signal_1569), .Q (new_AGEMA_signal_4003) ) ;
    buf_clk new_AGEMA_reg_buffer_2651 ( .C (clk), .D (SelectedKey[60]), .Q (new_AGEMA_signal_4011) ) ;
    buf_clk new_AGEMA_reg_buffer_2659 ( .C (clk), .D (new_AGEMA_signal_1572), .Q (new_AGEMA_signal_4019) ) ;
    buf_clk new_AGEMA_reg_buffer_2667 ( .C (clk), .D (SelectedKey[62]), .Q (new_AGEMA_signal_4027) ) ;
    buf_clk new_AGEMA_reg_buffer_2675 ( .C (clk), .D (new_AGEMA_signal_1290), .Q (new_AGEMA_signal_4035) ) ;
    buf_clk new_AGEMA_reg_buffer_2683 ( .C (clk), .D (AddKeyConstXOR_XORInst_0_0_n1), .Q (new_AGEMA_signal_4043) ) ;
    buf_clk new_AGEMA_reg_buffer_2691 ( .C (clk), .D (new_AGEMA_signal_1707), .Q (new_AGEMA_signal_4051) ) ;
    buf_clk new_AGEMA_reg_buffer_2699 ( .C (clk), .D (AddKeyConstXOR_XORInst_0_2_n1), .Q (new_AGEMA_signal_4059) ) ;
    buf_clk new_AGEMA_reg_buffer_2707 ( .C (clk), .D (new_AGEMA_signal_1709), .Q (new_AGEMA_signal_4067) ) ;
    buf_clk new_AGEMA_reg_buffer_2715 ( .C (clk), .D (AddKeyConstXOR_XORInst_1_0_n1), .Q (new_AGEMA_signal_4075) ) ;
    buf_clk new_AGEMA_reg_buffer_2723 ( .C (clk), .D (new_AGEMA_signal_1711), .Q (new_AGEMA_signal_4083) ) ;
    buf_clk new_AGEMA_reg_buffer_2731 ( .C (clk), .D (AddKeyConstXOR_XORInst_1_2_n1), .Q (new_AGEMA_signal_4091) ) ;
    buf_clk new_AGEMA_reg_buffer_2739 ( .C (clk), .D (new_AGEMA_signal_1713), .Q (new_AGEMA_signal_4099) ) ;
    buf_clk new_AGEMA_reg_buffer_2747 ( .C (clk), .D (SelectedKey[0]), .Q (new_AGEMA_signal_4107) ) ;
    buf_clk new_AGEMA_reg_buffer_2755 ( .C (clk), .D (new_AGEMA_signal_1245), .Q (new_AGEMA_signal_4115) ) ;
    buf_clk new_AGEMA_reg_buffer_2763 ( .C (clk), .D (SelectedKey[2]), .Q (new_AGEMA_signal_4123) ) ;
    buf_clk new_AGEMA_reg_buffer_2771 ( .C (clk), .D (new_AGEMA_signal_1248), .Q (new_AGEMA_signal_4131) ) ;
    buf_clk new_AGEMA_reg_buffer_2779 ( .C (clk), .D (SelectedKey[4]), .Q (new_AGEMA_signal_4139) ) ;
    buf_clk new_AGEMA_reg_buffer_2787 ( .C (clk), .D (new_AGEMA_signal_1443), .Q (new_AGEMA_signal_4147) ) ;
    buf_clk new_AGEMA_reg_buffer_2795 ( .C (clk), .D (SelectedKey[6]), .Q (new_AGEMA_signal_4155) ) ;
    buf_clk new_AGEMA_reg_buffer_2803 ( .C (clk), .D (new_AGEMA_signal_1449), .Q (new_AGEMA_signal_4163) ) ;
    buf_clk new_AGEMA_reg_buffer_2811 ( .C (clk), .D (SelectedKey[8]), .Q (new_AGEMA_signal_4171) ) ;
    buf_clk new_AGEMA_reg_buffer_2819 ( .C (clk), .D (new_AGEMA_signal_1455), .Q (new_AGEMA_signal_4179) ) ;
    buf_clk new_AGEMA_reg_buffer_2827 ( .C (clk), .D (SelectedKey[10]), .Q (new_AGEMA_signal_4187) ) ;
    buf_clk new_AGEMA_reg_buffer_2835 ( .C (clk), .D (new_AGEMA_signal_1461), .Q (new_AGEMA_signal_4195) ) ;
    buf_clk new_AGEMA_reg_buffer_2843 ( .C (clk), .D (SelectedKey[12]), .Q (new_AGEMA_signal_4203) ) ;
    buf_clk new_AGEMA_reg_buffer_2851 ( .C (clk), .D (new_AGEMA_signal_1467), .Q (new_AGEMA_signal_4211) ) ;
    buf_clk new_AGEMA_reg_buffer_2859 ( .C (clk), .D (SelectedKey[14]), .Q (new_AGEMA_signal_4219) ) ;
    buf_clk new_AGEMA_reg_buffer_2867 ( .C (clk), .D (new_AGEMA_signal_1473), .Q (new_AGEMA_signal_4227) ) ;
    buf_clk new_AGEMA_reg_buffer_2875 ( .C (clk), .D (SelectedKey[16]), .Q (new_AGEMA_signal_4235) ) ;
    buf_clk new_AGEMA_reg_buffer_2883 ( .C (clk), .D (new_AGEMA_signal_1479), .Q (new_AGEMA_signal_4243) ) ;
    buf_clk new_AGEMA_reg_buffer_2891 ( .C (clk), .D (SelectedKey[18]), .Q (new_AGEMA_signal_4251) ) ;
    buf_clk new_AGEMA_reg_buffer_2899 ( .C (clk), .D (new_AGEMA_signal_1485), .Q (new_AGEMA_signal_4259) ) ;
    buf_clk new_AGEMA_reg_buffer_2907 ( .C (clk), .D (SelectedKey[20]), .Q (new_AGEMA_signal_4267) ) ;
    buf_clk new_AGEMA_reg_buffer_2915 ( .C (clk), .D (new_AGEMA_signal_1491), .Q (new_AGEMA_signal_4275) ) ;
    buf_clk new_AGEMA_reg_buffer_2923 ( .C (clk), .D (SelectedKey[22]), .Q (new_AGEMA_signal_4283) ) ;
    buf_clk new_AGEMA_reg_buffer_2931 ( .C (clk), .D (new_AGEMA_signal_1251), .Q (new_AGEMA_signal_4291) ) ;
    buf_clk new_AGEMA_reg_buffer_2939 ( .C (clk), .D (SelectedKey[24]), .Q (new_AGEMA_signal_4299) ) ;
    buf_clk new_AGEMA_reg_buffer_2947 ( .C (clk), .D (new_AGEMA_signal_1257), .Q (new_AGEMA_signal_4307) ) ;
    buf_clk new_AGEMA_reg_buffer_2955 ( .C (clk), .D (SelectedKey[26]), .Q (new_AGEMA_signal_4315) ) ;
    buf_clk new_AGEMA_reg_buffer_2963 ( .C (clk), .D (new_AGEMA_signal_1263), .Q (new_AGEMA_signal_4323) ) ;
    buf_clk new_AGEMA_reg_buffer_2971 ( .C (clk), .D (SelectedKey[28]), .Q (new_AGEMA_signal_4331) ) ;
    buf_clk new_AGEMA_reg_buffer_2979 ( .C (clk), .D (new_AGEMA_signal_1497), .Q (new_AGEMA_signal_4339) ) ;
    buf_clk new_AGEMA_reg_buffer_2987 ( .C (clk), .D (SelectedKey[30]), .Q (new_AGEMA_signal_4347) ) ;
    buf_clk new_AGEMA_reg_buffer_2995 ( .C (clk), .D (new_AGEMA_signal_1503), .Q (new_AGEMA_signal_4355) ) ;
    buf_clk new_AGEMA_reg_buffer_3003 ( .C (clk), .D (SelectedKey[32]), .Q (new_AGEMA_signal_4363) ) ;
    buf_clk new_AGEMA_reg_buffer_3011 ( .C (clk), .D (new_AGEMA_signal_1509), .Q (new_AGEMA_signal_4371) ) ;
    buf_clk new_AGEMA_reg_buffer_3019 ( .C (clk), .D (SelectedKey[34]), .Q (new_AGEMA_signal_4379) ) ;
    buf_clk new_AGEMA_reg_buffer_3027 ( .C (clk), .D (new_AGEMA_signal_1512), .Q (new_AGEMA_signal_4387) ) ;
    buf_clk new_AGEMA_reg_buffer_3035 ( .C (clk), .D (SelectedKey[36]), .Q (new_AGEMA_signal_4395) ) ;
    buf_clk new_AGEMA_reg_buffer_3043 ( .C (clk), .D (new_AGEMA_signal_1272), .Q (new_AGEMA_signal_4403) ) ;
    buf_clk new_AGEMA_reg_buffer_3051 ( .C (clk), .D (SelectedKey[38]), .Q (new_AGEMA_signal_4411) ) ;
    buf_clk new_AGEMA_reg_buffer_3059 ( .C (clk), .D (new_AGEMA_signal_1521), .Q (new_AGEMA_signal_4419) ) ;
    buf_clk new_AGEMA_reg_buffer_3387 ( .C (clk), .D (FSMUpdate[6]), .Q (new_AGEMA_signal_4747) ) ;
    buf_clk new_AGEMA_reg_buffer_3395 ( .C (clk), .D (FSMUpdate[5]), .Q (new_AGEMA_signal_4755) ) ;
    buf_clk new_AGEMA_reg_buffer_3403 ( .C (clk), .D (FSMUpdate[4]), .Q (new_AGEMA_signal_4763) ) ;
    buf_clk new_AGEMA_reg_buffer_3411 ( .C (clk), .D (FSMUpdate[3]), .Q (new_AGEMA_signal_4771) ) ;
    buf_clk new_AGEMA_reg_buffer_3419 ( .C (clk), .D (FSMUpdate[2]), .Q (new_AGEMA_signal_4779) ) ;
    buf_clk new_AGEMA_reg_buffer_3427 ( .C (clk), .D (FSMUpdate[1]), .Q (new_AGEMA_signal_4787) ) ;
    buf_clk new_AGEMA_reg_buffer_3435 ( .C (clk), .D (FSMUpdate[0]), .Q (new_AGEMA_signal_4795) ) ;
    buf_clk new_AGEMA_reg_buffer_3443 ( .C (clk), .D (selectsNext[1]), .Q (new_AGEMA_signal_4803) ) ;
    buf_clk new_AGEMA_reg_buffer_3451 ( .C (clk), .D (selectsNext[0]), .Q (new_AGEMA_signal_4811) ) ;
    buf_clk new_AGEMA_reg_buffer_3459 ( .C (clk), .D (done_internal), .Q (new_AGEMA_signal_4819) ) ;

    /* cells in depth 2 */
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U14 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r (Fresh[0]), .c ({new_AGEMA_signal_1021, SubCellInst_SboxInst_0_n10}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U13 ( .a ({new_AGEMA_signal_1025, SubCellInst_SboxInst_0_n8}), .b ({new_AGEMA_signal_1024, SubCellInst_SboxInst_0_n7}), .clk (clk), .r (Fresh[1]), .c ({new_AGEMA_signal_1148, SubCellInst_SboxInst_0_n15}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U10 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_1026, SubCellInst_SboxInst_0_n9}), .clk (clk), .r (Fresh[2]), .c ({new_AGEMA_signal_1149, SubCellInst_SboxInst_0_n4}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U9 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_1025, SubCellInst_SboxInst_0_n8}), .clk (clk), .r (Fresh[3]), .c ({new_AGEMA_signal_1150, SubCellInst_SboxInst_0_n6}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U5 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r (Fresh[4]), .c ({new_AGEMA_signal_1023, SubCellInst_SboxInst_0_n1}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U3 ( .a ({new_AGEMA_signal_1026, SubCellInst_SboxInst_0_n9}), .b ({new_AGEMA_signal_1025, SubCellInst_SboxInst_0_n8}), .clk (clk), .r (Fresh[5]), .c ({new_AGEMA_signal_1152, SubCellInst_SboxInst_0_n13}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U14 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({ciphertext_s1[51], ciphertext_s0[51]}), .clk (clk), .r (Fresh[6]), .c ({new_AGEMA_signal_1029, SubCellInst_SboxInst_1_n10}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U13 ( .a ({new_AGEMA_signal_1033, SubCellInst_SboxInst_1_n8}), .b ({new_AGEMA_signal_1032, SubCellInst_SboxInst_1_n7}), .clk (clk), .r (Fresh[7]), .c ({new_AGEMA_signal_1154, SubCellInst_SboxInst_1_n15}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U10 ( .a ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({new_AGEMA_signal_1034, SubCellInst_SboxInst_1_n9}), .clk (clk), .r (Fresh[8]), .c ({new_AGEMA_signal_1155, SubCellInst_SboxInst_1_n4}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U9 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_1033, SubCellInst_SboxInst_1_n8}), .clk (clk), .r (Fresh[9]), .c ({new_AGEMA_signal_1156, SubCellInst_SboxInst_1_n6}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U5 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({ciphertext_s1[51], ciphertext_s0[51]}), .clk (clk), .r (Fresh[10]), .c ({new_AGEMA_signal_1031, SubCellInst_SboxInst_1_n1}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U3 ( .a ({new_AGEMA_signal_1034, SubCellInst_SboxInst_1_n9}), .b ({new_AGEMA_signal_1033, SubCellInst_SboxInst_1_n8}), .clk (clk), .r (Fresh[11]), .c ({new_AGEMA_signal_1158, SubCellInst_SboxInst_1_n13}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U14 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r (Fresh[12]), .c ({new_AGEMA_signal_1037, SubCellInst_SboxInst_2_n10}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U13 ( .a ({new_AGEMA_signal_1041, SubCellInst_SboxInst_2_n8}), .b ({new_AGEMA_signal_1040, SubCellInst_SboxInst_2_n7}), .clk (clk), .r (Fresh[13]), .c ({new_AGEMA_signal_1160, SubCellInst_SboxInst_2_n15}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U10 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({new_AGEMA_signal_1042, SubCellInst_SboxInst_2_n9}), .clk (clk), .r (Fresh[14]), .c ({new_AGEMA_signal_1161, SubCellInst_SboxInst_2_n4}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U9 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_1041, SubCellInst_SboxInst_2_n8}), .clk (clk), .r (Fresh[15]), .c ({new_AGEMA_signal_1162, SubCellInst_SboxInst_2_n6}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U5 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r (Fresh[16]), .c ({new_AGEMA_signal_1039, SubCellInst_SboxInst_2_n1}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U3 ( .a ({new_AGEMA_signal_1042, SubCellInst_SboxInst_2_n9}), .b ({new_AGEMA_signal_1041, SubCellInst_SboxInst_2_n8}), .clk (clk), .r (Fresh[17]), .c ({new_AGEMA_signal_1164, SubCellInst_SboxInst_2_n13}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U14 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .clk (clk), .r (Fresh[18]), .c ({new_AGEMA_signal_1045, SubCellInst_SboxInst_3_n10}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U13 ( .a ({new_AGEMA_signal_1049, SubCellInst_SboxInst_3_n8}), .b ({new_AGEMA_signal_1048, SubCellInst_SboxInst_3_n7}), .clk (clk), .r (Fresh[19]), .c ({new_AGEMA_signal_1166, SubCellInst_SboxInst_3_n15}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U10 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_1050, SubCellInst_SboxInst_3_n9}), .clk (clk), .r (Fresh[20]), .c ({new_AGEMA_signal_1167, SubCellInst_SboxInst_3_n4}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U9 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_1049, SubCellInst_SboxInst_3_n8}), .clk (clk), .r (Fresh[21]), .c ({new_AGEMA_signal_1168, SubCellInst_SboxInst_3_n6}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U5 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .clk (clk), .r (Fresh[22]), .c ({new_AGEMA_signal_1047, SubCellInst_SboxInst_3_n1}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U3 ( .a ({new_AGEMA_signal_1050, SubCellInst_SboxInst_3_n9}), .b ({new_AGEMA_signal_1049, SubCellInst_SboxInst_3_n8}), .clk (clk), .r (Fresh[23]), .c ({new_AGEMA_signal_1170, SubCellInst_SboxInst_3_n13}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U14 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({ciphertext_s1[35], ciphertext_s0[35]}), .clk (clk), .r (Fresh[24]), .c ({new_AGEMA_signal_1053, SubCellInst_SboxInst_4_n10}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U13 ( .a ({new_AGEMA_signal_1057, SubCellInst_SboxInst_4_n8}), .b ({new_AGEMA_signal_1056, SubCellInst_SboxInst_4_n7}), .clk (clk), .r (Fresh[25]), .c ({new_AGEMA_signal_1172, SubCellInst_SboxInst_4_n15}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U10 ( .a ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({new_AGEMA_signal_1058, SubCellInst_SboxInst_4_n9}), .clk (clk), .r (Fresh[26]), .c ({new_AGEMA_signal_1173, SubCellInst_SboxInst_4_n4}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U9 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_1057, SubCellInst_SboxInst_4_n8}), .clk (clk), .r (Fresh[27]), .c ({new_AGEMA_signal_1174, SubCellInst_SboxInst_4_n6}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U5 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({ciphertext_s1[35], ciphertext_s0[35]}), .clk (clk), .r (Fresh[28]), .c ({new_AGEMA_signal_1055, SubCellInst_SboxInst_4_n1}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U3 ( .a ({new_AGEMA_signal_1058, SubCellInst_SboxInst_4_n9}), .b ({new_AGEMA_signal_1057, SubCellInst_SboxInst_4_n8}), .clk (clk), .r (Fresh[29]), .c ({new_AGEMA_signal_1176, SubCellInst_SboxInst_4_n13}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U14 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r (Fresh[30]), .c ({new_AGEMA_signal_1061, SubCellInst_SboxInst_5_n10}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U13 ( .a ({new_AGEMA_signal_1065, SubCellInst_SboxInst_5_n8}), .b ({new_AGEMA_signal_1064, SubCellInst_SboxInst_5_n7}), .clk (clk), .r (Fresh[31]), .c ({new_AGEMA_signal_1178, SubCellInst_SboxInst_5_n15}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U10 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({new_AGEMA_signal_1066, SubCellInst_SboxInst_5_n9}), .clk (clk), .r (Fresh[32]), .c ({new_AGEMA_signal_1179, SubCellInst_SboxInst_5_n4}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U9 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_1065, SubCellInst_SboxInst_5_n8}), .clk (clk), .r (Fresh[33]), .c ({new_AGEMA_signal_1180, SubCellInst_SboxInst_5_n6}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U5 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r (Fresh[34]), .c ({new_AGEMA_signal_1063, SubCellInst_SboxInst_5_n1}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U3 ( .a ({new_AGEMA_signal_1066, SubCellInst_SboxInst_5_n9}), .b ({new_AGEMA_signal_1065, SubCellInst_SboxInst_5_n8}), .clk (clk), .r (Fresh[35]), .c ({new_AGEMA_signal_1182, SubCellInst_SboxInst_5_n13}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U14 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({ciphertext_s1[43], ciphertext_s0[43]}), .clk (clk), .r (Fresh[36]), .c ({new_AGEMA_signal_1069, SubCellInst_SboxInst_6_n10}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U13 ( .a ({new_AGEMA_signal_1073, SubCellInst_SboxInst_6_n8}), .b ({new_AGEMA_signal_1072, SubCellInst_SboxInst_6_n7}), .clk (clk), .r (Fresh[37]), .c ({new_AGEMA_signal_1184, SubCellInst_SboxInst_6_n15}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U10 ( .a ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({new_AGEMA_signal_1074, SubCellInst_SboxInst_6_n9}), .clk (clk), .r (Fresh[38]), .c ({new_AGEMA_signal_1185, SubCellInst_SboxInst_6_n4}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U9 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_1073, SubCellInst_SboxInst_6_n8}), .clk (clk), .r (Fresh[39]), .c ({new_AGEMA_signal_1186, SubCellInst_SboxInst_6_n6}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U5 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({ciphertext_s1[43], ciphertext_s0[43]}), .clk (clk), .r (Fresh[40]), .c ({new_AGEMA_signal_1071, SubCellInst_SboxInst_6_n1}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U3 ( .a ({new_AGEMA_signal_1074, SubCellInst_SboxInst_6_n9}), .b ({new_AGEMA_signal_1073, SubCellInst_SboxInst_6_n8}), .clk (clk), .r (Fresh[41]), .c ({new_AGEMA_signal_1188, SubCellInst_SboxInst_6_n13}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U14 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r (Fresh[42]), .c ({new_AGEMA_signal_1077, SubCellInst_SboxInst_7_n10}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U13 ( .a ({new_AGEMA_signal_1081, SubCellInst_SboxInst_7_n8}), .b ({new_AGEMA_signal_1080, SubCellInst_SboxInst_7_n7}), .clk (clk), .r (Fresh[43]), .c ({new_AGEMA_signal_1190, SubCellInst_SboxInst_7_n15}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U10 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({new_AGEMA_signal_1082, SubCellInst_SboxInst_7_n9}), .clk (clk), .r (Fresh[44]), .c ({new_AGEMA_signal_1191, SubCellInst_SboxInst_7_n4}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U9 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_1081, SubCellInst_SboxInst_7_n8}), .clk (clk), .r (Fresh[45]), .c ({new_AGEMA_signal_1192, SubCellInst_SboxInst_7_n6}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U5 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r (Fresh[46]), .c ({new_AGEMA_signal_1079, SubCellInst_SboxInst_7_n1}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U3 ( .a ({new_AGEMA_signal_1082, SubCellInst_SboxInst_7_n9}), .b ({new_AGEMA_signal_1081, SubCellInst_SboxInst_7_n8}), .clk (clk), .r (Fresh[47]), .c ({new_AGEMA_signal_1194, SubCellInst_SboxInst_7_n13}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U14 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({ciphertext_s1[19], ciphertext_s0[19]}), .clk (clk), .r (Fresh[48]), .c ({new_AGEMA_signal_1085, SubCellInst_SboxInst_8_n10}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U13 ( .a ({new_AGEMA_signal_1089, SubCellInst_SboxInst_8_n8}), .b ({new_AGEMA_signal_1088, SubCellInst_SboxInst_8_n7}), .clk (clk), .r (Fresh[49]), .c ({new_AGEMA_signal_1196, SubCellInst_SboxInst_8_n15}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U10 ( .a ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({new_AGEMA_signal_1090, SubCellInst_SboxInst_8_n9}), .clk (clk), .r (Fresh[50]), .c ({new_AGEMA_signal_1197, SubCellInst_SboxInst_8_n4}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U9 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_1089, SubCellInst_SboxInst_8_n8}), .clk (clk), .r (Fresh[51]), .c ({new_AGEMA_signal_1198, SubCellInst_SboxInst_8_n6}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U5 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({ciphertext_s1[19], ciphertext_s0[19]}), .clk (clk), .r (Fresh[52]), .c ({new_AGEMA_signal_1087, SubCellInst_SboxInst_8_n1}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U3 ( .a ({new_AGEMA_signal_1090, SubCellInst_SboxInst_8_n9}), .b ({new_AGEMA_signal_1089, SubCellInst_SboxInst_8_n8}), .clk (clk), .r (Fresh[53]), .c ({new_AGEMA_signal_1200, SubCellInst_SboxInst_8_n13}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U14 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r (Fresh[54]), .c ({new_AGEMA_signal_1093, SubCellInst_SboxInst_9_n10}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U13 ( .a ({new_AGEMA_signal_1097, SubCellInst_SboxInst_9_n8}), .b ({new_AGEMA_signal_1096, SubCellInst_SboxInst_9_n7}), .clk (clk), .r (Fresh[55]), .c ({new_AGEMA_signal_1202, SubCellInst_SboxInst_9_n15}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U10 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_1098, SubCellInst_SboxInst_9_n9}), .clk (clk), .r (Fresh[56]), .c ({new_AGEMA_signal_1203, SubCellInst_SboxInst_9_n4}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U9 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_1097, SubCellInst_SboxInst_9_n8}), .clk (clk), .r (Fresh[57]), .c ({new_AGEMA_signal_1204, SubCellInst_SboxInst_9_n6}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U5 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r (Fresh[58]), .c ({new_AGEMA_signal_1095, SubCellInst_SboxInst_9_n1}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U3 ( .a ({new_AGEMA_signal_1098, SubCellInst_SboxInst_9_n9}), .b ({new_AGEMA_signal_1097, SubCellInst_SboxInst_9_n8}), .clk (clk), .r (Fresh[59]), .c ({new_AGEMA_signal_1206, SubCellInst_SboxInst_9_n13}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U14 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .clk (clk), .r (Fresh[60]), .c ({new_AGEMA_signal_1101, SubCellInst_SboxInst_10_n10}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U13 ( .a ({new_AGEMA_signal_1105, SubCellInst_SboxInst_10_n8}), .b ({new_AGEMA_signal_1104, SubCellInst_SboxInst_10_n7}), .clk (clk), .r (Fresh[61]), .c ({new_AGEMA_signal_1208, SubCellInst_SboxInst_10_n15}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U10 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_1106, SubCellInst_SboxInst_10_n9}), .clk (clk), .r (Fresh[62]), .c ({new_AGEMA_signal_1209, SubCellInst_SboxInst_10_n4}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U9 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_1105, SubCellInst_SboxInst_10_n8}), .clk (clk), .r (Fresh[63]), .c ({new_AGEMA_signal_1210, SubCellInst_SboxInst_10_n6}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U5 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .clk (clk), .r (Fresh[64]), .c ({new_AGEMA_signal_1103, SubCellInst_SboxInst_10_n1}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U3 ( .a ({new_AGEMA_signal_1106, SubCellInst_SboxInst_10_n9}), .b ({new_AGEMA_signal_1105, SubCellInst_SboxInst_10_n8}), .clk (clk), .r (Fresh[65]), .c ({new_AGEMA_signal_1212, SubCellInst_SboxInst_10_n13}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U14 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r (Fresh[66]), .c ({new_AGEMA_signal_1109, SubCellInst_SboxInst_11_n10}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U13 ( .a ({new_AGEMA_signal_1113, SubCellInst_SboxInst_11_n8}), .b ({new_AGEMA_signal_1112, SubCellInst_SboxInst_11_n7}), .clk (clk), .r (Fresh[67]), .c ({new_AGEMA_signal_1214, SubCellInst_SboxInst_11_n15}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U10 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({new_AGEMA_signal_1114, SubCellInst_SboxInst_11_n9}), .clk (clk), .r (Fresh[68]), .c ({new_AGEMA_signal_1215, SubCellInst_SboxInst_11_n4}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U9 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_1113, SubCellInst_SboxInst_11_n8}), .clk (clk), .r (Fresh[69]), .c ({new_AGEMA_signal_1216, SubCellInst_SboxInst_11_n6}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U5 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r (Fresh[70]), .c ({new_AGEMA_signal_1111, SubCellInst_SboxInst_11_n1}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U3 ( .a ({new_AGEMA_signal_1114, SubCellInst_SboxInst_11_n9}), .b ({new_AGEMA_signal_1113, SubCellInst_SboxInst_11_n8}), .clk (clk), .r (Fresh[71]), .c ({new_AGEMA_signal_1218, SubCellInst_SboxInst_11_n13}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U14 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r (Fresh[72]), .c ({new_AGEMA_signal_1117, SubCellInst_SboxInst_12_n10}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U13 ( .a ({new_AGEMA_signal_1121, SubCellInst_SboxInst_12_n8}), .b ({new_AGEMA_signal_1120, SubCellInst_SboxInst_12_n7}), .clk (clk), .r (Fresh[73]), .c ({new_AGEMA_signal_1220, SubCellInst_SboxInst_12_n15}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U10 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({new_AGEMA_signal_1122, SubCellInst_SboxInst_12_n9}), .clk (clk), .r (Fresh[74]), .c ({new_AGEMA_signal_1221, SubCellInst_SboxInst_12_n4}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U9 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_1121, SubCellInst_SboxInst_12_n8}), .clk (clk), .r (Fresh[75]), .c ({new_AGEMA_signal_1222, SubCellInst_SboxInst_12_n6}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U5 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r (Fresh[76]), .c ({new_AGEMA_signal_1119, SubCellInst_SboxInst_12_n1}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U3 ( .a ({new_AGEMA_signal_1122, SubCellInst_SboxInst_12_n9}), .b ({new_AGEMA_signal_1121, SubCellInst_SboxInst_12_n8}), .clk (clk), .r (Fresh[77]), .c ({new_AGEMA_signal_1224, SubCellInst_SboxInst_12_n13}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U14 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({ciphertext_s1[11], ciphertext_s0[11]}), .clk (clk), .r (Fresh[78]), .c ({new_AGEMA_signal_1125, SubCellInst_SboxInst_13_n10}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U13 ( .a ({new_AGEMA_signal_1129, SubCellInst_SboxInst_13_n8}), .b ({new_AGEMA_signal_1128, SubCellInst_SboxInst_13_n7}), .clk (clk), .r (Fresh[79]), .c ({new_AGEMA_signal_1226, SubCellInst_SboxInst_13_n15}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U10 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({new_AGEMA_signal_1130, SubCellInst_SboxInst_13_n9}), .clk (clk), .r (Fresh[80]), .c ({new_AGEMA_signal_1227, SubCellInst_SboxInst_13_n4}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U9 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_1129, SubCellInst_SboxInst_13_n8}), .clk (clk), .r (Fresh[81]), .c ({new_AGEMA_signal_1228, SubCellInst_SboxInst_13_n6}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U5 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({ciphertext_s1[11], ciphertext_s0[11]}), .clk (clk), .r (Fresh[82]), .c ({new_AGEMA_signal_1127, SubCellInst_SboxInst_13_n1}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U3 ( .a ({new_AGEMA_signal_1130, SubCellInst_SboxInst_13_n9}), .b ({new_AGEMA_signal_1129, SubCellInst_SboxInst_13_n8}), .clk (clk), .r (Fresh[83]), .c ({new_AGEMA_signal_1230, SubCellInst_SboxInst_13_n13}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U14 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r (Fresh[84]), .c ({new_AGEMA_signal_1133, SubCellInst_SboxInst_14_n10}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U13 ( .a ({new_AGEMA_signal_1137, SubCellInst_SboxInst_14_n8}), .b ({new_AGEMA_signal_1136, SubCellInst_SboxInst_14_n7}), .clk (clk), .r (Fresh[85]), .c ({new_AGEMA_signal_1232, SubCellInst_SboxInst_14_n15}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U10 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({new_AGEMA_signal_1138, SubCellInst_SboxInst_14_n9}), .clk (clk), .r (Fresh[86]), .c ({new_AGEMA_signal_1233, SubCellInst_SboxInst_14_n4}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U9 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_1137, SubCellInst_SboxInst_14_n8}), .clk (clk), .r (Fresh[87]), .c ({new_AGEMA_signal_1234, SubCellInst_SboxInst_14_n6}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U5 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r (Fresh[88]), .c ({new_AGEMA_signal_1135, SubCellInst_SboxInst_14_n1}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U3 ( .a ({new_AGEMA_signal_1138, SubCellInst_SboxInst_14_n9}), .b ({new_AGEMA_signal_1137, SubCellInst_SboxInst_14_n8}), .clk (clk), .r (Fresh[89]), .c ({new_AGEMA_signal_1236, SubCellInst_SboxInst_14_n13}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U14 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({ciphertext_s1[3], ciphertext_s0[3]}), .clk (clk), .r (Fresh[90]), .c ({new_AGEMA_signal_1141, SubCellInst_SboxInst_15_n10}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U13 ( .a ({new_AGEMA_signal_1145, SubCellInst_SboxInst_15_n8}), .b ({new_AGEMA_signal_1144, SubCellInst_SboxInst_15_n7}), .clk (clk), .r (Fresh[91]), .c ({new_AGEMA_signal_1238, SubCellInst_SboxInst_15_n15}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U10 ( .a ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({new_AGEMA_signal_1146, SubCellInst_SboxInst_15_n9}), .clk (clk), .r (Fresh[92]), .c ({new_AGEMA_signal_1239, SubCellInst_SboxInst_15_n4}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U9 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_1145, SubCellInst_SboxInst_15_n8}), .clk (clk), .r (Fresh[93]), .c ({new_AGEMA_signal_1240, SubCellInst_SboxInst_15_n6}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U5 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({ciphertext_s1[3], ciphertext_s0[3]}), .clk (clk), .r (Fresh[94]), .c ({new_AGEMA_signal_1143, SubCellInst_SboxInst_15_n1}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U3 ( .a ({new_AGEMA_signal_1146, SubCellInst_SboxInst_15_n9}), .b ({new_AGEMA_signal_1145, SubCellInst_SboxInst_15_n8}), .clk (clk), .r (Fresh[95]), .c ({new_AGEMA_signal_1242, SubCellInst_SboxInst_15_n13}) ) ;
    buf_clk new_AGEMA_reg_buffer_820 ( .C (clk), .D (new_AGEMA_signal_2179), .Q (new_AGEMA_signal_2180) ) ;
    buf_clk new_AGEMA_reg_buffer_822 ( .C (clk), .D (new_AGEMA_signal_2181), .Q (new_AGEMA_signal_2182) ) ;
    buf_clk new_AGEMA_reg_buffer_824 ( .C (clk), .D (new_AGEMA_signal_2183), .Q (new_AGEMA_signal_2184) ) ;
    buf_clk new_AGEMA_reg_buffer_826 ( .C (clk), .D (new_AGEMA_signal_2185), .Q (new_AGEMA_signal_2186) ) ;
    buf_clk new_AGEMA_reg_buffer_828 ( .C (clk), .D (new_AGEMA_signal_2187), .Q (new_AGEMA_signal_2188) ) ;
    buf_clk new_AGEMA_reg_buffer_830 ( .C (clk), .D (new_AGEMA_signal_2189), .Q (new_AGEMA_signal_2190) ) ;
    buf_clk new_AGEMA_reg_buffer_832 ( .C (clk), .D (new_AGEMA_signal_2191), .Q (new_AGEMA_signal_2192) ) ;
    buf_clk new_AGEMA_reg_buffer_834 ( .C (clk), .D (new_AGEMA_signal_2193), .Q (new_AGEMA_signal_2194) ) ;
    buf_clk new_AGEMA_reg_buffer_836 ( .C (clk), .D (new_AGEMA_signal_2195), .Q (new_AGEMA_signal_2196) ) ;
    buf_clk new_AGEMA_reg_buffer_838 ( .C (clk), .D (new_AGEMA_signal_2197), .Q (new_AGEMA_signal_2198) ) ;
    buf_clk new_AGEMA_reg_buffer_840 ( .C (clk), .D (new_AGEMA_signal_2199), .Q (new_AGEMA_signal_2200) ) ;
    buf_clk new_AGEMA_reg_buffer_842 ( .C (clk), .D (new_AGEMA_signal_2201), .Q (new_AGEMA_signal_2202) ) ;
    buf_clk new_AGEMA_reg_buffer_844 ( .C (clk), .D (new_AGEMA_signal_2203), .Q (new_AGEMA_signal_2204) ) ;
    buf_clk new_AGEMA_reg_buffer_846 ( .C (clk), .D (new_AGEMA_signal_2205), .Q (new_AGEMA_signal_2206) ) ;
    buf_clk new_AGEMA_reg_buffer_848 ( .C (clk), .D (new_AGEMA_signal_2207), .Q (new_AGEMA_signal_2208) ) ;
    buf_clk new_AGEMA_reg_buffer_850 ( .C (clk), .D (new_AGEMA_signal_2209), .Q (new_AGEMA_signal_2210) ) ;
    buf_clk new_AGEMA_reg_buffer_852 ( .C (clk), .D (new_AGEMA_signal_2211), .Q (new_AGEMA_signal_2212) ) ;
    buf_clk new_AGEMA_reg_buffer_854 ( .C (clk), .D (new_AGEMA_signal_2213), .Q (new_AGEMA_signal_2214) ) ;
    buf_clk new_AGEMA_reg_buffer_856 ( .C (clk), .D (new_AGEMA_signal_2215), .Q (new_AGEMA_signal_2216) ) ;
    buf_clk new_AGEMA_reg_buffer_858 ( .C (clk), .D (new_AGEMA_signal_2217), .Q (new_AGEMA_signal_2218) ) ;
    buf_clk new_AGEMA_reg_buffer_860 ( .C (clk), .D (new_AGEMA_signal_2219), .Q (new_AGEMA_signal_2220) ) ;
    buf_clk new_AGEMA_reg_buffer_862 ( .C (clk), .D (new_AGEMA_signal_2221), .Q (new_AGEMA_signal_2222) ) ;
    buf_clk new_AGEMA_reg_buffer_864 ( .C (clk), .D (new_AGEMA_signal_2223), .Q (new_AGEMA_signal_2224) ) ;
    buf_clk new_AGEMA_reg_buffer_866 ( .C (clk), .D (new_AGEMA_signal_2225), .Q (new_AGEMA_signal_2226) ) ;
    buf_clk new_AGEMA_reg_buffer_868 ( .C (clk), .D (new_AGEMA_signal_2227), .Q (new_AGEMA_signal_2228) ) ;
    buf_clk new_AGEMA_reg_buffer_870 ( .C (clk), .D (new_AGEMA_signal_2229), .Q (new_AGEMA_signal_2230) ) ;
    buf_clk new_AGEMA_reg_buffer_872 ( .C (clk), .D (new_AGEMA_signal_2231), .Q (new_AGEMA_signal_2232) ) ;
    buf_clk new_AGEMA_reg_buffer_874 ( .C (clk), .D (new_AGEMA_signal_2233), .Q (new_AGEMA_signal_2234) ) ;
    buf_clk new_AGEMA_reg_buffer_876 ( .C (clk), .D (new_AGEMA_signal_2235), .Q (new_AGEMA_signal_2236) ) ;
    buf_clk new_AGEMA_reg_buffer_878 ( .C (clk), .D (new_AGEMA_signal_2237), .Q (new_AGEMA_signal_2238) ) ;
    buf_clk new_AGEMA_reg_buffer_880 ( .C (clk), .D (new_AGEMA_signal_2239), .Q (new_AGEMA_signal_2240) ) ;
    buf_clk new_AGEMA_reg_buffer_882 ( .C (clk), .D (new_AGEMA_signal_2241), .Q (new_AGEMA_signal_2242) ) ;
    buf_clk new_AGEMA_reg_buffer_884 ( .C (clk), .D (new_AGEMA_signal_2243), .Q (new_AGEMA_signal_2244) ) ;
    buf_clk new_AGEMA_reg_buffer_886 ( .C (clk), .D (new_AGEMA_signal_2245), .Q (new_AGEMA_signal_2246) ) ;
    buf_clk new_AGEMA_reg_buffer_888 ( .C (clk), .D (new_AGEMA_signal_2247), .Q (new_AGEMA_signal_2248) ) ;
    buf_clk new_AGEMA_reg_buffer_890 ( .C (clk), .D (new_AGEMA_signal_2249), .Q (new_AGEMA_signal_2250) ) ;
    buf_clk new_AGEMA_reg_buffer_892 ( .C (clk), .D (new_AGEMA_signal_2251), .Q (new_AGEMA_signal_2252) ) ;
    buf_clk new_AGEMA_reg_buffer_894 ( .C (clk), .D (new_AGEMA_signal_2253), .Q (new_AGEMA_signal_2254) ) ;
    buf_clk new_AGEMA_reg_buffer_896 ( .C (clk), .D (new_AGEMA_signal_2255), .Q (new_AGEMA_signal_2256) ) ;
    buf_clk new_AGEMA_reg_buffer_898 ( .C (clk), .D (new_AGEMA_signal_2257), .Q (new_AGEMA_signal_2258) ) ;
    buf_clk new_AGEMA_reg_buffer_900 ( .C (clk), .D (new_AGEMA_signal_2259), .Q (new_AGEMA_signal_2260) ) ;
    buf_clk new_AGEMA_reg_buffer_902 ( .C (clk), .D (new_AGEMA_signal_2261), .Q (new_AGEMA_signal_2262) ) ;
    buf_clk new_AGEMA_reg_buffer_904 ( .C (clk), .D (new_AGEMA_signal_2263), .Q (new_AGEMA_signal_2264) ) ;
    buf_clk new_AGEMA_reg_buffer_906 ( .C (clk), .D (new_AGEMA_signal_2265), .Q (new_AGEMA_signal_2266) ) ;
    buf_clk new_AGEMA_reg_buffer_908 ( .C (clk), .D (new_AGEMA_signal_2267), .Q (new_AGEMA_signal_2268) ) ;
    buf_clk new_AGEMA_reg_buffer_910 ( .C (clk), .D (new_AGEMA_signal_2269), .Q (new_AGEMA_signal_2270) ) ;
    buf_clk new_AGEMA_reg_buffer_912 ( .C (clk), .D (new_AGEMA_signal_2271), .Q (new_AGEMA_signal_2272) ) ;
    buf_clk new_AGEMA_reg_buffer_914 ( .C (clk), .D (new_AGEMA_signal_2273), .Q (new_AGEMA_signal_2274) ) ;
    buf_clk new_AGEMA_reg_buffer_916 ( .C (clk), .D (new_AGEMA_signal_2275), .Q (new_AGEMA_signal_2276) ) ;
    buf_clk new_AGEMA_reg_buffer_918 ( .C (clk), .D (new_AGEMA_signal_2277), .Q (new_AGEMA_signal_2278) ) ;
    buf_clk new_AGEMA_reg_buffer_920 ( .C (clk), .D (new_AGEMA_signal_2279), .Q (new_AGEMA_signal_2280) ) ;
    buf_clk new_AGEMA_reg_buffer_922 ( .C (clk), .D (new_AGEMA_signal_2281), .Q (new_AGEMA_signal_2282) ) ;
    buf_clk new_AGEMA_reg_buffer_924 ( .C (clk), .D (new_AGEMA_signal_2283), .Q (new_AGEMA_signal_2284) ) ;
    buf_clk new_AGEMA_reg_buffer_926 ( .C (clk), .D (new_AGEMA_signal_2285), .Q (new_AGEMA_signal_2286) ) ;
    buf_clk new_AGEMA_reg_buffer_928 ( .C (clk), .D (new_AGEMA_signal_2287), .Q (new_AGEMA_signal_2288) ) ;
    buf_clk new_AGEMA_reg_buffer_930 ( .C (clk), .D (new_AGEMA_signal_2289), .Q (new_AGEMA_signal_2290) ) ;
    buf_clk new_AGEMA_reg_buffer_932 ( .C (clk), .D (new_AGEMA_signal_2291), .Q (new_AGEMA_signal_2292) ) ;
    buf_clk new_AGEMA_reg_buffer_934 ( .C (clk), .D (new_AGEMA_signal_2293), .Q (new_AGEMA_signal_2294) ) ;
    buf_clk new_AGEMA_reg_buffer_936 ( .C (clk), .D (new_AGEMA_signal_2295), .Q (new_AGEMA_signal_2296) ) ;
    buf_clk new_AGEMA_reg_buffer_938 ( .C (clk), .D (new_AGEMA_signal_2297), .Q (new_AGEMA_signal_2298) ) ;
    buf_clk new_AGEMA_reg_buffer_940 ( .C (clk), .D (new_AGEMA_signal_2299), .Q (new_AGEMA_signal_2300) ) ;
    buf_clk new_AGEMA_reg_buffer_942 ( .C (clk), .D (new_AGEMA_signal_2301), .Q (new_AGEMA_signal_2302) ) ;
    buf_clk new_AGEMA_reg_buffer_944 ( .C (clk), .D (new_AGEMA_signal_2303), .Q (new_AGEMA_signal_2304) ) ;
    buf_clk new_AGEMA_reg_buffer_946 ( .C (clk), .D (new_AGEMA_signal_2305), .Q (new_AGEMA_signal_2306) ) ;
    buf_clk new_AGEMA_reg_buffer_948 ( .C (clk), .D (new_AGEMA_signal_2307), .Q (new_AGEMA_signal_2308) ) ;
    buf_clk new_AGEMA_reg_buffer_950 ( .C (clk), .D (new_AGEMA_signal_2309), .Q (new_AGEMA_signal_2310) ) ;
    buf_clk new_AGEMA_reg_buffer_952 ( .C (clk), .D (new_AGEMA_signal_2311), .Q (new_AGEMA_signal_2312) ) ;
    buf_clk new_AGEMA_reg_buffer_954 ( .C (clk), .D (new_AGEMA_signal_2313), .Q (new_AGEMA_signal_2314) ) ;
    buf_clk new_AGEMA_reg_buffer_956 ( .C (clk), .D (new_AGEMA_signal_2315), .Q (new_AGEMA_signal_2316) ) ;
    buf_clk new_AGEMA_reg_buffer_958 ( .C (clk), .D (new_AGEMA_signal_2317), .Q (new_AGEMA_signal_2318) ) ;
    buf_clk new_AGEMA_reg_buffer_960 ( .C (clk), .D (new_AGEMA_signal_2319), .Q (new_AGEMA_signal_2320) ) ;
    buf_clk new_AGEMA_reg_buffer_962 ( .C (clk), .D (new_AGEMA_signal_2321), .Q (new_AGEMA_signal_2322) ) ;
    buf_clk new_AGEMA_reg_buffer_964 ( .C (clk), .D (new_AGEMA_signal_2323), .Q (new_AGEMA_signal_2324) ) ;
    buf_clk new_AGEMA_reg_buffer_966 ( .C (clk), .D (new_AGEMA_signal_2325), .Q (new_AGEMA_signal_2326) ) ;
    buf_clk new_AGEMA_reg_buffer_968 ( .C (clk), .D (new_AGEMA_signal_2327), .Q (new_AGEMA_signal_2328) ) ;
    buf_clk new_AGEMA_reg_buffer_970 ( .C (clk), .D (new_AGEMA_signal_2329), .Q (new_AGEMA_signal_2330) ) ;
    buf_clk new_AGEMA_reg_buffer_972 ( .C (clk), .D (new_AGEMA_signal_2331), .Q (new_AGEMA_signal_2332) ) ;
    buf_clk new_AGEMA_reg_buffer_974 ( .C (clk), .D (new_AGEMA_signal_2333), .Q (new_AGEMA_signal_2334) ) ;
    buf_clk new_AGEMA_reg_buffer_976 ( .C (clk), .D (new_AGEMA_signal_2335), .Q (new_AGEMA_signal_2336) ) ;
    buf_clk new_AGEMA_reg_buffer_978 ( .C (clk), .D (new_AGEMA_signal_2337), .Q (new_AGEMA_signal_2338) ) ;
    buf_clk new_AGEMA_reg_buffer_980 ( .C (clk), .D (new_AGEMA_signal_2339), .Q (new_AGEMA_signal_2340) ) ;
    buf_clk new_AGEMA_reg_buffer_982 ( .C (clk), .D (new_AGEMA_signal_2341), .Q (new_AGEMA_signal_2342) ) ;
    buf_clk new_AGEMA_reg_buffer_984 ( .C (clk), .D (new_AGEMA_signal_2343), .Q (new_AGEMA_signal_2344) ) ;
    buf_clk new_AGEMA_reg_buffer_986 ( .C (clk), .D (new_AGEMA_signal_2345), .Q (new_AGEMA_signal_2346) ) ;
    buf_clk new_AGEMA_reg_buffer_988 ( .C (clk), .D (new_AGEMA_signal_2347), .Q (new_AGEMA_signal_2348) ) ;
    buf_clk new_AGEMA_reg_buffer_990 ( .C (clk), .D (new_AGEMA_signal_2349), .Q (new_AGEMA_signal_2350) ) ;
    buf_clk new_AGEMA_reg_buffer_992 ( .C (clk), .D (new_AGEMA_signal_2351), .Q (new_AGEMA_signal_2352) ) ;
    buf_clk new_AGEMA_reg_buffer_994 ( .C (clk), .D (new_AGEMA_signal_2353), .Q (new_AGEMA_signal_2354) ) ;
    buf_clk new_AGEMA_reg_buffer_996 ( .C (clk), .D (new_AGEMA_signal_2355), .Q (new_AGEMA_signal_2356) ) ;
    buf_clk new_AGEMA_reg_buffer_998 ( .C (clk), .D (new_AGEMA_signal_2357), .Q (new_AGEMA_signal_2358) ) ;
    buf_clk new_AGEMA_reg_buffer_1000 ( .C (clk), .D (new_AGEMA_signal_2359), .Q (new_AGEMA_signal_2360) ) ;
    buf_clk new_AGEMA_reg_buffer_1002 ( .C (clk), .D (new_AGEMA_signal_2361), .Q (new_AGEMA_signal_2362) ) ;
    buf_clk new_AGEMA_reg_buffer_1004 ( .C (clk), .D (new_AGEMA_signal_2363), .Q (new_AGEMA_signal_2364) ) ;
    buf_clk new_AGEMA_reg_buffer_1006 ( .C (clk), .D (new_AGEMA_signal_2365), .Q (new_AGEMA_signal_2366) ) ;
    buf_clk new_AGEMA_reg_buffer_1008 ( .C (clk), .D (new_AGEMA_signal_2367), .Q (new_AGEMA_signal_2368) ) ;
    buf_clk new_AGEMA_reg_buffer_1010 ( .C (clk), .D (new_AGEMA_signal_2369), .Q (new_AGEMA_signal_2370) ) ;
    buf_clk new_AGEMA_reg_buffer_1012 ( .C (clk), .D (new_AGEMA_signal_2371), .Q (new_AGEMA_signal_2372) ) ;
    buf_clk new_AGEMA_reg_buffer_1014 ( .C (clk), .D (new_AGEMA_signal_2373), .Q (new_AGEMA_signal_2374) ) ;
    buf_clk new_AGEMA_reg_buffer_1016 ( .C (clk), .D (new_AGEMA_signal_2375), .Q (new_AGEMA_signal_2376) ) ;
    buf_clk new_AGEMA_reg_buffer_1018 ( .C (clk), .D (new_AGEMA_signal_2377), .Q (new_AGEMA_signal_2378) ) ;
    buf_clk new_AGEMA_reg_buffer_1020 ( .C (clk), .D (new_AGEMA_signal_2379), .Q (new_AGEMA_signal_2380) ) ;
    buf_clk new_AGEMA_reg_buffer_1022 ( .C (clk), .D (new_AGEMA_signal_2381), .Q (new_AGEMA_signal_2382) ) ;
    buf_clk new_AGEMA_reg_buffer_1024 ( .C (clk), .D (new_AGEMA_signal_2383), .Q (new_AGEMA_signal_2384) ) ;
    buf_clk new_AGEMA_reg_buffer_1026 ( .C (clk), .D (new_AGEMA_signal_2385), .Q (new_AGEMA_signal_2386) ) ;
    buf_clk new_AGEMA_reg_buffer_1028 ( .C (clk), .D (new_AGEMA_signal_2387), .Q (new_AGEMA_signal_2388) ) ;
    buf_clk new_AGEMA_reg_buffer_1030 ( .C (clk), .D (new_AGEMA_signal_2389), .Q (new_AGEMA_signal_2390) ) ;
    buf_clk new_AGEMA_reg_buffer_1032 ( .C (clk), .D (new_AGEMA_signal_2391), .Q (new_AGEMA_signal_2392) ) ;
    buf_clk new_AGEMA_reg_buffer_1034 ( .C (clk), .D (new_AGEMA_signal_2393), .Q (new_AGEMA_signal_2394) ) ;
    buf_clk new_AGEMA_reg_buffer_1036 ( .C (clk), .D (new_AGEMA_signal_2395), .Q (new_AGEMA_signal_2396) ) ;
    buf_clk new_AGEMA_reg_buffer_1038 ( .C (clk), .D (new_AGEMA_signal_2397), .Q (new_AGEMA_signal_2398) ) ;
    buf_clk new_AGEMA_reg_buffer_1040 ( .C (clk), .D (new_AGEMA_signal_2399), .Q (new_AGEMA_signal_2400) ) ;
    buf_clk new_AGEMA_reg_buffer_1042 ( .C (clk), .D (new_AGEMA_signal_2401), .Q (new_AGEMA_signal_2402) ) ;
    buf_clk new_AGEMA_reg_buffer_1044 ( .C (clk), .D (new_AGEMA_signal_2403), .Q (new_AGEMA_signal_2404) ) ;
    buf_clk new_AGEMA_reg_buffer_1046 ( .C (clk), .D (new_AGEMA_signal_2405), .Q (new_AGEMA_signal_2406) ) ;
    buf_clk new_AGEMA_reg_buffer_1048 ( .C (clk), .D (new_AGEMA_signal_2407), .Q (new_AGEMA_signal_2408) ) ;
    buf_clk new_AGEMA_reg_buffer_1050 ( .C (clk), .D (new_AGEMA_signal_2409), .Q (new_AGEMA_signal_2410) ) ;
    buf_clk new_AGEMA_reg_buffer_1052 ( .C (clk), .D (new_AGEMA_signal_2411), .Q (new_AGEMA_signal_2412) ) ;
    buf_clk new_AGEMA_reg_buffer_1054 ( .C (clk), .D (new_AGEMA_signal_2413), .Q (new_AGEMA_signal_2414) ) ;
    buf_clk new_AGEMA_reg_buffer_1056 ( .C (clk), .D (new_AGEMA_signal_2415), .Q (new_AGEMA_signal_2416) ) ;
    buf_clk new_AGEMA_reg_buffer_1058 ( .C (clk), .D (new_AGEMA_signal_2417), .Q (new_AGEMA_signal_2418) ) ;
    buf_clk new_AGEMA_reg_buffer_1060 ( .C (clk), .D (new_AGEMA_signal_2419), .Q (new_AGEMA_signal_2420) ) ;
    buf_clk new_AGEMA_reg_buffer_1062 ( .C (clk), .D (new_AGEMA_signal_2421), .Q (new_AGEMA_signal_2422) ) ;
    buf_clk new_AGEMA_reg_buffer_1064 ( .C (clk), .D (new_AGEMA_signal_2423), .Q (new_AGEMA_signal_2424) ) ;
    buf_clk new_AGEMA_reg_buffer_1066 ( .C (clk), .D (new_AGEMA_signal_2425), .Q (new_AGEMA_signal_2426) ) ;
    buf_clk new_AGEMA_reg_buffer_1068 ( .C (clk), .D (new_AGEMA_signal_2427), .Q (new_AGEMA_signal_2428) ) ;
    buf_clk new_AGEMA_reg_buffer_1070 ( .C (clk), .D (new_AGEMA_signal_2429), .Q (new_AGEMA_signal_2430) ) ;
    buf_clk new_AGEMA_reg_buffer_1072 ( .C (clk), .D (new_AGEMA_signal_2431), .Q (new_AGEMA_signal_2432) ) ;
    buf_clk new_AGEMA_reg_buffer_1074 ( .C (clk), .D (new_AGEMA_signal_2433), .Q (new_AGEMA_signal_2434) ) ;
    buf_clk new_AGEMA_reg_buffer_1076 ( .C (clk), .D (new_AGEMA_signal_2435), .Q (new_AGEMA_signal_2436) ) ;
    buf_clk new_AGEMA_reg_buffer_1082 ( .C (clk), .D (new_AGEMA_signal_2441), .Q (new_AGEMA_signal_2442) ) ;
    buf_clk new_AGEMA_reg_buffer_1088 ( .C (clk), .D (new_AGEMA_signal_2447), .Q (new_AGEMA_signal_2448) ) ;
    buf_clk new_AGEMA_reg_buffer_1094 ( .C (clk), .D (new_AGEMA_signal_2453), .Q (new_AGEMA_signal_2454) ) ;
    buf_clk new_AGEMA_reg_buffer_1100 ( .C (clk), .D (new_AGEMA_signal_2459), .Q (new_AGEMA_signal_2460) ) ;
    buf_clk new_AGEMA_reg_buffer_1106 ( .C (clk), .D (new_AGEMA_signal_2465), .Q (new_AGEMA_signal_2466) ) ;
    buf_clk new_AGEMA_reg_buffer_1112 ( .C (clk), .D (new_AGEMA_signal_2471), .Q (new_AGEMA_signal_2472) ) ;
    buf_clk new_AGEMA_reg_buffer_1118 ( .C (clk), .D (new_AGEMA_signal_2477), .Q (new_AGEMA_signal_2478) ) ;
    buf_clk new_AGEMA_reg_buffer_1124 ( .C (clk), .D (new_AGEMA_signal_2483), .Q (new_AGEMA_signal_2484) ) ;
    buf_clk new_AGEMA_reg_buffer_1130 ( .C (clk), .D (new_AGEMA_signal_2489), .Q (new_AGEMA_signal_2490) ) ;
    buf_clk new_AGEMA_reg_buffer_1136 ( .C (clk), .D (new_AGEMA_signal_2495), .Q (new_AGEMA_signal_2496) ) ;
    buf_clk new_AGEMA_reg_buffer_1142 ( .C (clk), .D (new_AGEMA_signal_2501), .Q (new_AGEMA_signal_2502) ) ;
    buf_clk new_AGEMA_reg_buffer_1148 ( .C (clk), .D (new_AGEMA_signal_2507), .Q (new_AGEMA_signal_2508) ) ;
    buf_clk new_AGEMA_reg_buffer_1154 ( .C (clk), .D (new_AGEMA_signal_2513), .Q (new_AGEMA_signal_2514) ) ;
    buf_clk new_AGEMA_reg_buffer_1160 ( .C (clk), .D (new_AGEMA_signal_2519), .Q (new_AGEMA_signal_2520) ) ;
    buf_clk new_AGEMA_reg_buffer_1166 ( .C (clk), .D (new_AGEMA_signal_2525), .Q (new_AGEMA_signal_2526) ) ;
    buf_clk new_AGEMA_reg_buffer_1172 ( .C (clk), .D (new_AGEMA_signal_2531), .Q (new_AGEMA_signal_2532) ) ;
    buf_clk new_AGEMA_reg_buffer_1178 ( .C (clk), .D (new_AGEMA_signal_2537), .Q (new_AGEMA_signal_2538) ) ;
    buf_clk new_AGEMA_reg_buffer_1184 ( .C (clk), .D (new_AGEMA_signal_2543), .Q (new_AGEMA_signal_2544) ) ;
    buf_clk new_AGEMA_reg_buffer_1190 ( .C (clk), .D (new_AGEMA_signal_2549), .Q (new_AGEMA_signal_2550) ) ;
    buf_clk new_AGEMA_reg_buffer_1196 ( .C (clk), .D (new_AGEMA_signal_2555), .Q (new_AGEMA_signal_2556) ) ;
    buf_clk new_AGEMA_reg_buffer_1202 ( .C (clk), .D (new_AGEMA_signal_2561), .Q (new_AGEMA_signal_2562) ) ;
    buf_clk new_AGEMA_reg_buffer_1208 ( .C (clk), .D (new_AGEMA_signal_2567), .Q (new_AGEMA_signal_2568) ) ;
    buf_clk new_AGEMA_reg_buffer_1214 ( .C (clk), .D (new_AGEMA_signal_2573), .Q (new_AGEMA_signal_2574) ) ;
    buf_clk new_AGEMA_reg_buffer_1220 ( .C (clk), .D (new_AGEMA_signal_2579), .Q (new_AGEMA_signal_2580) ) ;
    buf_clk new_AGEMA_reg_buffer_1226 ( .C (clk), .D (new_AGEMA_signal_2585), .Q (new_AGEMA_signal_2586) ) ;
    buf_clk new_AGEMA_reg_buffer_1232 ( .C (clk), .D (new_AGEMA_signal_2591), .Q (new_AGEMA_signal_2592) ) ;
    buf_clk new_AGEMA_reg_buffer_1238 ( .C (clk), .D (new_AGEMA_signal_2597), .Q (new_AGEMA_signal_2598) ) ;
    buf_clk new_AGEMA_reg_buffer_1244 ( .C (clk), .D (new_AGEMA_signal_2603), .Q (new_AGEMA_signal_2604) ) ;
    buf_clk new_AGEMA_reg_buffer_1250 ( .C (clk), .D (new_AGEMA_signal_2609), .Q (new_AGEMA_signal_2610) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C (clk), .D (new_AGEMA_signal_2615), .Q (new_AGEMA_signal_2616) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C (clk), .D (new_AGEMA_signal_2621), .Q (new_AGEMA_signal_2622) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C (clk), .D (new_AGEMA_signal_2627), .Q (new_AGEMA_signal_2628) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C (clk), .D (new_AGEMA_signal_2633), .Q (new_AGEMA_signal_2634) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C (clk), .D (new_AGEMA_signal_2639), .Q (new_AGEMA_signal_2640) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C (clk), .D (new_AGEMA_signal_2645), .Q (new_AGEMA_signal_2646) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C (clk), .D (new_AGEMA_signal_2651), .Q (new_AGEMA_signal_2652) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C (clk), .D (new_AGEMA_signal_2657), .Q (new_AGEMA_signal_2658) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C (clk), .D (new_AGEMA_signal_2663), .Q (new_AGEMA_signal_2664) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C (clk), .D (new_AGEMA_signal_2669), .Q (new_AGEMA_signal_2670) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C (clk), .D (new_AGEMA_signal_2675), .Q (new_AGEMA_signal_2676) ) ;
    buf_clk new_AGEMA_reg_buffer_1322 ( .C (clk), .D (new_AGEMA_signal_2681), .Q (new_AGEMA_signal_2682) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C (clk), .D (new_AGEMA_signal_2687), .Q (new_AGEMA_signal_2688) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C (clk), .D (new_AGEMA_signal_2693), .Q (new_AGEMA_signal_2694) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C (clk), .D (new_AGEMA_signal_2699), .Q (new_AGEMA_signal_2700) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C (clk), .D (new_AGEMA_signal_2705), .Q (new_AGEMA_signal_2706) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C (clk), .D (new_AGEMA_signal_2711), .Q (new_AGEMA_signal_2712) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C (clk), .D (new_AGEMA_signal_2717), .Q (new_AGEMA_signal_2718) ) ;
    buf_clk new_AGEMA_reg_buffer_1364 ( .C (clk), .D (new_AGEMA_signal_2723), .Q (new_AGEMA_signal_2724) ) ;
    buf_clk new_AGEMA_reg_buffer_1370 ( .C (clk), .D (new_AGEMA_signal_2729), .Q (new_AGEMA_signal_2730) ) ;
    buf_clk new_AGEMA_reg_buffer_1376 ( .C (clk), .D (new_AGEMA_signal_2735), .Q (new_AGEMA_signal_2736) ) ;
    buf_clk new_AGEMA_reg_buffer_1382 ( .C (clk), .D (new_AGEMA_signal_2741), .Q (new_AGEMA_signal_2742) ) ;
    buf_clk new_AGEMA_reg_buffer_1388 ( .C (clk), .D (new_AGEMA_signal_2747), .Q (new_AGEMA_signal_2748) ) ;
    buf_clk new_AGEMA_reg_buffer_1394 ( .C (clk), .D (new_AGEMA_signal_2753), .Q (new_AGEMA_signal_2754) ) ;
    buf_clk new_AGEMA_reg_buffer_1400 ( .C (clk), .D (new_AGEMA_signal_2759), .Q (new_AGEMA_signal_2760) ) ;
    buf_clk new_AGEMA_reg_buffer_1406 ( .C (clk), .D (new_AGEMA_signal_2765), .Q (new_AGEMA_signal_2766) ) ;
    buf_clk new_AGEMA_reg_buffer_1412 ( .C (clk), .D (new_AGEMA_signal_2771), .Q (new_AGEMA_signal_2772) ) ;
    buf_clk new_AGEMA_reg_buffer_1418 ( .C (clk), .D (new_AGEMA_signal_2777), .Q (new_AGEMA_signal_2778) ) ;
    buf_clk new_AGEMA_reg_buffer_1424 ( .C (clk), .D (new_AGEMA_signal_2783), .Q (new_AGEMA_signal_2784) ) ;
    buf_clk new_AGEMA_reg_buffer_1430 ( .C (clk), .D (new_AGEMA_signal_2789), .Q (new_AGEMA_signal_2790) ) ;
    buf_clk new_AGEMA_reg_buffer_1436 ( .C (clk), .D (new_AGEMA_signal_2795), .Q (new_AGEMA_signal_2796) ) ;
    buf_clk new_AGEMA_reg_buffer_1442 ( .C (clk), .D (new_AGEMA_signal_2801), .Q (new_AGEMA_signal_2802) ) ;
    buf_clk new_AGEMA_reg_buffer_1448 ( .C (clk), .D (new_AGEMA_signal_2807), .Q (new_AGEMA_signal_2808) ) ;
    buf_clk new_AGEMA_reg_buffer_1454 ( .C (clk), .D (new_AGEMA_signal_2813), .Q (new_AGEMA_signal_2814) ) ;
    buf_clk new_AGEMA_reg_buffer_1460 ( .C (clk), .D (new_AGEMA_signal_2819), .Q (new_AGEMA_signal_2820) ) ;
    buf_clk new_AGEMA_reg_buffer_1466 ( .C (clk), .D (new_AGEMA_signal_2825), .Q (new_AGEMA_signal_2826) ) ;
    buf_clk new_AGEMA_reg_buffer_1472 ( .C (clk), .D (new_AGEMA_signal_2831), .Q (new_AGEMA_signal_2832) ) ;
    buf_clk new_AGEMA_reg_buffer_1478 ( .C (clk), .D (new_AGEMA_signal_2837), .Q (new_AGEMA_signal_2838) ) ;
    buf_clk new_AGEMA_reg_buffer_1484 ( .C (clk), .D (new_AGEMA_signal_2843), .Q (new_AGEMA_signal_2844) ) ;
    buf_clk new_AGEMA_reg_buffer_1490 ( .C (clk), .D (new_AGEMA_signal_2849), .Q (new_AGEMA_signal_2850) ) ;
    buf_clk new_AGEMA_reg_buffer_1496 ( .C (clk), .D (new_AGEMA_signal_2855), .Q (new_AGEMA_signal_2856) ) ;
    buf_clk new_AGEMA_reg_buffer_1502 ( .C (clk), .D (new_AGEMA_signal_2861), .Q (new_AGEMA_signal_2862) ) ;
    buf_clk new_AGEMA_reg_buffer_1508 ( .C (clk), .D (new_AGEMA_signal_2867), .Q (new_AGEMA_signal_2868) ) ;
    buf_clk new_AGEMA_reg_buffer_1514 ( .C (clk), .D (new_AGEMA_signal_2873), .Q (new_AGEMA_signal_2874) ) ;
    buf_clk new_AGEMA_reg_buffer_1520 ( .C (clk), .D (new_AGEMA_signal_2879), .Q (new_AGEMA_signal_2880) ) ;
    buf_clk new_AGEMA_reg_buffer_1526 ( .C (clk), .D (new_AGEMA_signal_2885), .Q (new_AGEMA_signal_2886) ) ;
    buf_clk new_AGEMA_reg_buffer_1532 ( .C (clk), .D (new_AGEMA_signal_2891), .Q (new_AGEMA_signal_2892) ) ;
    buf_clk new_AGEMA_reg_buffer_1538 ( .C (clk), .D (new_AGEMA_signal_2897), .Q (new_AGEMA_signal_2898) ) ;
    buf_clk new_AGEMA_reg_buffer_1544 ( .C (clk), .D (new_AGEMA_signal_2903), .Q (new_AGEMA_signal_2904) ) ;
    buf_clk new_AGEMA_reg_buffer_1550 ( .C (clk), .D (new_AGEMA_signal_2909), .Q (new_AGEMA_signal_2910) ) ;
    buf_clk new_AGEMA_reg_buffer_1556 ( .C (clk), .D (new_AGEMA_signal_2915), .Q (new_AGEMA_signal_2916) ) ;
    buf_clk new_AGEMA_reg_buffer_1562 ( .C (clk), .D (new_AGEMA_signal_2921), .Q (new_AGEMA_signal_2922) ) ;
    buf_clk new_AGEMA_reg_buffer_1568 ( .C (clk), .D (new_AGEMA_signal_2927), .Q (new_AGEMA_signal_2928) ) ;
    buf_clk new_AGEMA_reg_buffer_1574 ( .C (clk), .D (new_AGEMA_signal_2933), .Q (new_AGEMA_signal_2934) ) ;
    buf_clk new_AGEMA_reg_buffer_1580 ( .C (clk), .D (new_AGEMA_signal_2939), .Q (new_AGEMA_signal_2940) ) ;
    buf_clk new_AGEMA_reg_buffer_1586 ( .C (clk), .D (new_AGEMA_signal_2945), .Q (new_AGEMA_signal_2946) ) ;
    buf_clk new_AGEMA_reg_buffer_1592 ( .C (clk), .D (new_AGEMA_signal_2951), .Q (new_AGEMA_signal_2952) ) ;
    buf_clk new_AGEMA_reg_buffer_1598 ( .C (clk), .D (new_AGEMA_signal_2957), .Q (new_AGEMA_signal_2958) ) ;
    buf_clk new_AGEMA_reg_buffer_1604 ( .C (clk), .D (new_AGEMA_signal_2963), .Q (new_AGEMA_signal_2964) ) ;
    buf_clk new_AGEMA_reg_buffer_1610 ( .C (clk), .D (new_AGEMA_signal_2969), .Q (new_AGEMA_signal_2970) ) ;
    buf_clk new_AGEMA_reg_buffer_1616 ( .C (clk), .D (new_AGEMA_signal_2975), .Q (new_AGEMA_signal_2976) ) ;
    buf_clk new_AGEMA_reg_buffer_1622 ( .C (clk), .D (new_AGEMA_signal_2981), .Q (new_AGEMA_signal_2982) ) ;
    buf_clk new_AGEMA_reg_buffer_1628 ( .C (clk), .D (new_AGEMA_signal_2987), .Q (new_AGEMA_signal_2988) ) ;
    buf_clk new_AGEMA_reg_buffer_1634 ( .C (clk), .D (new_AGEMA_signal_2993), .Q (new_AGEMA_signal_2994) ) ;
    buf_clk new_AGEMA_reg_buffer_1640 ( .C (clk), .D (new_AGEMA_signal_2999), .Q (new_AGEMA_signal_3000) ) ;
    buf_clk new_AGEMA_reg_buffer_1646 ( .C (clk), .D (new_AGEMA_signal_3005), .Q (new_AGEMA_signal_3006) ) ;
    buf_clk new_AGEMA_reg_buffer_1652 ( .C (clk), .D (new_AGEMA_signal_3011), .Q (new_AGEMA_signal_3012) ) ;
    buf_clk new_AGEMA_reg_buffer_1658 ( .C (clk), .D (new_AGEMA_signal_3017), .Q (new_AGEMA_signal_3018) ) ;
    buf_clk new_AGEMA_reg_buffer_1664 ( .C (clk), .D (new_AGEMA_signal_3023), .Q (new_AGEMA_signal_3024) ) ;
    buf_clk new_AGEMA_reg_buffer_1670 ( .C (clk), .D (new_AGEMA_signal_3029), .Q (new_AGEMA_signal_3030) ) ;
    buf_clk new_AGEMA_reg_buffer_1676 ( .C (clk), .D (new_AGEMA_signal_3035), .Q (new_AGEMA_signal_3036) ) ;
    buf_clk new_AGEMA_reg_buffer_1682 ( .C (clk), .D (new_AGEMA_signal_3041), .Q (new_AGEMA_signal_3042) ) ;
    buf_clk new_AGEMA_reg_buffer_1688 ( .C (clk), .D (new_AGEMA_signal_3047), .Q (new_AGEMA_signal_3048) ) ;
    buf_clk new_AGEMA_reg_buffer_1694 ( .C (clk), .D (new_AGEMA_signal_3053), .Q (new_AGEMA_signal_3054) ) ;
    buf_clk new_AGEMA_reg_buffer_1700 ( .C (clk), .D (new_AGEMA_signal_3059), .Q (new_AGEMA_signal_3060) ) ;
    buf_clk new_AGEMA_reg_buffer_1706 ( .C (clk), .D (new_AGEMA_signal_3065), .Q (new_AGEMA_signal_3066) ) ;
    buf_clk new_AGEMA_reg_buffer_1712 ( .C (clk), .D (new_AGEMA_signal_3071), .Q (new_AGEMA_signal_3072) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C (clk), .D (new_AGEMA_signal_3077), .Q (new_AGEMA_signal_3078) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C (clk), .D (new_AGEMA_signal_3083), .Q (new_AGEMA_signal_3084) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C (clk), .D (new_AGEMA_signal_3089), .Q (new_AGEMA_signal_3090) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C (clk), .D (new_AGEMA_signal_3095), .Q (new_AGEMA_signal_3096) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C (clk), .D (new_AGEMA_signal_3101), .Q (new_AGEMA_signal_3102) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C (clk), .D (new_AGEMA_signal_3107), .Q (new_AGEMA_signal_3108) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C (clk), .D (new_AGEMA_signal_3113), .Q (new_AGEMA_signal_3114) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C (clk), .D (new_AGEMA_signal_3119), .Q (new_AGEMA_signal_3120) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C (clk), .D (new_AGEMA_signal_3125), .Q (new_AGEMA_signal_3126) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C (clk), .D (new_AGEMA_signal_3131), .Q (new_AGEMA_signal_3132) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C (clk), .D (new_AGEMA_signal_3137), .Q (new_AGEMA_signal_3138) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C (clk), .D (new_AGEMA_signal_3143), .Q (new_AGEMA_signal_3144) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C (clk), .D (new_AGEMA_signal_3149), .Q (new_AGEMA_signal_3150) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C (clk), .D (new_AGEMA_signal_3155), .Q (new_AGEMA_signal_3156) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C (clk), .D (new_AGEMA_signal_3161), .Q (new_AGEMA_signal_3162) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C (clk), .D (new_AGEMA_signal_3167), .Q (new_AGEMA_signal_3168) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C (clk), .D (new_AGEMA_signal_3173), .Q (new_AGEMA_signal_3174) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C (clk), .D (new_AGEMA_signal_3179), .Q (new_AGEMA_signal_3180) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C (clk), .D (new_AGEMA_signal_3185), .Q (new_AGEMA_signal_3186) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C (clk), .D (new_AGEMA_signal_3191), .Q (new_AGEMA_signal_3192) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C (clk), .D (new_AGEMA_signal_3197), .Q (new_AGEMA_signal_3198) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C (clk), .D (new_AGEMA_signal_3203), .Q (new_AGEMA_signal_3204) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C (clk), .D (new_AGEMA_signal_3403), .Q (new_AGEMA_signal_3404) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C (clk), .D (new_AGEMA_signal_3411), .Q (new_AGEMA_signal_3412) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C (clk), .D (new_AGEMA_signal_3419), .Q (new_AGEMA_signal_3420) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C (clk), .D (new_AGEMA_signal_3427), .Q (new_AGEMA_signal_3428) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C (clk), .D (new_AGEMA_signal_3435), .Q (new_AGEMA_signal_3436) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C (clk), .D (new_AGEMA_signal_3443), .Q (new_AGEMA_signal_3444) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C (clk), .D (new_AGEMA_signal_3451), .Q (new_AGEMA_signal_3452) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C (clk), .D (new_AGEMA_signal_3459), .Q (new_AGEMA_signal_3460) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C (clk), .D (new_AGEMA_signal_3467), .Q (new_AGEMA_signal_3468) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C (clk), .D (new_AGEMA_signal_3475), .Q (new_AGEMA_signal_3476) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C (clk), .D (new_AGEMA_signal_3483), .Q (new_AGEMA_signal_3484) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C (clk), .D (new_AGEMA_signal_3491), .Q (new_AGEMA_signal_3492) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C (clk), .D (new_AGEMA_signal_3499), .Q (new_AGEMA_signal_3500) ) ;
    buf_clk new_AGEMA_reg_buffer_2148 ( .C (clk), .D (new_AGEMA_signal_3507), .Q (new_AGEMA_signal_3508) ) ;
    buf_clk new_AGEMA_reg_buffer_2156 ( .C (clk), .D (new_AGEMA_signal_3515), .Q (new_AGEMA_signal_3516) ) ;
    buf_clk new_AGEMA_reg_buffer_2164 ( .C (clk), .D (new_AGEMA_signal_3523), .Q (new_AGEMA_signal_3524) ) ;
    buf_clk new_AGEMA_reg_buffer_2172 ( .C (clk), .D (new_AGEMA_signal_3531), .Q (new_AGEMA_signal_3532) ) ;
    buf_clk new_AGEMA_reg_buffer_2180 ( .C (clk), .D (new_AGEMA_signal_3539), .Q (new_AGEMA_signal_3540) ) ;
    buf_clk new_AGEMA_reg_buffer_2188 ( .C (clk), .D (new_AGEMA_signal_3547), .Q (new_AGEMA_signal_3548) ) ;
    buf_clk new_AGEMA_reg_buffer_2196 ( .C (clk), .D (new_AGEMA_signal_3555), .Q (new_AGEMA_signal_3556) ) ;
    buf_clk new_AGEMA_reg_buffer_2204 ( .C (clk), .D (new_AGEMA_signal_3563), .Q (new_AGEMA_signal_3564) ) ;
    buf_clk new_AGEMA_reg_buffer_2212 ( .C (clk), .D (new_AGEMA_signal_3571), .Q (new_AGEMA_signal_3572) ) ;
    buf_clk new_AGEMA_reg_buffer_2220 ( .C (clk), .D (new_AGEMA_signal_3579), .Q (new_AGEMA_signal_3580) ) ;
    buf_clk new_AGEMA_reg_buffer_2228 ( .C (clk), .D (new_AGEMA_signal_3587), .Q (new_AGEMA_signal_3588) ) ;
    buf_clk new_AGEMA_reg_buffer_2236 ( .C (clk), .D (new_AGEMA_signal_3595), .Q (new_AGEMA_signal_3596) ) ;
    buf_clk new_AGEMA_reg_buffer_2244 ( .C (clk), .D (new_AGEMA_signal_3603), .Q (new_AGEMA_signal_3604) ) ;
    buf_clk new_AGEMA_reg_buffer_2252 ( .C (clk), .D (new_AGEMA_signal_3611), .Q (new_AGEMA_signal_3612) ) ;
    buf_clk new_AGEMA_reg_buffer_2260 ( .C (clk), .D (new_AGEMA_signal_3619), .Q (new_AGEMA_signal_3620) ) ;
    buf_clk new_AGEMA_reg_buffer_2268 ( .C (clk), .D (new_AGEMA_signal_3627), .Q (new_AGEMA_signal_3628) ) ;
    buf_clk new_AGEMA_reg_buffer_2276 ( .C (clk), .D (new_AGEMA_signal_3635), .Q (new_AGEMA_signal_3636) ) ;
    buf_clk new_AGEMA_reg_buffer_2284 ( .C (clk), .D (new_AGEMA_signal_3643), .Q (new_AGEMA_signal_3644) ) ;
    buf_clk new_AGEMA_reg_buffer_2292 ( .C (clk), .D (new_AGEMA_signal_3651), .Q (new_AGEMA_signal_3652) ) ;
    buf_clk new_AGEMA_reg_buffer_2300 ( .C (clk), .D (new_AGEMA_signal_3659), .Q (new_AGEMA_signal_3660) ) ;
    buf_clk new_AGEMA_reg_buffer_2308 ( .C (clk), .D (new_AGEMA_signal_3667), .Q (new_AGEMA_signal_3668) ) ;
    buf_clk new_AGEMA_reg_buffer_2316 ( .C (clk), .D (new_AGEMA_signal_3675), .Q (new_AGEMA_signal_3676) ) ;
    buf_clk new_AGEMA_reg_buffer_2324 ( .C (clk), .D (new_AGEMA_signal_3683), .Q (new_AGEMA_signal_3684) ) ;
    buf_clk new_AGEMA_reg_buffer_2332 ( .C (clk), .D (new_AGEMA_signal_3691), .Q (new_AGEMA_signal_3692) ) ;
    buf_clk new_AGEMA_reg_buffer_2340 ( .C (clk), .D (new_AGEMA_signal_3699), .Q (new_AGEMA_signal_3700) ) ;
    buf_clk new_AGEMA_reg_buffer_2348 ( .C (clk), .D (new_AGEMA_signal_3707), .Q (new_AGEMA_signal_3708) ) ;
    buf_clk new_AGEMA_reg_buffer_2356 ( .C (clk), .D (new_AGEMA_signal_3715), .Q (new_AGEMA_signal_3716) ) ;
    buf_clk new_AGEMA_reg_buffer_2364 ( .C (clk), .D (new_AGEMA_signal_3723), .Q (new_AGEMA_signal_3724) ) ;
    buf_clk new_AGEMA_reg_buffer_2372 ( .C (clk), .D (new_AGEMA_signal_3731), .Q (new_AGEMA_signal_3732) ) ;
    buf_clk new_AGEMA_reg_buffer_2380 ( .C (clk), .D (new_AGEMA_signal_3739), .Q (new_AGEMA_signal_3740) ) ;
    buf_clk new_AGEMA_reg_buffer_2388 ( .C (clk), .D (new_AGEMA_signal_3747), .Q (new_AGEMA_signal_3748) ) ;
    buf_clk new_AGEMA_reg_buffer_2396 ( .C (clk), .D (new_AGEMA_signal_3755), .Q (new_AGEMA_signal_3756) ) ;
    buf_clk new_AGEMA_reg_buffer_2404 ( .C (clk), .D (new_AGEMA_signal_3763), .Q (new_AGEMA_signal_3764) ) ;
    buf_clk new_AGEMA_reg_buffer_2412 ( .C (clk), .D (new_AGEMA_signal_3771), .Q (new_AGEMA_signal_3772) ) ;
    buf_clk new_AGEMA_reg_buffer_2420 ( .C (clk), .D (new_AGEMA_signal_3779), .Q (new_AGEMA_signal_3780) ) ;
    buf_clk new_AGEMA_reg_buffer_2428 ( .C (clk), .D (new_AGEMA_signal_3787), .Q (new_AGEMA_signal_3788) ) ;
    buf_clk new_AGEMA_reg_buffer_2436 ( .C (clk), .D (new_AGEMA_signal_3795), .Q (new_AGEMA_signal_3796) ) ;
    buf_clk new_AGEMA_reg_buffer_2444 ( .C (clk), .D (new_AGEMA_signal_3803), .Q (new_AGEMA_signal_3804) ) ;
    buf_clk new_AGEMA_reg_buffer_2452 ( .C (clk), .D (new_AGEMA_signal_3811), .Q (new_AGEMA_signal_3812) ) ;
    buf_clk new_AGEMA_reg_buffer_2460 ( .C (clk), .D (new_AGEMA_signal_3819), .Q (new_AGEMA_signal_3820) ) ;
    buf_clk new_AGEMA_reg_buffer_2468 ( .C (clk), .D (new_AGEMA_signal_3827), .Q (new_AGEMA_signal_3828) ) ;
    buf_clk new_AGEMA_reg_buffer_2476 ( .C (clk), .D (new_AGEMA_signal_3835), .Q (new_AGEMA_signal_3836) ) ;
    buf_clk new_AGEMA_reg_buffer_2484 ( .C (clk), .D (new_AGEMA_signal_3843), .Q (new_AGEMA_signal_3844) ) ;
    buf_clk new_AGEMA_reg_buffer_2492 ( .C (clk), .D (new_AGEMA_signal_3851), .Q (new_AGEMA_signal_3852) ) ;
    buf_clk new_AGEMA_reg_buffer_2500 ( .C (clk), .D (new_AGEMA_signal_3859), .Q (new_AGEMA_signal_3860) ) ;
    buf_clk new_AGEMA_reg_buffer_2508 ( .C (clk), .D (new_AGEMA_signal_3867), .Q (new_AGEMA_signal_3868) ) ;
    buf_clk new_AGEMA_reg_buffer_2516 ( .C (clk), .D (new_AGEMA_signal_3875), .Q (new_AGEMA_signal_3876) ) ;
    buf_clk new_AGEMA_reg_buffer_2524 ( .C (clk), .D (new_AGEMA_signal_3883), .Q (new_AGEMA_signal_3884) ) ;
    buf_clk new_AGEMA_reg_buffer_2532 ( .C (clk), .D (new_AGEMA_signal_3891), .Q (new_AGEMA_signal_3892) ) ;
    buf_clk new_AGEMA_reg_buffer_2540 ( .C (clk), .D (new_AGEMA_signal_3899), .Q (new_AGEMA_signal_3900) ) ;
    buf_clk new_AGEMA_reg_buffer_2548 ( .C (clk), .D (new_AGEMA_signal_3907), .Q (new_AGEMA_signal_3908) ) ;
    buf_clk new_AGEMA_reg_buffer_2556 ( .C (clk), .D (new_AGEMA_signal_3915), .Q (new_AGEMA_signal_3916) ) ;
    buf_clk new_AGEMA_reg_buffer_2564 ( .C (clk), .D (new_AGEMA_signal_3923), .Q (new_AGEMA_signal_3924) ) ;
    buf_clk new_AGEMA_reg_buffer_2572 ( .C (clk), .D (new_AGEMA_signal_3931), .Q (new_AGEMA_signal_3932) ) ;
    buf_clk new_AGEMA_reg_buffer_2580 ( .C (clk), .D (new_AGEMA_signal_3939), .Q (new_AGEMA_signal_3940) ) ;
    buf_clk new_AGEMA_reg_buffer_2588 ( .C (clk), .D (new_AGEMA_signal_3947), .Q (new_AGEMA_signal_3948) ) ;
    buf_clk new_AGEMA_reg_buffer_2596 ( .C (clk), .D (new_AGEMA_signal_3955), .Q (new_AGEMA_signal_3956) ) ;
    buf_clk new_AGEMA_reg_buffer_2604 ( .C (clk), .D (new_AGEMA_signal_3963), .Q (new_AGEMA_signal_3964) ) ;
    buf_clk new_AGEMA_reg_buffer_2612 ( .C (clk), .D (new_AGEMA_signal_3971), .Q (new_AGEMA_signal_3972) ) ;
    buf_clk new_AGEMA_reg_buffer_2620 ( .C (clk), .D (new_AGEMA_signal_3979), .Q (new_AGEMA_signal_3980) ) ;
    buf_clk new_AGEMA_reg_buffer_2628 ( .C (clk), .D (new_AGEMA_signal_3987), .Q (new_AGEMA_signal_3988) ) ;
    buf_clk new_AGEMA_reg_buffer_2636 ( .C (clk), .D (new_AGEMA_signal_3995), .Q (new_AGEMA_signal_3996) ) ;
    buf_clk new_AGEMA_reg_buffer_2644 ( .C (clk), .D (new_AGEMA_signal_4003), .Q (new_AGEMA_signal_4004) ) ;
    buf_clk new_AGEMA_reg_buffer_2652 ( .C (clk), .D (new_AGEMA_signal_4011), .Q (new_AGEMA_signal_4012) ) ;
    buf_clk new_AGEMA_reg_buffer_2660 ( .C (clk), .D (new_AGEMA_signal_4019), .Q (new_AGEMA_signal_4020) ) ;
    buf_clk new_AGEMA_reg_buffer_2668 ( .C (clk), .D (new_AGEMA_signal_4027), .Q (new_AGEMA_signal_4028) ) ;
    buf_clk new_AGEMA_reg_buffer_2676 ( .C (clk), .D (new_AGEMA_signal_4035), .Q (new_AGEMA_signal_4036) ) ;
    buf_clk new_AGEMA_reg_buffer_2684 ( .C (clk), .D (new_AGEMA_signal_4043), .Q (new_AGEMA_signal_4044) ) ;
    buf_clk new_AGEMA_reg_buffer_2692 ( .C (clk), .D (new_AGEMA_signal_4051), .Q (new_AGEMA_signal_4052) ) ;
    buf_clk new_AGEMA_reg_buffer_2700 ( .C (clk), .D (new_AGEMA_signal_4059), .Q (new_AGEMA_signal_4060) ) ;
    buf_clk new_AGEMA_reg_buffer_2708 ( .C (clk), .D (new_AGEMA_signal_4067), .Q (new_AGEMA_signal_4068) ) ;
    buf_clk new_AGEMA_reg_buffer_2716 ( .C (clk), .D (new_AGEMA_signal_4075), .Q (new_AGEMA_signal_4076) ) ;
    buf_clk new_AGEMA_reg_buffer_2724 ( .C (clk), .D (new_AGEMA_signal_4083), .Q (new_AGEMA_signal_4084) ) ;
    buf_clk new_AGEMA_reg_buffer_2732 ( .C (clk), .D (new_AGEMA_signal_4091), .Q (new_AGEMA_signal_4092) ) ;
    buf_clk new_AGEMA_reg_buffer_2740 ( .C (clk), .D (new_AGEMA_signal_4099), .Q (new_AGEMA_signal_4100) ) ;
    buf_clk new_AGEMA_reg_buffer_2748 ( .C (clk), .D (new_AGEMA_signal_4107), .Q (new_AGEMA_signal_4108) ) ;
    buf_clk new_AGEMA_reg_buffer_2756 ( .C (clk), .D (new_AGEMA_signal_4115), .Q (new_AGEMA_signal_4116) ) ;
    buf_clk new_AGEMA_reg_buffer_2764 ( .C (clk), .D (new_AGEMA_signal_4123), .Q (new_AGEMA_signal_4124) ) ;
    buf_clk new_AGEMA_reg_buffer_2772 ( .C (clk), .D (new_AGEMA_signal_4131), .Q (new_AGEMA_signal_4132) ) ;
    buf_clk new_AGEMA_reg_buffer_2780 ( .C (clk), .D (new_AGEMA_signal_4139), .Q (new_AGEMA_signal_4140) ) ;
    buf_clk new_AGEMA_reg_buffer_2788 ( .C (clk), .D (new_AGEMA_signal_4147), .Q (new_AGEMA_signal_4148) ) ;
    buf_clk new_AGEMA_reg_buffer_2796 ( .C (clk), .D (new_AGEMA_signal_4155), .Q (new_AGEMA_signal_4156) ) ;
    buf_clk new_AGEMA_reg_buffer_2804 ( .C (clk), .D (new_AGEMA_signal_4163), .Q (new_AGEMA_signal_4164) ) ;
    buf_clk new_AGEMA_reg_buffer_2812 ( .C (clk), .D (new_AGEMA_signal_4171), .Q (new_AGEMA_signal_4172) ) ;
    buf_clk new_AGEMA_reg_buffer_2820 ( .C (clk), .D (new_AGEMA_signal_4179), .Q (new_AGEMA_signal_4180) ) ;
    buf_clk new_AGEMA_reg_buffer_2828 ( .C (clk), .D (new_AGEMA_signal_4187), .Q (new_AGEMA_signal_4188) ) ;
    buf_clk new_AGEMA_reg_buffer_2836 ( .C (clk), .D (new_AGEMA_signal_4195), .Q (new_AGEMA_signal_4196) ) ;
    buf_clk new_AGEMA_reg_buffer_2844 ( .C (clk), .D (new_AGEMA_signal_4203), .Q (new_AGEMA_signal_4204) ) ;
    buf_clk new_AGEMA_reg_buffer_2852 ( .C (clk), .D (new_AGEMA_signal_4211), .Q (new_AGEMA_signal_4212) ) ;
    buf_clk new_AGEMA_reg_buffer_2860 ( .C (clk), .D (new_AGEMA_signal_4219), .Q (new_AGEMA_signal_4220) ) ;
    buf_clk new_AGEMA_reg_buffer_2868 ( .C (clk), .D (new_AGEMA_signal_4227), .Q (new_AGEMA_signal_4228) ) ;
    buf_clk new_AGEMA_reg_buffer_2876 ( .C (clk), .D (new_AGEMA_signal_4235), .Q (new_AGEMA_signal_4236) ) ;
    buf_clk new_AGEMA_reg_buffer_2884 ( .C (clk), .D (new_AGEMA_signal_4243), .Q (new_AGEMA_signal_4244) ) ;
    buf_clk new_AGEMA_reg_buffer_2892 ( .C (clk), .D (new_AGEMA_signal_4251), .Q (new_AGEMA_signal_4252) ) ;
    buf_clk new_AGEMA_reg_buffer_2900 ( .C (clk), .D (new_AGEMA_signal_4259), .Q (new_AGEMA_signal_4260) ) ;
    buf_clk new_AGEMA_reg_buffer_2908 ( .C (clk), .D (new_AGEMA_signal_4267), .Q (new_AGEMA_signal_4268) ) ;
    buf_clk new_AGEMA_reg_buffer_2916 ( .C (clk), .D (new_AGEMA_signal_4275), .Q (new_AGEMA_signal_4276) ) ;
    buf_clk new_AGEMA_reg_buffer_2924 ( .C (clk), .D (new_AGEMA_signal_4283), .Q (new_AGEMA_signal_4284) ) ;
    buf_clk new_AGEMA_reg_buffer_2932 ( .C (clk), .D (new_AGEMA_signal_4291), .Q (new_AGEMA_signal_4292) ) ;
    buf_clk new_AGEMA_reg_buffer_2940 ( .C (clk), .D (new_AGEMA_signal_4299), .Q (new_AGEMA_signal_4300) ) ;
    buf_clk new_AGEMA_reg_buffer_2948 ( .C (clk), .D (new_AGEMA_signal_4307), .Q (new_AGEMA_signal_4308) ) ;
    buf_clk new_AGEMA_reg_buffer_2956 ( .C (clk), .D (new_AGEMA_signal_4315), .Q (new_AGEMA_signal_4316) ) ;
    buf_clk new_AGEMA_reg_buffer_2964 ( .C (clk), .D (new_AGEMA_signal_4323), .Q (new_AGEMA_signal_4324) ) ;
    buf_clk new_AGEMA_reg_buffer_2972 ( .C (clk), .D (new_AGEMA_signal_4331), .Q (new_AGEMA_signal_4332) ) ;
    buf_clk new_AGEMA_reg_buffer_2980 ( .C (clk), .D (new_AGEMA_signal_4339), .Q (new_AGEMA_signal_4340) ) ;
    buf_clk new_AGEMA_reg_buffer_2988 ( .C (clk), .D (new_AGEMA_signal_4347), .Q (new_AGEMA_signal_4348) ) ;
    buf_clk new_AGEMA_reg_buffer_2996 ( .C (clk), .D (new_AGEMA_signal_4355), .Q (new_AGEMA_signal_4356) ) ;
    buf_clk new_AGEMA_reg_buffer_3004 ( .C (clk), .D (new_AGEMA_signal_4363), .Q (new_AGEMA_signal_4364) ) ;
    buf_clk new_AGEMA_reg_buffer_3012 ( .C (clk), .D (new_AGEMA_signal_4371), .Q (new_AGEMA_signal_4372) ) ;
    buf_clk new_AGEMA_reg_buffer_3020 ( .C (clk), .D (new_AGEMA_signal_4379), .Q (new_AGEMA_signal_4380) ) ;
    buf_clk new_AGEMA_reg_buffer_3028 ( .C (clk), .D (new_AGEMA_signal_4387), .Q (new_AGEMA_signal_4388) ) ;
    buf_clk new_AGEMA_reg_buffer_3036 ( .C (clk), .D (new_AGEMA_signal_4395), .Q (new_AGEMA_signal_4396) ) ;
    buf_clk new_AGEMA_reg_buffer_3044 ( .C (clk), .D (new_AGEMA_signal_4403), .Q (new_AGEMA_signal_4404) ) ;
    buf_clk new_AGEMA_reg_buffer_3052 ( .C (clk), .D (new_AGEMA_signal_4411), .Q (new_AGEMA_signal_4412) ) ;
    buf_clk new_AGEMA_reg_buffer_3060 ( .C (clk), .D (new_AGEMA_signal_4419), .Q (new_AGEMA_signal_4420) ) ;
    buf_clk new_AGEMA_reg_buffer_3388 ( .C (clk), .D (new_AGEMA_signal_4747), .Q (new_AGEMA_signal_4748) ) ;
    buf_clk new_AGEMA_reg_buffer_3396 ( .C (clk), .D (new_AGEMA_signal_4755), .Q (new_AGEMA_signal_4756) ) ;
    buf_clk new_AGEMA_reg_buffer_3404 ( .C (clk), .D (new_AGEMA_signal_4763), .Q (new_AGEMA_signal_4764) ) ;
    buf_clk new_AGEMA_reg_buffer_3412 ( .C (clk), .D (new_AGEMA_signal_4771), .Q (new_AGEMA_signal_4772) ) ;
    buf_clk new_AGEMA_reg_buffer_3420 ( .C (clk), .D (new_AGEMA_signal_4779), .Q (new_AGEMA_signal_4780) ) ;
    buf_clk new_AGEMA_reg_buffer_3428 ( .C (clk), .D (new_AGEMA_signal_4787), .Q (new_AGEMA_signal_4788) ) ;
    buf_clk new_AGEMA_reg_buffer_3436 ( .C (clk), .D (new_AGEMA_signal_4795), .Q (new_AGEMA_signal_4796) ) ;
    buf_clk new_AGEMA_reg_buffer_3444 ( .C (clk), .D (new_AGEMA_signal_4803), .Q (new_AGEMA_signal_4804) ) ;
    buf_clk new_AGEMA_reg_buffer_3452 ( .C (clk), .D (new_AGEMA_signal_4811), .Q (new_AGEMA_signal_4812) ) ;
    buf_clk new_AGEMA_reg_buffer_3460 ( .C (clk), .D (new_AGEMA_signal_4819), .Q (new_AGEMA_signal_4820) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_1077 ( .C (clk), .D (new_AGEMA_signal_2436), .Q (new_AGEMA_signal_2437) ) ;
    buf_clk new_AGEMA_reg_buffer_1083 ( .C (clk), .D (new_AGEMA_signal_2442), .Q (new_AGEMA_signal_2443) ) ;
    buf_clk new_AGEMA_reg_buffer_1089 ( .C (clk), .D (new_AGEMA_signal_2448), .Q (new_AGEMA_signal_2449) ) ;
    buf_clk new_AGEMA_reg_buffer_1095 ( .C (clk), .D (new_AGEMA_signal_2454), .Q (new_AGEMA_signal_2455) ) ;
    buf_clk new_AGEMA_reg_buffer_1101 ( .C (clk), .D (new_AGEMA_signal_2460), .Q (new_AGEMA_signal_2461) ) ;
    buf_clk new_AGEMA_reg_buffer_1107 ( .C (clk), .D (new_AGEMA_signal_2466), .Q (new_AGEMA_signal_2467) ) ;
    buf_clk new_AGEMA_reg_buffer_1113 ( .C (clk), .D (new_AGEMA_signal_2472), .Q (new_AGEMA_signal_2473) ) ;
    buf_clk new_AGEMA_reg_buffer_1119 ( .C (clk), .D (new_AGEMA_signal_2478), .Q (new_AGEMA_signal_2479) ) ;
    buf_clk new_AGEMA_reg_buffer_1125 ( .C (clk), .D (new_AGEMA_signal_2484), .Q (new_AGEMA_signal_2485) ) ;
    buf_clk new_AGEMA_reg_buffer_1131 ( .C (clk), .D (new_AGEMA_signal_2490), .Q (new_AGEMA_signal_2491) ) ;
    buf_clk new_AGEMA_reg_buffer_1137 ( .C (clk), .D (new_AGEMA_signal_2496), .Q (new_AGEMA_signal_2497) ) ;
    buf_clk new_AGEMA_reg_buffer_1143 ( .C (clk), .D (new_AGEMA_signal_2502), .Q (new_AGEMA_signal_2503) ) ;
    buf_clk new_AGEMA_reg_buffer_1149 ( .C (clk), .D (new_AGEMA_signal_2508), .Q (new_AGEMA_signal_2509) ) ;
    buf_clk new_AGEMA_reg_buffer_1155 ( .C (clk), .D (new_AGEMA_signal_2514), .Q (new_AGEMA_signal_2515) ) ;
    buf_clk new_AGEMA_reg_buffer_1161 ( .C (clk), .D (new_AGEMA_signal_2520), .Q (new_AGEMA_signal_2521) ) ;
    buf_clk new_AGEMA_reg_buffer_1167 ( .C (clk), .D (new_AGEMA_signal_2526), .Q (new_AGEMA_signal_2527) ) ;
    buf_clk new_AGEMA_reg_buffer_1173 ( .C (clk), .D (new_AGEMA_signal_2532), .Q (new_AGEMA_signal_2533) ) ;
    buf_clk new_AGEMA_reg_buffer_1179 ( .C (clk), .D (new_AGEMA_signal_2538), .Q (new_AGEMA_signal_2539) ) ;
    buf_clk new_AGEMA_reg_buffer_1185 ( .C (clk), .D (new_AGEMA_signal_2544), .Q (new_AGEMA_signal_2545) ) ;
    buf_clk new_AGEMA_reg_buffer_1191 ( .C (clk), .D (new_AGEMA_signal_2550), .Q (new_AGEMA_signal_2551) ) ;
    buf_clk new_AGEMA_reg_buffer_1197 ( .C (clk), .D (new_AGEMA_signal_2556), .Q (new_AGEMA_signal_2557) ) ;
    buf_clk new_AGEMA_reg_buffer_1203 ( .C (clk), .D (new_AGEMA_signal_2562), .Q (new_AGEMA_signal_2563) ) ;
    buf_clk new_AGEMA_reg_buffer_1209 ( .C (clk), .D (new_AGEMA_signal_2568), .Q (new_AGEMA_signal_2569) ) ;
    buf_clk new_AGEMA_reg_buffer_1215 ( .C (clk), .D (new_AGEMA_signal_2574), .Q (new_AGEMA_signal_2575) ) ;
    buf_clk new_AGEMA_reg_buffer_1221 ( .C (clk), .D (new_AGEMA_signal_2580), .Q (new_AGEMA_signal_2581) ) ;
    buf_clk new_AGEMA_reg_buffer_1227 ( .C (clk), .D (new_AGEMA_signal_2586), .Q (new_AGEMA_signal_2587) ) ;
    buf_clk new_AGEMA_reg_buffer_1233 ( .C (clk), .D (new_AGEMA_signal_2592), .Q (new_AGEMA_signal_2593) ) ;
    buf_clk new_AGEMA_reg_buffer_1239 ( .C (clk), .D (new_AGEMA_signal_2598), .Q (new_AGEMA_signal_2599) ) ;
    buf_clk new_AGEMA_reg_buffer_1245 ( .C (clk), .D (new_AGEMA_signal_2604), .Q (new_AGEMA_signal_2605) ) ;
    buf_clk new_AGEMA_reg_buffer_1251 ( .C (clk), .D (new_AGEMA_signal_2610), .Q (new_AGEMA_signal_2611) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C (clk), .D (new_AGEMA_signal_2616), .Q (new_AGEMA_signal_2617) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C (clk), .D (new_AGEMA_signal_2622), .Q (new_AGEMA_signal_2623) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C (clk), .D (new_AGEMA_signal_2628), .Q (new_AGEMA_signal_2629) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C (clk), .D (new_AGEMA_signal_2634), .Q (new_AGEMA_signal_2635) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C (clk), .D (new_AGEMA_signal_2640), .Q (new_AGEMA_signal_2641) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C (clk), .D (new_AGEMA_signal_2646), .Q (new_AGEMA_signal_2647) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C (clk), .D (new_AGEMA_signal_2652), .Q (new_AGEMA_signal_2653) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C (clk), .D (new_AGEMA_signal_2658), .Q (new_AGEMA_signal_2659) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C (clk), .D (new_AGEMA_signal_2664), .Q (new_AGEMA_signal_2665) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C (clk), .D (new_AGEMA_signal_2670), .Q (new_AGEMA_signal_2671) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C (clk), .D (new_AGEMA_signal_2676), .Q (new_AGEMA_signal_2677) ) ;
    buf_clk new_AGEMA_reg_buffer_1323 ( .C (clk), .D (new_AGEMA_signal_2682), .Q (new_AGEMA_signal_2683) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C (clk), .D (new_AGEMA_signal_2688), .Q (new_AGEMA_signal_2689) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C (clk), .D (new_AGEMA_signal_2694), .Q (new_AGEMA_signal_2695) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C (clk), .D (new_AGEMA_signal_2700), .Q (new_AGEMA_signal_2701) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C (clk), .D (new_AGEMA_signal_2706), .Q (new_AGEMA_signal_2707) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C (clk), .D (new_AGEMA_signal_2712), .Q (new_AGEMA_signal_2713) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C (clk), .D (new_AGEMA_signal_2718), .Q (new_AGEMA_signal_2719) ) ;
    buf_clk new_AGEMA_reg_buffer_1365 ( .C (clk), .D (new_AGEMA_signal_2724), .Q (new_AGEMA_signal_2725) ) ;
    buf_clk new_AGEMA_reg_buffer_1371 ( .C (clk), .D (new_AGEMA_signal_2730), .Q (new_AGEMA_signal_2731) ) ;
    buf_clk new_AGEMA_reg_buffer_1377 ( .C (clk), .D (new_AGEMA_signal_2736), .Q (new_AGEMA_signal_2737) ) ;
    buf_clk new_AGEMA_reg_buffer_1383 ( .C (clk), .D (new_AGEMA_signal_2742), .Q (new_AGEMA_signal_2743) ) ;
    buf_clk new_AGEMA_reg_buffer_1389 ( .C (clk), .D (new_AGEMA_signal_2748), .Q (new_AGEMA_signal_2749) ) ;
    buf_clk new_AGEMA_reg_buffer_1395 ( .C (clk), .D (new_AGEMA_signal_2754), .Q (new_AGEMA_signal_2755) ) ;
    buf_clk new_AGEMA_reg_buffer_1401 ( .C (clk), .D (new_AGEMA_signal_2760), .Q (new_AGEMA_signal_2761) ) ;
    buf_clk new_AGEMA_reg_buffer_1407 ( .C (clk), .D (new_AGEMA_signal_2766), .Q (new_AGEMA_signal_2767) ) ;
    buf_clk new_AGEMA_reg_buffer_1413 ( .C (clk), .D (new_AGEMA_signal_2772), .Q (new_AGEMA_signal_2773) ) ;
    buf_clk new_AGEMA_reg_buffer_1419 ( .C (clk), .D (new_AGEMA_signal_2778), .Q (new_AGEMA_signal_2779) ) ;
    buf_clk new_AGEMA_reg_buffer_1425 ( .C (clk), .D (new_AGEMA_signal_2784), .Q (new_AGEMA_signal_2785) ) ;
    buf_clk new_AGEMA_reg_buffer_1431 ( .C (clk), .D (new_AGEMA_signal_2790), .Q (new_AGEMA_signal_2791) ) ;
    buf_clk new_AGEMA_reg_buffer_1437 ( .C (clk), .D (new_AGEMA_signal_2796), .Q (new_AGEMA_signal_2797) ) ;
    buf_clk new_AGEMA_reg_buffer_1443 ( .C (clk), .D (new_AGEMA_signal_2802), .Q (new_AGEMA_signal_2803) ) ;
    buf_clk new_AGEMA_reg_buffer_1449 ( .C (clk), .D (new_AGEMA_signal_2808), .Q (new_AGEMA_signal_2809) ) ;
    buf_clk new_AGEMA_reg_buffer_1455 ( .C (clk), .D (new_AGEMA_signal_2814), .Q (new_AGEMA_signal_2815) ) ;
    buf_clk new_AGEMA_reg_buffer_1461 ( .C (clk), .D (new_AGEMA_signal_2820), .Q (new_AGEMA_signal_2821) ) ;
    buf_clk new_AGEMA_reg_buffer_1467 ( .C (clk), .D (new_AGEMA_signal_2826), .Q (new_AGEMA_signal_2827) ) ;
    buf_clk new_AGEMA_reg_buffer_1473 ( .C (clk), .D (new_AGEMA_signal_2832), .Q (new_AGEMA_signal_2833) ) ;
    buf_clk new_AGEMA_reg_buffer_1479 ( .C (clk), .D (new_AGEMA_signal_2838), .Q (new_AGEMA_signal_2839) ) ;
    buf_clk new_AGEMA_reg_buffer_1485 ( .C (clk), .D (new_AGEMA_signal_2844), .Q (new_AGEMA_signal_2845) ) ;
    buf_clk new_AGEMA_reg_buffer_1491 ( .C (clk), .D (new_AGEMA_signal_2850), .Q (new_AGEMA_signal_2851) ) ;
    buf_clk new_AGEMA_reg_buffer_1497 ( .C (clk), .D (new_AGEMA_signal_2856), .Q (new_AGEMA_signal_2857) ) ;
    buf_clk new_AGEMA_reg_buffer_1503 ( .C (clk), .D (new_AGEMA_signal_2862), .Q (new_AGEMA_signal_2863) ) ;
    buf_clk new_AGEMA_reg_buffer_1509 ( .C (clk), .D (new_AGEMA_signal_2868), .Q (new_AGEMA_signal_2869) ) ;
    buf_clk new_AGEMA_reg_buffer_1515 ( .C (clk), .D (new_AGEMA_signal_2874), .Q (new_AGEMA_signal_2875) ) ;
    buf_clk new_AGEMA_reg_buffer_1521 ( .C (clk), .D (new_AGEMA_signal_2880), .Q (new_AGEMA_signal_2881) ) ;
    buf_clk new_AGEMA_reg_buffer_1527 ( .C (clk), .D (new_AGEMA_signal_2886), .Q (new_AGEMA_signal_2887) ) ;
    buf_clk new_AGEMA_reg_buffer_1533 ( .C (clk), .D (new_AGEMA_signal_2892), .Q (new_AGEMA_signal_2893) ) ;
    buf_clk new_AGEMA_reg_buffer_1539 ( .C (clk), .D (new_AGEMA_signal_2898), .Q (new_AGEMA_signal_2899) ) ;
    buf_clk new_AGEMA_reg_buffer_1545 ( .C (clk), .D (new_AGEMA_signal_2904), .Q (new_AGEMA_signal_2905) ) ;
    buf_clk new_AGEMA_reg_buffer_1551 ( .C (clk), .D (new_AGEMA_signal_2910), .Q (new_AGEMA_signal_2911) ) ;
    buf_clk new_AGEMA_reg_buffer_1557 ( .C (clk), .D (new_AGEMA_signal_2916), .Q (new_AGEMA_signal_2917) ) ;
    buf_clk new_AGEMA_reg_buffer_1563 ( .C (clk), .D (new_AGEMA_signal_2922), .Q (new_AGEMA_signal_2923) ) ;
    buf_clk new_AGEMA_reg_buffer_1569 ( .C (clk), .D (new_AGEMA_signal_2928), .Q (new_AGEMA_signal_2929) ) ;
    buf_clk new_AGEMA_reg_buffer_1575 ( .C (clk), .D (new_AGEMA_signal_2934), .Q (new_AGEMA_signal_2935) ) ;
    buf_clk new_AGEMA_reg_buffer_1581 ( .C (clk), .D (new_AGEMA_signal_2940), .Q (new_AGEMA_signal_2941) ) ;
    buf_clk new_AGEMA_reg_buffer_1587 ( .C (clk), .D (new_AGEMA_signal_2946), .Q (new_AGEMA_signal_2947) ) ;
    buf_clk new_AGEMA_reg_buffer_1593 ( .C (clk), .D (new_AGEMA_signal_2952), .Q (new_AGEMA_signal_2953) ) ;
    buf_clk new_AGEMA_reg_buffer_1599 ( .C (clk), .D (new_AGEMA_signal_2958), .Q (new_AGEMA_signal_2959) ) ;
    buf_clk new_AGEMA_reg_buffer_1605 ( .C (clk), .D (new_AGEMA_signal_2964), .Q (new_AGEMA_signal_2965) ) ;
    buf_clk new_AGEMA_reg_buffer_1611 ( .C (clk), .D (new_AGEMA_signal_2970), .Q (new_AGEMA_signal_2971) ) ;
    buf_clk new_AGEMA_reg_buffer_1617 ( .C (clk), .D (new_AGEMA_signal_2976), .Q (new_AGEMA_signal_2977) ) ;
    buf_clk new_AGEMA_reg_buffer_1623 ( .C (clk), .D (new_AGEMA_signal_2982), .Q (new_AGEMA_signal_2983) ) ;
    buf_clk new_AGEMA_reg_buffer_1629 ( .C (clk), .D (new_AGEMA_signal_2988), .Q (new_AGEMA_signal_2989) ) ;
    buf_clk new_AGEMA_reg_buffer_1635 ( .C (clk), .D (new_AGEMA_signal_2994), .Q (new_AGEMA_signal_2995) ) ;
    buf_clk new_AGEMA_reg_buffer_1641 ( .C (clk), .D (new_AGEMA_signal_3000), .Q (new_AGEMA_signal_3001) ) ;
    buf_clk new_AGEMA_reg_buffer_1647 ( .C (clk), .D (new_AGEMA_signal_3006), .Q (new_AGEMA_signal_3007) ) ;
    buf_clk new_AGEMA_reg_buffer_1653 ( .C (clk), .D (new_AGEMA_signal_3012), .Q (new_AGEMA_signal_3013) ) ;
    buf_clk new_AGEMA_reg_buffer_1659 ( .C (clk), .D (new_AGEMA_signal_3018), .Q (new_AGEMA_signal_3019) ) ;
    buf_clk new_AGEMA_reg_buffer_1665 ( .C (clk), .D (new_AGEMA_signal_3024), .Q (new_AGEMA_signal_3025) ) ;
    buf_clk new_AGEMA_reg_buffer_1671 ( .C (clk), .D (new_AGEMA_signal_3030), .Q (new_AGEMA_signal_3031) ) ;
    buf_clk new_AGEMA_reg_buffer_1677 ( .C (clk), .D (new_AGEMA_signal_3036), .Q (new_AGEMA_signal_3037) ) ;
    buf_clk new_AGEMA_reg_buffer_1683 ( .C (clk), .D (new_AGEMA_signal_3042), .Q (new_AGEMA_signal_3043) ) ;
    buf_clk new_AGEMA_reg_buffer_1689 ( .C (clk), .D (new_AGEMA_signal_3048), .Q (new_AGEMA_signal_3049) ) ;
    buf_clk new_AGEMA_reg_buffer_1695 ( .C (clk), .D (new_AGEMA_signal_3054), .Q (new_AGEMA_signal_3055) ) ;
    buf_clk new_AGEMA_reg_buffer_1701 ( .C (clk), .D (new_AGEMA_signal_3060), .Q (new_AGEMA_signal_3061) ) ;
    buf_clk new_AGEMA_reg_buffer_1707 ( .C (clk), .D (new_AGEMA_signal_3066), .Q (new_AGEMA_signal_3067) ) ;
    buf_clk new_AGEMA_reg_buffer_1713 ( .C (clk), .D (new_AGEMA_signal_3072), .Q (new_AGEMA_signal_3073) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C (clk), .D (new_AGEMA_signal_3078), .Q (new_AGEMA_signal_3079) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C (clk), .D (new_AGEMA_signal_3084), .Q (new_AGEMA_signal_3085) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C (clk), .D (new_AGEMA_signal_3090), .Q (new_AGEMA_signal_3091) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C (clk), .D (new_AGEMA_signal_3096), .Q (new_AGEMA_signal_3097) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C (clk), .D (new_AGEMA_signal_3102), .Q (new_AGEMA_signal_3103) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C (clk), .D (new_AGEMA_signal_3108), .Q (new_AGEMA_signal_3109) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C (clk), .D (new_AGEMA_signal_3114), .Q (new_AGEMA_signal_3115) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C (clk), .D (new_AGEMA_signal_3120), .Q (new_AGEMA_signal_3121) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C (clk), .D (new_AGEMA_signal_3126), .Q (new_AGEMA_signal_3127) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C (clk), .D (new_AGEMA_signal_3132), .Q (new_AGEMA_signal_3133) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C (clk), .D (new_AGEMA_signal_3138), .Q (new_AGEMA_signal_3139) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C (clk), .D (new_AGEMA_signal_3144), .Q (new_AGEMA_signal_3145) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C (clk), .D (new_AGEMA_signal_3150), .Q (new_AGEMA_signal_3151) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C (clk), .D (new_AGEMA_signal_3156), .Q (new_AGEMA_signal_3157) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C (clk), .D (new_AGEMA_signal_3162), .Q (new_AGEMA_signal_3163) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C (clk), .D (new_AGEMA_signal_3168), .Q (new_AGEMA_signal_3169) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C (clk), .D (new_AGEMA_signal_3174), .Q (new_AGEMA_signal_3175) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C (clk), .D (new_AGEMA_signal_3180), .Q (new_AGEMA_signal_3181) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C (clk), .D (new_AGEMA_signal_3186), .Q (new_AGEMA_signal_3187) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C (clk), .D (new_AGEMA_signal_3192), .Q (new_AGEMA_signal_3193) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C (clk), .D (new_AGEMA_signal_3198), .Q (new_AGEMA_signal_3199) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C (clk), .D (new_AGEMA_signal_3204), .Q (new_AGEMA_signal_3205) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C (clk), .D (SubCellInst_SboxInst_0_n15), .Q (new_AGEMA_signal_3209) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C (clk), .D (new_AGEMA_signal_1148), .Q (new_AGEMA_signal_3211) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C (clk), .D (new_AGEMA_signal_2180), .Q (new_AGEMA_signal_3213) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C (clk), .D (new_AGEMA_signal_2182), .Q (new_AGEMA_signal_3215) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C (clk), .D (SubCellInst_SboxInst_0_n6), .Q (new_AGEMA_signal_3217) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C (clk), .D (new_AGEMA_signal_1150), .Q (new_AGEMA_signal_3219) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C (clk), .D (SubCellInst_SboxInst_1_n15), .Q (new_AGEMA_signal_3221) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C (clk), .D (new_AGEMA_signal_1154), .Q (new_AGEMA_signal_3223) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C (clk), .D (new_AGEMA_signal_2196), .Q (new_AGEMA_signal_3225) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C (clk), .D (new_AGEMA_signal_2198), .Q (new_AGEMA_signal_3227) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C (clk), .D (SubCellInst_SboxInst_1_n6), .Q (new_AGEMA_signal_3229) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C (clk), .D (new_AGEMA_signal_1156), .Q (new_AGEMA_signal_3231) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C (clk), .D (SubCellInst_SboxInst_2_n15), .Q (new_AGEMA_signal_3233) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C (clk), .D (new_AGEMA_signal_1160), .Q (new_AGEMA_signal_3235) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C (clk), .D (new_AGEMA_signal_2212), .Q (new_AGEMA_signal_3237) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C (clk), .D (new_AGEMA_signal_2214), .Q (new_AGEMA_signal_3239) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C (clk), .D (SubCellInst_SboxInst_2_n6), .Q (new_AGEMA_signal_3241) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C (clk), .D (new_AGEMA_signal_1162), .Q (new_AGEMA_signal_3243) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C (clk), .D (SubCellInst_SboxInst_3_n15), .Q (new_AGEMA_signal_3245) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C (clk), .D (new_AGEMA_signal_1166), .Q (new_AGEMA_signal_3247) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C (clk), .D (new_AGEMA_signal_2228), .Q (new_AGEMA_signal_3249) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C (clk), .D (new_AGEMA_signal_2230), .Q (new_AGEMA_signal_3251) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C (clk), .D (SubCellInst_SboxInst_3_n6), .Q (new_AGEMA_signal_3253) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C (clk), .D (new_AGEMA_signal_1168), .Q (new_AGEMA_signal_3255) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C (clk), .D (SubCellInst_SboxInst_4_n15), .Q (new_AGEMA_signal_3257) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C (clk), .D (new_AGEMA_signal_1172), .Q (new_AGEMA_signal_3259) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C (clk), .D (new_AGEMA_signal_2244), .Q (new_AGEMA_signal_3261) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C (clk), .D (new_AGEMA_signal_2246), .Q (new_AGEMA_signal_3263) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C (clk), .D (SubCellInst_SboxInst_4_n6), .Q (new_AGEMA_signal_3265) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C (clk), .D (new_AGEMA_signal_1174), .Q (new_AGEMA_signal_3267) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C (clk), .D (SubCellInst_SboxInst_5_n15), .Q (new_AGEMA_signal_3269) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C (clk), .D (new_AGEMA_signal_1178), .Q (new_AGEMA_signal_3271) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C (clk), .D (new_AGEMA_signal_2260), .Q (new_AGEMA_signal_3273) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C (clk), .D (new_AGEMA_signal_2262), .Q (new_AGEMA_signal_3275) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C (clk), .D (SubCellInst_SboxInst_5_n6), .Q (new_AGEMA_signal_3277) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C (clk), .D (new_AGEMA_signal_1180), .Q (new_AGEMA_signal_3279) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C (clk), .D (SubCellInst_SboxInst_6_n15), .Q (new_AGEMA_signal_3281) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C (clk), .D (new_AGEMA_signal_1184), .Q (new_AGEMA_signal_3283) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C (clk), .D (new_AGEMA_signal_2276), .Q (new_AGEMA_signal_3285) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C (clk), .D (new_AGEMA_signal_2278), .Q (new_AGEMA_signal_3287) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C (clk), .D (SubCellInst_SboxInst_6_n6), .Q (new_AGEMA_signal_3289) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C (clk), .D (new_AGEMA_signal_1186), .Q (new_AGEMA_signal_3291) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C (clk), .D (SubCellInst_SboxInst_7_n15), .Q (new_AGEMA_signal_3293) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C (clk), .D (new_AGEMA_signal_1190), .Q (new_AGEMA_signal_3295) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C (clk), .D (new_AGEMA_signal_2292), .Q (new_AGEMA_signal_3297) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C (clk), .D (new_AGEMA_signal_2294), .Q (new_AGEMA_signal_3299) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C (clk), .D (SubCellInst_SboxInst_7_n6), .Q (new_AGEMA_signal_3301) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C (clk), .D (new_AGEMA_signal_1192), .Q (new_AGEMA_signal_3303) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C (clk), .D (SubCellInst_SboxInst_8_n15), .Q (new_AGEMA_signal_3305) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C (clk), .D (new_AGEMA_signal_1196), .Q (new_AGEMA_signal_3307) ) ;
    buf_clk new_AGEMA_reg_buffer_1949 ( .C (clk), .D (new_AGEMA_signal_2308), .Q (new_AGEMA_signal_3309) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C (clk), .D (new_AGEMA_signal_2310), .Q (new_AGEMA_signal_3311) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C (clk), .D (SubCellInst_SboxInst_8_n6), .Q (new_AGEMA_signal_3313) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C (clk), .D (new_AGEMA_signal_1198), .Q (new_AGEMA_signal_3315) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C (clk), .D (SubCellInst_SboxInst_9_n15), .Q (new_AGEMA_signal_3317) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C (clk), .D (new_AGEMA_signal_1202), .Q (new_AGEMA_signal_3319) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C (clk), .D (new_AGEMA_signal_2324), .Q (new_AGEMA_signal_3321) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C (clk), .D (new_AGEMA_signal_2326), .Q (new_AGEMA_signal_3323) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C (clk), .D (SubCellInst_SboxInst_9_n6), .Q (new_AGEMA_signal_3325) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C (clk), .D (new_AGEMA_signal_1204), .Q (new_AGEMA_signal_3327) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C (clk), .D (SubCellInst_SboxInst_10_n15), .Q (new_AGEMA_signal_3329) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C (clk), .D (new_AGEMA_signal_1208), .Q (new_AGEMA_signal_3331) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C (clk), .D (new_AGEMA_signal_2340), .Q (new_AGEMA_signal_3333) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C (clk), .D (new_AGEMA_signal_2342), .Q (new_AGEMA_signal_3335) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C (clk), .D (SubCellInst_SboxInst_10_n6), .Q (new_AGEMA_signal_3337) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C (clk), .D (new_AGEMA_signal_1210), .Q (new_AGEMA_signal_3339) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C (clk), .D (SubCellInst_SboxInst_11_n15), .Q (new_AGEMA_signal_3341) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C (clk), .D (new_AGEMA_signal_1214), .Q (new_AGEMA_signal_3343) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C (clk), .D (new_AGEMA_signal_2356), .Q (new_AGEMA_signal_3345) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C (clk), .D (new_AGEMA_signal_2358), .Q (new_AGEMA_signal_3347) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C (clk), .D (SubCellInst_SboxInst_11_n6), .Q (new_AGEMA_signal_3349) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C (clk), .D (new_AGEMA_signal_1216), .Q (new_AGEMA_signal_3351) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C (clk), .D (SubCellInst_SboxInst_12_n15), .Q (new_AGEMA_signal_3353) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C (clk), .D (new_AGEMA_signal_1220), .Q (new_AGEMA_signal_3355) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C (clk), .D (new_AGEMA_signal_2372), .Q (new_AGEMA_signal_3357) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C (clk), .D (new_AGEMA_signal_2374), .Q (new_AGEMA_signal_3359) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C (clk), .D (SubCellInst_SboxInst_12_n6), .Q (new_AGEMA_signal_3361) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C (clk), .D (new_AGEMA_signal_1222), .Q (new_AGEMA_signal_3363) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C (clk), .D (SubCellInst_SboxInst_13_n15), .Q (new_AGEMA_signal_3365) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C (clk), .D (new_AGEMA_signal_1226), .Q (new_AGEMA_signal_3367) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C (clk), .D (new_AGEMA_signal_2388), .Q (new_AGEMA_signal_3369) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C (clk), .D (new_AGEMA_signal_2390), .Q (new_AGEMA_signal_3371) ) ;
    buf_clk new_AGEMA_reg_buffer_2013 ( .C (clk), .D (SubCellInst_SboxInst_13_n6), .Q (new_AGEMA_signal_3373) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C (clk), .D (new_AGEMA_signal_1228), .Q (new_AGEMA_signal_3375) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C (clk), .D (SubCellInst_SboxInst_14_n15), .Q (new_AGEMA_signal_3377) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C (clk), .D (new_AGEMA_signal_1232), .Q (new_AGEMA_signal_3379) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C (clk), .D (new_AGEMA_signal_2404), .Q (new_AGEMA_signal_3381) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C (clk), .D (new_AGEMA_signal_2406), .Q (new_AGEMA_signal_3383) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C (clk), .D (SubCellInst_SboxInst_14_n6), .Q (new_AGEMA_signal_3385) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C (clk), .D (new_AGEMA_signal_1234), .Q (new_AGEMA_signal_3387) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C (clk), .D (SubCellInst_SboxInst_15_n15), .Q (new_AGEMA_signal_3389) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C (clk), .D (new_AGEMA_signal_1238), .Q (new_AGEMA_signal_3391) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C (clk), .D (new_AGEMA_signal_2420), .Q (new_AGEMA_signal_3393) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C (clk), .D (new_AGEMA_signal_2422), .Q (new_AGEMA_signal_3395) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C (clk), .D (SubCellInst_SboxInst_15_n6), .Q (new_AGEMA_signal_3397) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C (clk), .D (new_AGEMA_signal_1240), .Q (new_AGEMA_signal_3399) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C (clk), .D (new_AGEMA_signal_3404), .Q (new_AGEMA_signal_3405) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C (clk), .D (new_AGEMA_signal_3412), .Q (new_AGEMA_signal_3413) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C (clk), .D (new_AGEMA_signal_3420), .Q (new_AGEMA_signal_3421) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C (clk), .D (new_AGEMA_signal_3428), .Q (new_AGEMA_signal_3429) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C (clk), .D (new_AGEMA_signal_3436), .Q (new_AGEMA_signal_3437) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C (clk), .D (new_AGEMA_signal_3444), .Q (new_AGEMA_signal_3445) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C (clk), .D (new_AGEMA_signal_3452), .Q (new_AGEMA_signal_3453) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C (clk), .D (new_AGEMA_signal_3460), .Q (new_AGEMA_signal_3461) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C (clk), .D (new_AGEMA_signal_3468), .Q (new_AGEMA_signal_3469) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C (clk), .D (new_AGEMA_signal_3476), .Q (new_AGEMA_signal_3477) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C (clk), .D (new_AGEMA_signal_3484), .Q (new_AGEMA_signal_3485) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C (clk), .D (new_AGEMA_signal_3492), .Q (new_AGEMA_signal_3493) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C (clk), .D (new_AGEMA_signal_3500), .Q (new_AGEMA_signal_3501) ) ;
    buf_clk new_AGEMA_reg_buffer_2149 ( .C (clk), .D (new_AGEMA_signal_3508), .Q (new_AGEMA_signal_3509) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C (clk), .D (new_AGEMA_signal_3516), .Q (new_AGEMA_signal_3517) ) ;
    buf_clk new_AGEMA_reg_buffer_2165 ( .C (clk), .D (new_AGEMA_signal_3524), .Q (new_AGEMA_signal_3525) ) ;
    buf_clk new_AGEMA_reg_buffer_2173 ( .C (clk), .D (new_AGEMA_signal_3532), .Q (new_AGEMA_signal_3533) ) ;
    buf_clk new_AGEMA_reg_buffer_2181 ( .C (clk), .D (new_AGEMA_signal_3540), .Q (new_AGEMA_signal_3541) ) ;
    buf_clk new_AGEMA_reg_buffer_2189 ( .C (clk), .D (new_AGEMA_signal_3548), .Q (new_AGEMA_signal_3549) ) ;
    buf_clk new_AGEMA_reg_buffer_2197 ( .C (clk), .D (new_AGEMA_signal_3556), .Q (new_AGEMA_signal_3557) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C (clk), .D (new_AGEMA_signal_3564), .Q (new_AGEMA_signal_3565) ) ;
    buf_clk new_AGEMA_reg_buffer_2213 ( .C (clk), .D (new_AGEMA_signal_3572), .Q (new_AGEMA_signal_3573) ) ;
    buf_clk new_AGEMA_reg_buffer_2221 ( .C (clk), .D (new_AGEMA_signal_3580), .Q (new_AGEMA_signal_3581) ) ;
    buf_clk new_AGEMA_reg_buffer_2229 ( .C (clk), .D (new_AGEMA_signal_3588), .Q (new_AGEMA_signal_3589) ) ;
    buf_clk new_AGEMA_reg_buffer_2237 ( .C (clk), .D (new_AGEMA_signal_3596), .Q (new_AGEMA_signal_3597) ) ;
    buf_clk new_AGEMA_reg_buffer_2245 ( .C (clk), .D (new_AGEMA_signal_3604), .Q (new_AGEMA_signal_3605) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C (clk), .D (new_AGEMA_signal_3612), .Q (new_AGEMA_signal_3613) ) ;
    buf_clk new_AGEMA_reg_buffer_2261 ( .C (clk), .D (new_AGEMA_signal_3620), .Q (new_AGEMA_signal_3621) ) ;
    buf_clk new_AGEMA_reg_buffer_2269 ( .C (clk), .D (new_AGEMA_signal_3628), .Q (new_AGEMA_signal_3629) ) ;
    buf_clk new_AGEMA_reg_buffer_2277 ( .C (clk), .D (new_AGEMA_signal_3636), .Q (new_AGEMA_signal_3637) ) ;
    buf_clk new_AGEMA_reg_buffer_2285 ( .C (clk), .D (new_AGEMA_signal_3644), .Q (new_AGEMA_signal_3645) ) ;
    buf_clk new_AGEMA_reg_buffer_2293 ( .C (clk), .D (new_AGEMA_signal_3652), .Q (new_AGEMA_signal_3653) ) ;
    buf_clk new_AGEMA_reg_buffer_2301 ( .C (clk), .D (new_AGEMA_signal_3660), .Q (new_AGEMA_signal_3661) ) ;
    buf_clk new_AGEMA_reg_buffer_2309 ( .C (clk), .D (new_AGEMA_signal_3668), .Q (new_AGEMA_signal_3669) ) ;
    buf_clk new_AGEMA_reg_buffer_2317 ( .C (clk), .D (new_AGEMA_signal_3676), .Q (new_AGEMA_signal_3677) ) ;
    buf_clk new_AGEMA_reg_buffer_2325 ( .C (clk), .D (new_AGEMA_signal_3684), .Q (new_AGEMA_signal_3685) ) ;
    buf_clk new_AGEMA_reg_buffer_2333 ( .C (clk), .D (new_AGEMA_signal_3692), .Q (new_AGEMA_signal_3693) ) ;
    buf_clk new_AGEMA_reg_buffer_2341 ( .C (clk), .D (new_AGEMA_signal_3700), .Q (new_AGEMA_signal_3701) ) ;
    buf_clk new_AGEMA_reg_buffer_2349 ( .C (clk), .D (new_AGEMA_signal_3708), .Q (new_AGEMA_signal_3709) ) ;
    buf_clk new_AGEMA_reg_buffer_2357 ( .C (clk), .D (new_AGEMA_signal_3716), .Q (new_AGEMA_signal_3717) ) ;
    buf_clk new_AGEMA_reg_buffer_2365 ( .C (clk), .D (new_AGEMA_signal_3724), .Q (new_AGEMA_signal_3725) ) ;
    buf_clk new_AGEMA_reg_buffer_2373 ( .C (clk), .D (new_AGEMA_signal_3732), .Q (new_AGEMA_signal_3733) ) ;
    buf_clk new_AGEMA_reg_buffer_2381 ( .C (clk), .D (new_AGEMA_signal_3740), .Q (new_AGEMA_signal_3741) ) ;
    buf_clk new_AGEMA_reg_buffer_2389 ( .C (clk), .D (new_AGEMA_signal_3748), .Q (new_AGEMA_signal_3749) ) ;
    buf_clk new_AGEMA_reg_buffer_2397 ( .C (clk), .D (new_AGEMA_signal_3756), .Q (new_AGEMA_signal_3757) ) ;
    buf_clk new_AGEMA_reg_buffer_2405 ( .C (clk), .D (new_AGEMA_signal_3764), .Q (new_AGEMA_signal_3765) ) ;
    buf_clk new_AGEMA_reg_buffer_2413 ( .C (clk), .D (new_AGEMA_signal_3772), .Q (new_AGEMA_signal_3773) ) ;
    buf_clk new_AGEMA_reg_buffer_2421 ( .C (clk), .D (new_AGEMA_signal_3780), .Q (new_AGEMA_signal_3781) ) ;
    buf_clk new_AGEMA_reg_buffer_2429 ( .C (clk), .D (new_AGEMA_signal_3788), .Q (new_AGEMA_signal_3789) ) ;
    buf_clk new_AGEMA_reg_buffer_2437 ( .C (clk), .D (new_AGEMA_signal_3796), .Q (new_AGEMA_signal_3797) ) ;
    buf_clk new_AGEMA_reg_buffer_2445 ( .C (clk), .D (new_AGEMA_signal_3804), .Q (new_AGEMA_signal_3805) ) ;
    buf_clk new_AGEMA_reg_buffer_2453 ( .C (clk), .D (new_AGEMA_signal_3812), .Q (new_AGEMA_signal_3813) ) ;
    buf_clk new_AGEMA_reg_buffer_2461 ( .C (clk), .D (new_AGEMA_signal_3820), .Q (new_AGEMA_signal_3821) ) ;
    buf_clk new_AGEMA_reg_buffer_2469 ( .C (clk), .D (new_AGEMA_signal_3828), .Q (new_AGEMA_signal_3829) ) ;
    buf_clk new_AGEMA_reg_buffer_2477 ( .C (clk), .D (new_AGEMA_signal_3836), .Q (new_AGEMA_signal_3837) ) ;
    buf_clk new_AGEMA_reg_buffer_2485 ( .C (clk), .D (new_AGEMA_signal_3844), .Q (new_AGEMA_signal_3845) ) ;
    buf_clk new_AGEMA_reg_buffer_2493 ( .C (clk), .D (new_AGEMA_signal_3852), .Q (new_AGEMA_signal_3853) ) ;
    buf_clk new_AGEMA_reg_buffer_2501 ( .C (clk), .D (new_AGEMA_signal_3860), .Q (new_AGEMA_signal_3861) ) ;
    buf_clk new_AGEMA_reg_buffer_2509 ( .C (clk), .D (new_AGEMA_signal_3868), .Q (new_AGEMA_signal_3869) ) ;
    buf_clk new_AGEMA_reg_buffer_2517 ( .C (clk), .D (new_AGEMA_signal_3876), .Q (new_AGEMA_signal_3877) ) ;
    buf_clk new_AGEMA_reg_buffer_2525 ( .C (clk), .D (new_AGEMA_signal_3884), .Q (new_AGEMA_signal_3885) ) ;
    buf_clk new_AGEMA_reg_buffer_2533 ( .C (clk), .D (new_AGEMA_signal_3892), .Q (new_AGEMA_signal_3893) ) ;
    buf_clk new_AGEMA_reg_buffer_2541 ( .C (clk), .D (new_AGEMA_signal_3900), .Q (new_AGEMA_signal_3901) ) ;
    buf_clk new_AGEMA_reg_buffer_2549 ( .C (clk), .D (new_AGEMA_signal_3908), .Q (new_AGEMA_signal_3909) ) ;
    buf_clk new_AGEMA_reg_buffer_2557 ( .C (clk), .D (new_AGEMA_signal_3916), .Q (new_AGEMA_signal_3917) ) ;
    buf_clk new_AGEMA_reg_buffer_2565 ( .C (clk), .D (new_AGEMA_signal_3924), .Q (new_AGEMA_signal_3925) ) ;
    buf_clk new_AGEMA_reg_buffer_2573 ( .C (clk), .D (new_AGEMA_signal_3932), .Q (new_AGEMA_signal_3933) ) ;
    buf_clk new_AGEMA_reg_buffer_2581 ( .C (clk), .D (new_AGEMA_signal_3940), .Q (new_AGEMA_signal_3941) ) ;
    buf_clk new_AGEMA_reg_buffer_2589 ( .C (clk), .D (new_AGEMA_signal_3948), .Q (new_AGEMA_signal_3949) ) ;
    buf_clk new_AGEMA_reg_buffer_2597 ( .C (clk), .D (new_AGEMA_signal_3956), .Q (new_AGEMA_signal_3957) ) ;
    buf_clk new_AGEMA_reg_buffer_2605 ( .C (clk), .D (new_AGEMA_signal_3964), .Q (new_AGEMA_signal_3965) ) ;
    buf_clk new_AGEMA_reg_buffer_2613 ( .C (clk), .D (new_AGEMA_signal_3972), .Q (new_AGEMA_signal_3973) ) ;
    buf_clk new_AGEMA_reg_buffer_2621 ( .C (clk), .D (new_AGEMA_signal_3980), .Q (new_AGEMA_signal_3981) ) ;
    buf_clk new_AGEMA_reg_buffer_2629 ( .C (clk), .D (new_AGEMA_signal_3988), .Q (new_AGEMA_signal_3989) ) ;
    buf_clk new_AGEMA_reg_buffer_2637 ( .C (clk), .D (new_AGEMA_signal_3996), .Q (new_AGEMA_signal_3997) ) ;
    buf_clk new_AGEMA_reg_buffer_2645 ( .C (clk), .D (new_AGEMA_signal_4004), .Q (new_AGEMA_signal_4005) ) ;
    buf_clk new_AGEMA_reg_buffer_2653 ( .C (clk), .D (new_AGEMA_signal_4012), .Q (new_AGEMA_signal_4013) ) ;
    buf_clk new_AGEMA_reg_buffer_2661 ( .C (clk), .D (new_AGEMA_signal_4020), .Q (new_AGEMA_signal_4021) ) ;
    buf_clk new_AGEMA_reg_buffer_2669 ( .C (clk), .D (new_AGEMA_signal_4028), .Q (new_AGEMA_signal_4029) ) ;
    buf_clk new_AGEMA_reg_buffer_2677 ( .C (clk), .D (new_AGEMA_signal_4036), .Q (new_AGEMA_signal_4037) ) ;
    buf_clk new_AGEMA_reg_buffer_2685 ( .C (clk), .D (new_AGEMA_signal_4044), .Q (new_AGEMA_signal_4045) ) ;
    buf_clk new_AGEMA_reg_buffer_2693 ( .C (clk), .D (new_AGEMA_signal_4052), .Q (new_AGEMA_signal_4053) ) ;
    buf_clk new_AGEMA_reg_buffer_2701 ( .C (clk), .D (new_AGEMA_signal_4060), .Q (new_AGEMA_signal_4061) ) ;
    buf_clk new_AGEMA_reg_buffer_2709 ( .C (clk), .D (new_AGEMA_signal_4068), .Q (new_AGEMA_signal_4069) ) ;
    buf_clk new_AGEMA_reg_buffer_2717 ( .C (clk), .D (new_AGEMA_signal_4076), .Q (new_AGEMA_signal_4077) ) ;
    buf_clk new_AGEMA_reg_buffer_2725 ( .C (clk), .D (new_AGEMA_signal_4084), .Q (new_AGEMA_signal_4085) ) ;
    buf_clk new_AGEMA_reg_buffer_2733 ( .C (clk), .D (new_AGEMA_signal_4092), .Q (new_AGEMA_signal_4093) ) ;
    buf_clk new_AGEMA_reg_buffer_2741 ( .C (clk), .D (new_AGEMA_signal_4100), .Q (new_AGEMA_signal_4101) ) ;
    buf_clk new_AGEMA_reg_buffer_2749 ( .C (clk), .D (new_AGEMA_signal_4108), .Q (new_AGEMA_signal_4109) ) ;
    buf_clk new_AGEMA_reg_buffer_2757 ( .C (clk), .D (new_AGEMA_signal_4116), .Q (new_AGEMA_signal_4117) ) ;
    buf_clk new_AGEMA_reg_buffer_2765 ( .C (clk), .D (new_AGEMA_signal_4124), .Q (new_AGEMA_signal_4125) ) ;
    buf_clk new_AGEMA_reg_buffer_2773 ( .C (clk), .D (new_AGEMA_signal_4132), .Q (new_AGEMA_signal_4133) ) ;
    buf_clk new_AGEMA_reg_buffer_2781 ( .C (clk), .D (new_AGEMA_signal_4140), .Q (new_AGEMA_signal_4141) ) ;
    buf_clk new_AGEMA_reg_buffer_2789 ( .C (clk), .D (new_AGEMA_signal_4148), .Q (new_AGEMA_signal_4149) ) ;
    buf_clk new_AGEMA_reg_buffer_2797 ( .C (clk), .D (new_AGEMA_signal_4156), .Q (new_AGEMA_signal_4157) ) ;
    buf_clk new_AGEMA_reg_buffer_2805 ( .C (clk), .D (new_AGEMA_signal_4164), .Q (new_AGEMA_signal_4165) ) ;
    buf_clk new_AGEMA_reg_buffer_2813 ( .C (clk), .D (new_AGEMA_signal_4172), .Q (new_AGEMA_signal_4173) ) ;
    buf_clk new_AGEMA_reg_buffer_2821 ( .C (clk), .D (new_AGEMA_signal_4180), .Q (new_AGEMA_signal_4181) ) ;
    buf_clk new_AGEMA_reg_buffer_2829 ( .C (clk), .D (new_AGEMA_signal_4188), .Q (new_AGEMA_signal_4189) ) ;
    buf_clk new_AGEMA_reg_buffer_2837 ( .C (clk), .D (new_AGEMA_signal_4196), .Q (new_AGEMA_signal_4197) ) ;
    buf_clk new_AGEMA_reg_buffer_2845 ( .C (clk), .D (new_AGEMA_signal_4204), .Q (new_AGEMA_signal_4205) ) ;
    buf_clk new_AGEMA_reg_buffer_2853 ( .C (clk), .D (new_AGEMA_signal_4212), .Q (new_AGEMA_signal_4213) ) ;
    buf_clk new_AGEMA_reg_buffer_2861 ( .C (clk), .D (new_AGEMA_signal_4220), .Q (new_AGEMA_signal_4221) ) ;
    buf_clk new_AGEMA_reg_buffer_2869 ( .C (clk), .D (new_AGEMA_signal_4228), .Q (new_AGEMA_signal_4229) ) ;
    buf_clk new_AGEMA_reg_buffer_2877 ( .C (clk), .D (new_AGEMA_signal_4236), .Q (new_AGEMA_signal_4237) ) ;
    buf_clk new_AGEMA_reg_buffer_2885 ( .C (clk), .D (new_AGEMA_signal_4244), .Q (new_AGEMA_signal_4245) ) ;
    buf_clk new_AGEMA_reg_buffer_2893 ( .C (clk), .D (new_AGEMA_signal_4252), .Q (new_AGEMA_signal_4253) ) ;
    buf_clk new_AGEMA_reg_buffer_2901 ( .C (clk), .D (new_AGEMA_signal_4260), .Q (new_AGEMA_signal_4261) ) ;
    buf_clk new_AGEMA_reg_buffer_2909 ( .C (clk), .D (new_AGEMA_signal_4268), .Q (new_AGEMA_signal_4269) ) ;
    buf_clk new_AGEMA_reg_buffer_2917 ( .C (clk), .D (new_AGEMA_signal_4276), .Q (new_AGEMA_signal_4277) ) ;
    buf_clk new_AGEMA_reg_buffer_2925 ( .C (clk), .D (new_AGEMA_signal_4284), .Q (new_AGEMA_signal_4285) ) ;
    buf_clk new_AGEMA_reg_buffer_2933 ( .C (clk), .D (new_AGEMA_signal_4292), .Q (new_AGEMA_signal_4293) ) ;
    buf_clk new_AGEMA_reg_buffer_2941 ( .C (clk), .D (new_AGEMA_signal_4300), .Q (new_AGEMA_signal_4301) ) ;
    buf_clk new_AGEMA_reg_buffer_2949 ( .C (clk), .D (new_AGEMA_signal_4308), .Q (new_AGEMA_signal_4309) ) ;
    buf_clk new_AGEMA_reg_buffer_2957 ( .C (clk), .D (new_AGEMA_signal_4316), .Q (new_AGEMA_signal_4317) ) ;
    buf_clk new_AGEMA_reg_buffer_2965 ( .C (clk), .D (new_AGEMA_signal_4324), .Q (new_AGEMA_signal_4325) ) ;
    buf_clk new_AGEMA_reg_buffer_2973 ( .C (clk), .D (new_AGEMA_signal_4332), .Q (new_AGEMA_signal_4333) ) ;
    buf_clk new_AGEMA_reg_buffer_2981 ( .C (clk), .D (new_AGEMA_signal_4340), .Q (new_AGEMA_signal_4341) ) ;
    buf_clk new_AGEMA_reg_buffer_2989 ( .C (clk), .D (new_AGEMA_signal_4348), .Q (new_AGEMA_signal_4349) ) ;
    buf_clk new_AGEMA_reg_buffer_2997 ( .C (clk), .D (new_AGEMA_signal_4356), .Q (new_AGEMA_signal_4357) ) ;
    buf_clk new_AGEMA_reg_buffer_3005 ( .C (clk), .D (new_AGEMA_signal_4364), .Q (new_AGEMA_signal_4365) ) ;
    buf_clk new_AGEMA_reg_buffer_3013 ( .C (clk), .D (new_AGEMA_signal_4372), .Q (new_AGEMA_signal_4373) ) ;
    buf_clk new_AGEMA_reg_buffer_3021 ( .C (clk), .D (new_AGEMA_signal_4380), .Q (new_AGEMA_signal_4381) ) ;
    buf_clk new_AGEMA_reg_buffer_3029 ( .C (clk), .D (new_AGEMA_signal_4388), .Q (new_AGEMA_signal_4389) ) ;
    buf_clk new_AGEMA_reg_buffer_3037 ( .C (clk), .D (new_AGEMA_signal_4396), .Q (new_AGEMA_signal_4397) ) ;
    buf_clk new_AGEMA_reg_buffer_3045 ( .C (clk), .D (new_AGEMA_signal_4404), .Q (new_AGEMA_signal_4405) ) ;
    buf_clk new_AGEMA_reg_buffer_3053 ( .C (clk), .D (new_AGEMA_signal_4412), .Q (new_AGEMA_signal_4413) ) ;
    buf_clk new_AGEMA_reg_buffer_3061 ( .C (clk), .D (new_AGEMA_signal_4420), .Q (new_AGEMA_signal_4421) ) ;
    buf_clk new_AGEMA_reg_buffer_3071 ( .C (clk), .D (SubCellInst_SboxInst_0_n13), .Q (new_AGEMA_signal_4431) ) ;
    buf_clk new_AGEMA_reg_buffer_3075 ( .C (clk), .D (new_AGEMA_signal_1152), .Q (new_AGEMA_signal_4435) ) ;
    buf_clk new_AGEMA_reg_buffer_3083 ( .C (clk), .D (SubCellInst_SboxInst_1_n13), .Q (new_AGEMA_signal_4443) ) ;
    buf_clk new_AGEMA_reg_buffer_3087 ( .C (clk), .D (new_AGEMA_signal_1158), .Q (new_AGEMA_signal_4447) ) ;
    buf_clk new_AGEMA_reg_buffer_3095 ( .C (clk), .D (SubCellInst_SboxInst_2_n13), .Q (new_AGEMA_signal_4455) ) ;
    buf_clk new_AGEMA_reg_buffer_3099 ( .C (clk), .D (new_AGEMA_signal_1164), .Q (new_AGEMA_signal_4459) ) ;
    buf_clk new_AGEMA_reg_buffer_3107 ( .C (clk), .D (SubCellInst_SboxInst_3_n13), .Q (new_AGEMA_signal_4467) ) ;
    buf_clk new_AGEMA_reg_buffer_3111 ( .C (clk), .D (new_AGEMA_signal_1170), .Q (new_AGEMA_signal_4471) ) ;
    buf_clk new_AGEMA_reg_buffer_3119 ( .C (clk), .D (SubCellInst_SboxInst_4_n13), .Q (new_AGEMA_signal_4479) ) ;
    buf_clk new_AGEMA_reg_buffer_3123 ( .C (clk), .D (new_AGEMA_signal_1176), .Q (new_AGEMA_signal_4483) ) ;
    buf_clk new_AGEMA_reg_buffer_3131 ( .C (clk), .D (SubCellInst_SboxInst_5_n13), .Q (new_AGEMA_signal_4491) ) ;
    buf_clk new_AGEMA_reg_buffer_3135 ( .C (clk), .D (new_AGEMA_signal_1182), .Q (new_AGEMA_signal_4495) ) ;
    buf_clk new_AGEMA_reg_buffer_3143 ( .C (clk), .D (SubCellInst_SboxInst_6_n13), .Q (new_AGEMA_signal_4503) ) ;
    buf_clk new_AGEMA_reg_buffer_3147 ( .C (clk), .D (new_AGEMA_signal_1188), .Q (new_AGEMA_signal_4507) ) ;
    buf_clk new_AGEMA_reg_buffer_3155 ( .C (clk), .D (SubCellInst_SboxInst_7_n13), .Q (new_AGEMA_signal_4515) ) ;
    buf_clk new_AGEMA_reg_buffer_3159 ( .C (clk), .D (new_AGEMA_signal_1194), .Q (new_AGEMA_signal_4519) ) ;
    buf_clk new_AGEMA_reg_buffer_3167 ( .C (clk), .D (SubCellInst_SboxInst_8_n13), .Q (new_AGEMA_signal_4527) ) ;
    buf_clk new_AGEMA_reg_buffer_3171 ( .C (clk), .D (new_AGEMA_signal_1200), .Q (new_AGEMA_signal_4531) ) ;
    buf_clk new_AGEMA_reg_buffer_3179 ( .C (clk), .D (SubCellInst_SboxInst_9_n13), .Q (new_AGEMA_signal_4539) ) ;
    buf_clk new_AGEMA_reg_buffer_3183 ( .C (clk), .D (new_AGEMA_signal_1206), .Q (new_AGEMA_signal_4543) ) ;
    buf_clk new_AGEMA_reg_buffer_3191 ( .C (clk), .D (SubCellInst_SboxInst_10_n13), .Q (new_AGEMA_signal_4551) ) ;
    buf_clk new_AGEMA_reg_buffer_3195 ( .C (clk), .D (new_AGEMA_signal_1212), .Q (new_AGEMA_signal_4555) ) ;
    buf_clk new_AGEMA_reg_buffer_3203 ( .C (clk), .D (SubCellInst_SboxInst_11_n13), .Q (new_AGEMA_signal_4563) ) ;
    buf_clk new_AGEMA_reg_buffer_3207 ( .C (clk), .D (new_AGEMA_signal_1218), .Q (new_AGEMA_signal_4567) ) ;
    buf_clk new_AGEMA_reg_buffer_3215 ( .C (clk), .D (SubCellInst_SboxInst_12_n13), .Q (new_AGEMA_signal_4575) ) ;
    buf_clk new_AGEMA_reg_buffer_3219 ( .C (clk), .D (new_AGEMA_signal_1224), .Q (new_AGEMA_signal_4579) ) ;
    buf_clk new_AGEMA_reg_buffer_3227 ( .C (clk), .D (SubCellInst_SboxInst_13_n13), .Q (new_AGEMA_signal_4587) ) ;
    buf_clk new_AGEMA_reg_buffer_3231 ( .C (clk), .D (new_AGEMA_signal_1230), .Q (new_AGEMA_signal_4591) ) ;
    buf_clk new_AGEMA_reg_buffer_3239 ( .C (clk), .D (SubCellInst_SboxInst_14_n13), .Q (new_AGEMA_signal_4599) ) ;
    buf_clk new_AGEMA_reg_buffer_3243 ( .C (clk), .D (new_AGEMA_signal_1236), .Q (new_AGEMA_signal_4603) ) ;
    buf_clk new_AGEMA_reg_buffer_3251 ( .C (clk), .D (SubCellInst_SboxInst_15_n13), .Q (new_AGEMA_signal_4611) ) ;
    buf_clk new_AGEMA_reg_buffer_3255 ( .C (clk), .D (new_AGEMA_signal_1242), .Q (new_AGEMA_signal_4615) ) ;
    buf_clk new_AGEMA_reg_buffer_3389 ( .C (clk), .D (new_AGEMA_signal_4748), .Q (new_AGEMA_signal_4749) ) ;
    buf_clk new_AGEMA_reg_buffer_3397 ( .C (clk), .D (new_AGEMA_signal_4756), .Q (new_AGEMA_signal_4757) ) ;
    buf_clk new_AGEMA_reg_buffer_3405 ( .C (clk), .D (new_AGEMA_signal_4764), .Q (new_AGEMA_signal_4765) ) ;
    buf_clk new_AGEMA_reg_buffer_3413 ( .C (clk), .D (new_AGEMA_signal_4772), .Q (new_AGEMA_signal_4773) ) ;
    buf_clk new_AGEMA_reg_buffer_3421 ( .C (clk), .D (new_AGEMA_signal_4780), .Q (new_AGEMA_signal_4781) ) ;
    buf_clk new_AGEMA_reg_buffer_3429 ( .C (clk), .D (new_AGEMA_signal_4788), .Q (new_AGEMA_signal_4789) ) ;
    buf_clk new_AGEMA_reg_buffer_3437 ( .C (clk), .D (new_AGEMA_signal_4796), .Q (new_AGEMA_signal_4797) ) ;
    buf_clk new_AGEMA_reg_buffer_3445 ( .C (clk), .D (new_AGEMA_signal_4804), .Q (new_AGEMA_signal_4805) ) ;
    buf_clk new_AGEMA_reg_buffer_3453 ( .C (clk), .D (new_AGEMA_signal_4812), .Q (new_AGEMA_signal_4813) ) ;
    buf_clk new_AGEMA_reg_buffer_3461 ( .C (clk), .D (new_AGEMA_signal_4820), .Q (new_AGEMA_signal_4821) ) ;

    /* cells in depth 4 */
    or_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U18 ( .a ({new_AGEMA_signal_1152, SubCellInst_SboxInst_0_n13}), .b ({new_AGEMA_signal_2182, new_AGEMA_signal_2180}), .clk (clk), .r (Fresh[96]), .c ({new_AGEMA_signal_1292, SubCellInst_SboxInst_0_n14}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U15 ( .a ({new_AGEMA_signal_1021, SubCellInst_SboxInst_0_n10}), .b ({new_AGEMA_signal_2186, new_AGEMA_signal_2184}), .clk (clk), .r (Fresh[97]), .c ({new_AGEMA_signal_1147, SubCellInst_SboxInst_0_n11}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U11 ( .a ({new_AGEMA_signal_2190, new_AGEMA_signal_2188}), .b ({new_AGEMA_signal_1149, SubCellInst_SboxInst_0_n4}), .clk (clk), .r (Fresh[98]), .c ({new_AGEMA_signal_1294, SubCellInst_SboxInst_0_n5}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U6 ( .a ({new_AGEMA_signal_2194, new_AGEMA_signal_2192}), .b ({new_AGEMA_signal_1023, SubCellInst_SboxInst_0_n1}), .clk (clk), .r (Fresh[99]), .c ({new_AGEMA_signal_1151, SubCellInst_SboxInst_0_n2}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U18 ( .a ({new_AGEMA_signal_1158, SubCellInst_SboxInst_1_n13}), .b ({new_AGEMA_signal_2198, new_AGEMA_signal_2196}), .clk (clk), .r (Fresh[100]), .c ({new_AGEMA_signal_1297, SubCellInst_SboxInst_1_n14}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U15 ( .a ({new_AGEMA_signal_1029, SubCellInst_SboxInst_1_n10}), .b ({new_AGEMA_signal_2202, new_AGEMA_signal_2200}), .clk (clk), .r (Fresh[101]), .c ({new_AGEMA_signal_1153, SubCellInst_SboxInst_1_n11}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U11 ( .a ({new_AGEMA_signal_2206, new_AGEMA_signal_2204}), .b ({new_AGEMA_signal_1155, SubCellInst_SboxInst_1_n4}), .clk (clk), .r (Fresh[102]), .c ({new_AGEMA_signal_1299, SubCellInst_SboxInst_1_n5}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U6 ( .a ({new_AGEMA_signal_2210, new_AGEMA_signal_2208}), .b ({new_AGEMA_signal_1031, SubCellInst_SboxInst_1_n1}), .clk (clk), .r (Fresh[103]), .c ({new_AGEMA_signal_1157, SubCellInst_SboxInst_1_n2}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U18 ( .a ({new_AGEMA_signal_1164, SubCellInst_SboxInst_2_n13}), .b ({new_AGEMA_signal_2214, new_AGEMA_signal_2212}), .clk (clk), .r (Fresh[104]), .c ({new_AGEMA_signal_1302, SubCellInst_SboxInst_2_n14}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U15 ( .a ({new_AGEMA_signal_1037, SubCellInst_SboxInst_2_n10}), .b ({new_AGEMA_signal_2218, new_AGEMA_signal_2216}), .clk (clk), .r (Fresh[105]), .c ({new_AGEMA_signal_1159, SubCellInst_SboxInst_2_n11}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U11 ( .a ({new_AGEMA_signal_2222, new_AGEMA_signal_2220}), .b ({new_AGEMA_signal_1161, SubCellInst_SboxInst_2_n4}), .clk (clk), .r (Fresh[106]), .c ({new_AGEMA_signal_1304, SubCellInst_SboxInst_2_n5}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U6 ( .a ({new_AGEMA_signal_2226, new_AGEMA_signal_2224}), .b ({new_AGEMA_signal_1039, SubCellInst_SboxInst_2_n1}), .clk (clk), .r (Fresh[107]), .c ({new_AGEMA_signal_1163, SubCellInst_SboxInst_2_n2}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U18 ( .a ({new_AGEMA_signal_1170, SubCellInst_SboxInst_3_n13}), .b ({new_AGEMA_signal_2230, new_AGEMA_signal_2228}), .clk (clk), .r (Fresh[108]), .c ({new_AGEMA_signal_1307, SubCellInst_SboxInst_3_n14}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U15 ( .a ({new_AGEMA_signal_1045, SubCellInst_SboxInst_3_n10}), .b ({new_AGEMA_signal_2234, new_AGEMA_signal_2232}), .clk (clk), .r (Fresh[109]), .c ({new_AGEMA_signal_1165, SubCellInst_SboxInst_3_n11}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U11 ( .a ({new_AGEMA_signal_2238, new_AGEMA_signal_2236}), .b ({new_AGEMA_signal_1167, SubCellInst_SboxInst_3_n4}), .clk (clk), .r (Fresh[110]), .c ({new_AGEMA_signal_1309, SubCellInst_SboxInst_3_n5}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U6 ( .a ({new_AGEMA_signal_2242, new_AGEMA_signal_2240}), .b ({new_AGEMA_signal_1047, SubCellInst_SboxInst_3_n1}), .clk (clk), .r (Fresh[111]), .c ({new_AGEMA_signal_1169, SubCellInst_SboxInst_3_n2}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U18 ( .a ({new_AGEMA_signal_1176, SubCellInst_SboxInst_4_n13}), .b ({new_AGEMA_signal_2246, new_AGEMA_signal_2244}), .clk (clk), .r (Fresh[112]), .c ({new_AGEMA_signal_1312, SubCellInst_SboxInst_4_n14}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U15 ( .a ({new_AGEMA_signal_1053, SubCellInst_SboxInst_4_n10}), .b ({new_AGEMA_signal_2250, new_AGEMA_signal_2248}), .clk (clk), .r (Fresh[113]), .c ({new_AGEMA_signal_1171, SubCellInst_SboxInst_4_n11}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U11 ( .a ({new_AGEMA_signal_2254, new_AGEMA_signal_2252}), .b ({new_AGEMA_signal_1173, SubCellInst_SboxInst_4_n4}), .clk (clk), .r (Fresh[114]), .c ({new_AGEMA_signal_1314, SubCellInst_SboxInst_4_n5}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U6 ( .a ({new_AGEMA_signal_2258, new_AGEMA_signal_2256}), .b ({new_AGEMA_signal_1055, SubCellInst_SboxInst_4_n1}), .clk (clk), .r (Fresh[115]), .c ({new_AGEMA_signal_1175, SubCellInst_SboxInst_4_n2}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U18 ( .a ({new_AGEMA_signal_1182, SubCellInst_SboxInst_5_n13}), .b ({new_AGEMA_signal_2262, new_AGEMA_signal_2260}), .clk (clk), .r (Fresh[116]), .c ({new_AGEMA_signal_1317, SubCellInst_SboxInst_5_n14}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U15 ( .a ({new_AGEMA_signal_1061, SubCellInst_SboxInst_5_n10}), .b ({new_AGEMA_signal_2266, new_AGEMA_signal_2264}), .clk (clk), .r (Fresh[117]), .c ({new_AGEMA_signal_1177, SubCellInst_SboxInst_5_n11}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U11 ( .a ({new_AGEMA_signal_2270, new_AGEMA_signal_2268}), .b ({new_AGEMA_signal_1179, SubCellInst_SboxInst_5_n4}), .clk (clk), .r (Fresh[118]), .c ({new_AGEMA_signal_1319, SubCellInst_SboxInst_5_n5}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U6 ( .a ({new_AGEMA_signal_2274, new_AGEMA_signal_2272}), .b ({new_AGEMA_signal_1063, SubCellInst_SboxInst_5_n1}), .clk (clk), .r (Fresh[119]), .c ({new_AGEMA_signal_1181, SubCellInst_SboxInst_5_n2}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U18 ( .a ({new_AGEMA_signal_1188, SubCellInst_SboxInst_6_n13}), .b ({new_AGEMA_signal_2278, new_AGEMA_signal_2276}), .clk (clk), .r (Fresh[120]), .c ({new_AGEMA_signal_1322, SubCellInst_SboxInst_6_n14}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U15 ( .a ({new_AGEMA_signal_1069, SubCellInst_SboxInst_6_n10}), .b ({new_AGEMA_signal_2282, new_AGEMA_signal_2280}), .clk (clk), .r (Fresh[121]), .c ({new_AGEMA_signal_1183, SubCellInst_SboxInst_6_n11}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U11 ( .a ({new_AGEMA_signal_2286, new_AGEMA_signal_2284}), .b ({new_AGEMA_signal_1185, SubCellInst_SboxInst_6_n4}), .clk (clk), .r (Fresh[122]), .c ({new_AGEMA_signal_1324, SubCellInst_SboxInst_6_n5}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U6 ( .a ({new_AGEMA_signal_2290, new_AGEMA_signal_2288}), .b ({new_AGEMA_signal_1071, SubCellInst_SboxInst_6_n1}), .clk (clk), .r (Fresh[123]), .c ({new_AGEMA_signal_1187, SubCellInst_SboxInst_6_n2}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U18 ( .a ({new_AGEMA_signal_1194, SubCellInst_SboxInst_7_n13}), .b ({new_AGEMA_signal_2294, new_AGEMA_signal_2292}), .clk (clk), .r (Fresh[124]), .c ({new_AGEMA_signal_1327, SubCellInst_SboxInst_7_n14}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U15 ( .a ({new_AGEMA_signal_1077, SubCellInst_SboxInst_7_n10}), .b ({new_AGEMA_signal_2298, new_AGEMA_signal_2296}), .clk (clk), .r (Fresh[125]), .c ({new_AGEMA_signal_1189, SubCellInst_SboxInst_7_n11}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U11 ( .a ({new_AGEMA_signal_2302, new_AGEMA_signal_2300}), .b ({new_AGEMA_signal_1191, SubCellInst_SboxInst_7_n4}), .clk (clk), .r (Fresh[126]), .c ({new_AGEMA_signal_1329, SubCellInst_SboxInst_7_n5}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U6 ( .a ({new_AGEMA_signal_2306, new_AGEMA_signal_2304}), .b ({new_AGEMA_signal_1079, SubCellInst_SboxInst_7_n1}), .clk (clk), .r (Fresh[127]), .c ({new_AGEMA_signal_1193, SubCellInst_SboxInst_7_n2}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U18 ( .a ({new_AGEMA_signal_1200, SubCellInst_SboxInst_8_n13}), .b ({new_AGEMA_signal_2310, new_AGEMA_signal_2308}), .clk (clk), .r (Fresh[128]), .c ({new_AGEMA_signal_1332, SubCellInst_SboxInst_8_n14}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U15 ( .a ({new_AGEMA_signal_1085, SubCellInst_SboxInst_8_n10}), .b ({new_AGEMA_signal_2314, new_AGEMA_signal_2312}), .clk (clk), .r (Fresh[129]), .c ({new_AGEMA_signal_1195, SubCellInst_SboxInst_8_n11}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U11 ( .a ({new_AGEMA_signal_2318, new_AGEMA_signal_2316}), .b ({new_AGEMA_signal_1197, SubCellInst_SboxInst_8_n4}), .clk (clk), .r (Fresh[130]), .c ({new_AGEMA_signal_1334, SubCellInst_SboxInst_8_n5}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U6 ( .a ({new_AGEMA_signal_2322, new_AGEMA_signal_2320}), .b ({new_AGEMA_signal_1087, SubCellInst_SboxInst_8_n1}), .clk (clk), .r (Fresh[131]), .c ({new_AGEMA_signal_1199, SubCellInst_SboxInst_8_n2}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U18 ( .a ({new_AGEMA_signal_1206, SubCellInst_SboxInst_9_n13}), .b ({new_AGEMA_signal_2326, new_AGEMA_signal_2324}), .clk (clk), .r (Fresh[132]), .c ({new_AGEMA_signal_1337, SubCellInst_SboxInst_9_n14}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U15 ( .a ({new_AGEMA_signal_1093, SubCellInst_SboxInst_9_n10}), .b ({new_AGEMA_signal_2330, new_AGEMA_signal_2328}), .clk (clk), .r (Fresh[133]), .c ({new_AGEMA_signal_1201, SubCellInst_SboxInst_9_n11}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U11 ( .a ({new_AGEMA_signal_2334, new_AGEMA_signal_2332}), .b ({new_AGEMA_signal_1203, SubCellInst_SboxInst_9_n4}), .clk (clk), .r (Fresh[134]), .c ({new_AGEMA_signal_1339, SubCellInst_SboxInst_9_n5}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U6 ( .a ({new_AGEMA_signal_2338, new_AGEMA_signal_2336}), .b ({new_AGEMA_signal_1095, SubCellInst_SboxInst_9_n1}), .clk (clk), .r (Fresh[135]), .c ({new_AGEMA_signal_1205, SubCellInst_SboxInst_9_n2}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U18 ( .a ({new_AGEMA_signal_1212, SubCellInst_SboxInst_10_n13}), .b ({new_AGEMA_signal_2342, new_AGEMA_signal_2340}), .clk (clk), .r (Fresh[136]), .c ({new_AGEMA_signal_1342, SubCellInst_SboxInst_10_n14}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U15 ( .a ({new_AGEMA_signal_1101, SubCellInst_SboxInst_10_n10}), .b ({new_AGEMA_signal_2346, new_AGEMA_signal_2344}), .clk (clk), .r (Fresh[137]), .c ({new_AGEMA_signal_1207, SubCellInst_SboxInst_10_n11}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U11 ( .a ({new_AGEMA_signal_2350, new_AGEMA_signal_2348}), .b ({new_AGEMA_signal_1209, SubCellInst_SboxInst_10_n4}), .clk (clk), .r (Fresh[138]), .c ({new_AGEMA_signal_1344, SubCellInst_SboxInst_10_n5}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U6 ( .a ({new_AGEMA_signal_2354, new_AGEMA_signal_2352}), .b ({new_AGEMA_signal_1103, SubCellInst_SboxInst_10_n1}), .clk (clk), .r (Fresh[139]), .c ({new_AGEMA_signal_1211, SubCellInst_SboxInst_10_n2}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U18 ( .a ({new_AGEMA_signal_1218, SubCellInst_SboxInst_11_n13}), .b ({new_AGEMA_signal_2358, new_AGEMA_signal_2356}), .clk (clk), .r (Fresh[140]), .c ({new_AGEMA_signal_1347, SubCellInst_SboxInst_11_n14}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U15 ( .a ({new_AGEMA_signal_1109, SubCellInst_SboxInst_11_n10}), .b ({new_AGEMA_signal_2362, new_AGEMA_signal_2360}), .clk (clk), .r (Fresh[141]), .c ({new_AGEMA_signal_1213, SubCellInst_SboxInst_11_n11}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U11 ( .a ({new_AGEMA_signal_2366, new_AGEMA_signal_2364}), .b ({new_AGEMA_signal_1215, SubCellInst_SboxInst_11_n4}), .clk (clk), .r (Fresh[142]), .c ({new_AGEMA_signal_1349, SubCellInst_SboxInst_11_n5}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U6 ( .a ({new_AGEMA_signal_2370, new_AGEMA_signal_2368}), .b ({new_AGEMA_signal_1111, SubCellInst_SboxInst_11_n1}), .clk (clk), .r (Fresh[143]), .c ({new_AGEMA_signal_1217, SubCellInst_SboxInst_11_n2}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U18 ( .a ({new_AGEMA_signal_1224, SubCellInst_SboxInst_12_n13}), .b ({new_AGEMA_signal_2374, new_AGEMA_signal_2372}), .clk (clk), .r (Fresh[144]), .c ({new_AGEMA_signal_1352, SubCellInst_SboxInst_12_n14}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U15 ( .a ({new_AGEMA_signal_1117, SubCellInst_SboxInst_12_n10}), .b ({new_AGEMA_signal_2378, new_AGEMA_signal_2376}), .clk (clk), .r (Fresh[145]), .c ({new_AGEMA_signal_1219, SubCellInst_SboxInst_12_n11}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U11 ( .a ({new_AGEMA_signal_2382, new_AGEMA_signal_2380}), .b ({new_AGEMA_signal_1221, SubCellInst_SboxInst_12_n4}), .clk (clk), .r (Fresh[146]), .c ({new_AGEMA_signal_1354, SubCellInst_SboxInst_12_n5}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U6 ( .a ({new_AGEMA_signal_2386, new_AGEMA_signal_2384}), .b ({new_AGEMA_signal_1119, SubCellInst_SboxInst_12_n1}), .clk (clk), .r (Fresh[147]), .c ({new_AGEMA_signal_1223, SubCellInst_SboxInst_12_n2}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U18 ( .a ({new_AGEMA_signal_1230, SubCellInst_SboxInst_13_n13}), .b ({new_AGEMA_signal_2390, new_AGEMA_signal_2388}), .clk (clk), .r (Fresh[148]), .c ({new_AGEMA_signal_1357, SubCellInst_SboxInst_13_n14}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U15 ( .a ({new_AGEMA_signal_1125, SubCellInst_SboxInst_13_n10}), .b ({new_AGEMA_signal_2394, new_AGEMA_signal_2392}), .clk (clk), .r (Fresh[149]), .c ({new_AGEMA_signal_1225, SubCellInst_SboxInst_13_n11}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U11 ( .a ({new_AGEMA_signal_2398, new_AGEMA_signal_2396}), .b ({new_AGEMA_signal_1227, SubCellInst_SboxInst_13_n4}), .clk (clk), .r (Fresh[150]), .c ({new_AGEMA_signal_1359, SubCellInst_SboxInst_13_n5}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U6 ( .a ({new_AGEMA_signal_2402, new_AGEMA_signal_2400}), .b ({new_AGEMA_signal_1127, SubCellInst_SboxInst_13_n1}), .clk (clk), .r (Fresh[151]), .c ({new_AGEMA_signal_1229, SubCellInst_SboxInst_13_n2}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U18 ( .a ({new_AGEMA_signal_1236, SubCellInst_SboxInst_14_n13}), .b ({new_AGEMA_signal_2406, new_AGEMA_signal_2404}), .clk (clk), .r (Fresh[152]), .c ({new_AGEMA_signal_1362, SubCellInst_SboxInst_14_n14}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U15 ( .a ({new_AGEMA_signal_1133, SubCellInst_SboxInst_14_n10}), .b ({new_AGEMA_signal_2410, new_AGEMA_signal_2408}), .clk (clk), .r (Fresh[153]), .c ({new_AGEMA_signal_1231, SubCellInst_SboxInst_14_n11}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U11 ( .a ({new_AGEMA_signal_2414, new_AGEMA_signal_2412}), .b ({new_AGEMA_signal_1233, SubCellInst_SboxInst_14_n4}), .clk (clk), .r (Fresh[154]), .c ({new_AGEMA_signal_1364, SubCellInst_SboxInst_14_n5}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U6 ( .a ({new_AGEMA_signal_2418, new_AGEMA_signal_2416}), .b ({new_AGEMA_signal_1135, SubCellInst_SboxInst_14_n1}), .clk (clk), .r (Fresh[155]), .c ({new_AGEMA_signal_1235, SubCellInst_SboxInst_14_n2}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U18 ( .a ({new_AGEMA_signal_1242, SubCellInst_SboxInst_15_n13}), .b ({new_AGEMA_signal_2422, new_AGEMA_signal_2420}), .clk (clk), .r (Fresh[156]), .c ({new_AGEMA_signal_1367, SubCellInst_SboxInst_15_n14}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U15 ( .a ({new_AGEMA_signal_1141, SubCellInst_SboxInst_15_n10}), .b ({new_AGEMA_signal_2426, new_AGEMA_signal_2424}), .clk (clk), .r (Fresh[157]), .c ({new_AGEMA_signal_1237, SubCellInst_SboxInst_15_n11}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U11 ( .a ({new_AGEMA_signal_2430, new_AGEMA_signal_2428}), .b ({new_AGEMA_signal_1239, SubCellInst_SboxInst_15_n4}), .clk (clk), .r (Fresh[158]), .c ({new_AGEMA_signal_1369, SubCellInst_SboxInst_15_n5}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U6 ( .a ({new_AGEMA_signal_2434, new_AGEMA_signal_2432}), .b ({new_AGEMA_signal_1143, SubCellInst_SboxInst_15_n1}), .clk (clk), .r (Fresh[159]), .c ({new_AGEMA_signal_1241, SubCellInst_SboxInst_15_n2}) ) ;
    buf_clk new_AGEMA_reg_buffer_1078 ( .C (clk), .D (new_AGEMA_signal_2437), .Q (new_AGEMA_signal_2438) ) ;
    buf_clk new_AGEMA_reg_buffer_1084 ( .C (clk), .D (new_AGEMA_signal_2443), .Q (new_AGEMA_signal_2444) ) ;
    buf_clk new_AGEMA_reg_buffer_1090 ( .C (clk), .D (new_AGEMA_signal_2449), .Q (new_AGEMA_signal_2450) ) ;
    buf_clk new_AGEMA_reg_buffer_1096 ( .C (clk), .D (new_AGEMA_signal_2455), .Q (new_AGEMA_signal_2456) ) ;
    buf_clk new_AGEMA_reg_buffer_1102 ( .C (clk), .D (new_AGEMA_signal_2461), .Q (new_AGEMA_signal_2462) ) ;
    buf_clk new_AGEMA_reg_buffer_1108 ( .C (clk), .D (new_AGEMA_signal_2467), .Q (new_AGEMA_signal_2468) ) ;
    buf_clk new_AGEMA_reg_buffer_1114 ( .C (clk), .D (new_AGEMA_signal_2473), .Q (new_AGEMA_signal_2474) ) ;
    buf_clk new_AGEMA_reg_buffer_1120 ( .C (clk), .D (new_AGEMA_signal_2479), .Q (new_AGEMA_signal_2480) ) ;
    buf_clk new_AGEMA_reg_buffer_1126 ( .C (clk), .D (new_AGEMA_signal_2485), .Q (new_AGEMA_signal_2486) ) ;
    buf_clk new_AGEMA_reg_buffer_1132 ( .C (clk), .D (new_AGEMA_signal_2491), .Q (new_AGEMA_signal_2492) ) ;
    buf_clk new_AGEMA_reg_buffer_1138 ( .C (clk), .D (new_AGEMA_signal_2497), .Q (new_AGEMA_signal_2498) ) ;
    buf_clk new_AGEMA_reg_buffer_1144 ( .C (clk), .D (new_AGEMA_signal_2503), .Q (new_AGEMA_signal_2504) ) ;
    buf_clk new_AGEMA_reg_buffer_1150 ( .C (clk), .D (new_AGEMA_signal_2509), .Q (new_AGEMA_signal_2510) ) ;
    buf_clk new_AGEMA_reg_buffer_1156 ( .C (clk), .D (new_AGEMA_signal_2515), .Q (new_AGEMA_signal_2516) ) ;
    buf_clk new_AGEMA_reg_buffer_1162 ( .C (clk), .D (new_AGEMA_signal_2521), .Q (new_AGEMA_signal_2522) ) ;
    buf_clk new_AGEMA_reg_buffer_1168 ( .C (clk), .D (new_AGEMA_signal_2527), .Q (new_AGEMA_signal_2528) ) ;
    buf_clk new_AGEMA_reg_buffer_1174 ( .C (clk), .D (new_AGEMA_signal_2533), .Q (new_AGEMA_signal_2534) ) ;
    buf_clk new_AGEMA_reg_buffer_1180 ( .C (clk), .D (new_AGEMA_signal_2539), .Q (new_AGEMA_signal_2540) ) ;
    buf_clk new_AGEMA_reg_buffer_1186 ( .C (clk), .D (new_AGEMA_signal_2545), .Q (new_AGEMA_signal_2546) ) ;
    buf_clk new_AGEMA_reg_buffer_1192 ( .C (clk), .D (new_AGEMA_signal_2551), .Q (new_AGEMA_signal_2552) ) ;
    buf_clk new_AGEMA_reg_buffer_1198 ( .C (clk), .D (new_AGEMA_signal_2557), .Q (new_AGEMA_signal_2558) ) ;
    buf_clk new_AGEMA_reg_buffer_1204 ( .C (clk), .D (new_AGEMA_signal_2563), .Q (new_AGEMA_signal_2564) ) ;
    buf_clk new_AGEMA_reg_buffer_1210 ( .C (clk), .D (new_AGEMA_signal_2569), .Q (new_AGEMA_signal_2570) ) ;
    buf_clk new_AGEMA_reg_buffer_1216 ( .C (clk), .D (new_AGEMA_signal_2575), .Q (new_AGEMA_signal_2576) ) ;
    buf_clk new_AGEMA_reg_buffer_1222 ( .C (clk), .D (new_AGEMA_signal_2581), .Q (new_AGEMA_signal_2582) ) ;
    buf_clk new_AGEMA_reg_buffer_1228 ( .C (clk), .D (new_AGEMA_signal_2587), .Q (new_AGEMA_signal_2588) ) ;
    buf_clk new_AGEMA_reg_buffer_1234 ( .C (clk), .D (new_AGEMA_signal_2593), .Q (new_AGEMA_signal_2594) ) ;
    buf_clk new_AGEMA_reg_buffer_1240 ( .C (clk), .D (new_AGEMA_signal_2599), .Q (new_AGEMA_signal_2600) ) ;
    buf_clk new_AGEMA_reg_buffer_1246 ( .C (clk), .D (new_AGEMA_signal_2605), .Q (new_AGEMA_signal_2606) ) ;
    buf_clk new_AGEMA_reg_buffer_1252 ( .C (clk), .D (new_AGEMA_signal_2611), .Q (new_AGEMA_signal_2612) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C (clk), .D (new_AGEMA_signal_2617), .Q (new_AGEMA_signal_2618) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C (clk), .D (new_AGEMA_signal_2623), .Q (new_AGEMA_signal_2624) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C (clk), .D (new_AGEMA_signal_2629), .Q (new_AGEMA_signal_2630) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C (clk), .D (new_AGEMA_signal_2635), .Q (new_AGEMA_signal_2636) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C (clk), .D (new_AGEMA_signal_2641), .Q (new_AGEMA_signal_2642) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C (clk), .D (new_AGEMA_signal_2647), .Q (new_AGEMA_signal_2648) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C (clk), .D (new_AGEMA_signal_2653), .Q (new_AGEMA_signal_2654) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C (clk), .D (new_AGEMA_signal_2659), .Q (new_AGEMA_signal_2660) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C (clk), .D (new_AGEMA_signal_2665), .Q (new_AGEMA_signal_2666) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C (clk), .D (new_AGEMA_signal_2671), .Q (new_AGEMA_signal_2672) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C (clk), .D (new_AGEMA_signal_2677), .Q (new_AGEMA_signal_2678) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C (clk), .D (new_AGEMA_signal_2683), .Q (new_AGEMA_signal_2684) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C (clk), .D (new_AGEMA_signal_2689), .Q (new_AGEMA_signal_2690) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C (clk), .D (new_AGEMA_signal_2695), .Q (new_AGEMA_signal_2696) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C (clk), .D (new_AGEMA_signal_2701), .Q (new_AGEMA_signal_2702) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C (clk), .D (new_AGEMA_signal_2707), .Q (new_AGEMA_signal_2708) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C (clk), .D (new_AGEMA_signal_2713), .Q (new_AGEMA_signal_2714) ) ;
    buf_clk new_AGEMA_reg_buffer_1360 ( .C (clk), .D (new_AGEMA_signal_2719), .Q (new_AGEMA_signal_2720) ) ;
    buf_clk new_AGEMA_reg_buffer_1366 ( .C (clk), .D (new_AGEMA_signal_2725), .Q (new_AGEMA_signal_2726) ) ;
    buf_clk new_AGEMA_reg_buffer_1372 ( .C (clk), .D (new_AGEMA_signal_2731), .Q (new_AGEMA_signal_2732) ) ;
    buf_clk new_AGEMA_reg_buffer_1378 ( .C (clk), .D (new_AGEMA_signal_2737), .Q (new_AGEMA_signal_2738) ) ;
    buf_clk new_AGEMA_reg_buffer_1384 ( .C (clk), .D (new_AGEMA_signal_2743), .Q (new_AGEMA_signal_2744) ) ;
    buf_clk new_AGEMA_reg_buffer_1390 ( .C (clk), .D (new_AGEMA_signal_2749), .Q (new_AGEMA_signal_2750) ) ;
    buf_clk new_AGEMA_reg_buffer_1396 ( .C (clk), .D (new_AGEMA_signal_2755), .Q (new_AGEMA_signal_2756) ) ;
    buf_clk new_AGEMA_reg_buffer_1402 ( .C (clk), .D (new_AGEMA_signal_2761), .Q (new_AGEMA_signal_2762) ) ;
    buf_clk new_AGEMA_reg_buffer_1408 ( .C (clk), .D (new_AGEMA_signal_2767), .Q (new_AGEMA_signal_2768) ) ;
    buf_clk new_AGEMA_reg_buffer_1414 ( .C (clk), .D (new_AGEMA_signal_2773), .Q (new_AGEMA_signal_2774) ) ;
    buf_clk new_AGEMA_reg_buffer_1420 ( .C (clk), .D (new_AGEMA_signal_2779), .Q (new_AGEMA_signal_2780) ) ;
    buf_clk new_AGEMA_reg_buffer_1426 ( .C (clk), .D (new_AGEMA_signal_2785), .Q (new_AGEMA_signal_2786) ) ;
    buf_clk new_AGEMA_reg_buffer_1432 ( .C (clk), .D (new_AGEMA_signal_2791), .Q (new_AGEMA_signal_2792) ) ;
    buf_clk new_AGEMA_reg_buffer_1438 ( .C (clk), .D (new_AGEMA_signal_2797), .Q (new_AGEMA_signal_2798) ) ;
    buf_clk new_AGEMA_reg_buffer_1444 ( .C (clk), .D (new_AGEMA_signal_2803), .Q (new_AGEMA_signal_2804) ) ;
    buf_clk new_AGEMA_reg_buffer_1450 ( .C (clk), .D (new_AGEMA_signal_2809), .Q (new_AGEMA_signal_2810) ) ;
    buf_clk new_AGEMA_reg_buffer_1456 ( .C (clk), .D (new_AGEMA_signal_2815), .Q (new_AGEMA_signal_2816) ) ;
    buf_clk new_AGEMA_reg_buffer_1462 ( .C (clk), .D (new_AGEMA_signal_2821), .Q (new_AGEMA_signal_2822) ) ;
    buf_clk new_AGEMA_reg_buffer_1468 ( .C (clk), .D (new_AGEMA_signal_2827), .Q (new_AGEMA_signal_2828) ) ;
    buf_clk new_AGEMA_reg_buffer_1474 ( .C (clk), .D (new_AGEMA_signal_2833), .Q (new_AGEMA_signal_2834) ) ;
    buf_clk new_AGEMA_reg_buffer_1480 ( .C (clk), .D (new_AGEMA_signal_2839), .Q (new_AGEMA_signal_2840) ) ;
    buf_clk new_AGEMA_reg_buffer_1486 ( .C (clk), .D (new_AGEMA_signal_2845), .Q (new_AGEMA_signal_2846) ) ;
    buf_clk new_AGEMA_reg_buffer_1492 ( .C (clk), .D (new_AGEMA_signal_2851), .Q (new_AGEMA_signal_2852) ) ;
    buf_clk new_AGEMA_reg_buffer_1498 ( .C (clk), .D (new_AGEMA_signal_2857), .Q (new_AGEMA_signal_2858) ) ;
    buf_clk new_AGEMA_reg_buffer_1504 ( .C (clk), .D (new_AGEMA_signal_2863), .Q (new_AGEMA_signal_2864) ) ;
    buf_clk new_AGEMA_reg_buffer_1510 ( .C (clk), .D (new_AGEMA_signal_2869), .Q (new_AGEMA_signal_2870) ) ;
    buf_clk new_AGEMA_reg_buffer_1516 ( .C (clk), .D (new_AGEMA_signal_2875), .Q (new_AGEMA_signal_2876) ) ;
    buf_clk new_AGEMA_reg_buffer_1522 ( .C (clk), .D (new_AGEMA_signal_2881), .Q (new_AGEMA_signal_2882) ) ;
    buf_clk new_AGEMA_reg_buffer_1528 ( .C (clk), .D (new_AGEMA_signal_2887), .Q (new_AGEMA_signal_2888) ) ;
    buf_clk new_AGEMA_reg_buffer_1534 ( .C (clk), .D (new_AGEMA_signal_2893), .Q (new_AGEMA_signal_2894) ) ;
    buf_clk new_AGEMA_reg_buffer_1540 ( .C (clk), .D (new_AGEMA_signal_2899), .Q (new_AGEMA_signal_2900) ) ;
    buf_clk new_AGEMA_reg_buffer_1546 ( .C (clk), .D (new_AGEMA_signal_2905), .Q (new_AGEMA_signal_2906) ) ;
    buf_clk new_AGEMA_reg_buffer_1552 ( .C (clk), .D (new_AGEMA_signal_2911), .Q (new_AGEMA_signal_2912) ) ;
    buf_clk new_AGEMA_reg_buffer_1558 ( .C (clk), .D (new_AGEMA_signal_2917), .Q (new_AGEMA_signal_2918) ) ;
    buf_clk new_AGEMA_reg_buffer_1564 ( .C (clk), .D (new_AGEMA_signal_2923), .Q (new_AGEMA_signal_2924) ) ;
    buf_clk new_AGEMA_reg_buffer_1570 ( .C (clk), .D (new_AGEMA_signal_2929), .Q (new_AGEMA_signal_2930) ) ;
    buf_clk new_AGEMA_reg_buffer_1576 ( .C (clk), .D (new_AGEMA_signal_2935), .Q (new_AGEMA_signal_2936) ) ;
    buf_clk new_AGEMA_reg_buffer_1582 ( .C (clk), .D (new_AGEMA_signal_2941), .Q (new_AGEMA_signal_2942) ) ;
    buf_clk new_AGEMA_reg_buffer_1588 ( .C (clk), .D (new_AGEMA_signal_2947), .Q (new_AGEMA_signal_2948) ) ;
    buf_clk new_AGEMA_reg_buffer_1594 ( .C (clk), .D (new_AGEMA_signal_2953), .Q (new_AGEMA_signal_2954) ) ;
    buf_clk new_AGEMA_reg_buffer_1600 ( .C (clk), .D (new_AGEMA_signal_2959), .Q (new_AGEMA_signal_2960) ) ;
    buf_clk new_AGEMA_reg_buffer_1606 ( .C (clk), .D (new_AGEMA_signal_2965), .Q (new_AGEMA_signal_2966) ) ;
    buf_clk new_AGEMA_reg_buffer_1612 ( .C (clk), .D (new_AGEMA_signal_2971), .Q (new_AGEMA_signal_2972) ) ;
    buf_clk new_AGEMA_reg_buffer_1618 ( .C (clk), .D (new_AGEMA_signal_2977), .Q (new_AGEMA_signal_2978) ) ;
    buf_clk new_AGEMA_reg_buffer_1624 ( .C (clk), .D (new_AGEMA_signal_2983), .Q (new_AGEMA_signal_2984) ) ;
    buf_clk new_AGEMA_reg_buffer_1630 ( .C (clk), .D (new_AGEMA_signal_2989), .Q (new_AGEMA_signal_2990) ) ;
    buf_clk new_AGEMA_reg_buffer_1636 ( .C (clk), .D (new_AGEMA_signal_2995), .Q (new_AGEMA_signal_2996) ) ;
    buf_clk new_AGEMA_reg_buffer_1642 ( .C (clk), .D (new_AGEMA_signal_3001), .Q (new_AGEMA_signal_3002) ) ;
    buf_clk new_AGEMA_reg_buffer_1648 ( .C (clk), .D (new_AGEMA_signal_3007), .Q (new_AGEMA_signal_3008) ) ;
    buf_clk new_AGEMA_reg_buffer_1654 ( .C (clk), .D (new_AGEMA_signal_3013), .Q (new_AGEMA_signal_3014) ) ;
    buf_clk new_AGEMA_reg_buffer_1660 ( .C (clk), .D (new_AGEMA_signal_3019), .Q (new_AGEMA_signal_3020) ) ;
    buf_clk new_AGEMA_reg_buffer_1666 ( .C (clk), .D (new_AGEMA_signal_3025), .Q (new_AGEMA_signal_3026) ) ;
    buf_clk new_AGEMA_reg_buffer_1672 ( .C (clk), .D (new_AGEMA_signal_3031), .Q (new_AGEMA_signal_3032) ) ;
    buf_clk new_AGEMA_reg_buffer_1678 ( .C (clk), .D (new_AGEMA_signal_3037), .Q (new_AGEMA_signal_3038) ) ;
    buf_clk new_AGEMA_reg_buffer_1684 ( .C (clk), .D (new_AGEMA_signal_3043), .Q (new_AGEMA_signal_3044) ) ;
    buf_clk new_AGEMA_reg_buffer_1690 ( .C (clk), .D (new_AGEMA_signal_3049), .Q (new_AGEMA_signal_3050) ) ;
    buf_clk new_AGEMA_reg_buffer_1696 ( .C (clk), .D (new_AGEMA_signal_3055), .Q (new_AGEMA_signal_3056) ) ;
    buf_clk new_AGEMA_reg_buffer_1702 ( .C (clk), .D (new_AGEMA_signal_3061), .Q (new_AGEMA_signal_3062) ) ;
    buf_clk new_AGEMA_reg_buffer_1708 ( .C (clk), .D (new_AGEMA_signal_3067), .Q (new_AGEMA_signal_3068) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C (clk), .D (new_AGEMA_signal_3073), .Q (new_AGEMA_signal_3074) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C (clk), .D (new_AGEMA_signal_3079), .Q (new_AGEMA_signal_3080) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C (clk), .D (new_AGEMA_signal_3085), .Q (new_AGEMA_signal_3086) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C (clk), .D (new_AGEMA_signal_3091), .Q (new_AGEMA_signal_3092) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C (clk), .D (new_AGEMA_signal_3097), .Q (new_AGEMA_signal_3098) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C (clk), .D (new_AGEMA_signal_3103), .Q (new_AGEMA_signal_3104) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C (clk), .D (new_AGEMA_signal_3109), .Q (new_AGEMA_signal_3110) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C (clk), .D (new_AGEMA_signal_3115), .Q (new_AGEMA_signal_3116) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C (clk), .D (new_AGEMA_signal_3121), .Q (new_AGEMA_signal_3122) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C (clk), .D (new_AGEMA_signal_3127), .Q (new_AGEMA_signal_3128) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C (clk), .D (new_AGEMA_signal_3133), .Q (new_AGEMA_signal_3134) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C (clk), .D (new_AGEMA_signal_3139), .Q (new_AGEMA_signal_3140) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C (clk), .D (new_AGEMA_signal_3145), .Q (new_AGEMA_signal_3146) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C (clk), .D (new_AGEMA_signal_3151), .Q (new_AGEMA_signal_3152) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C (clk), .D (new_AGEMA_signal_3157), .Q (new_AGEMA_signal_3158) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C (clk), .D (new_AGEMA_signal_3163), .Q (new_AGEMA_signal_3164) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C (clk), .D (new_AGEMA_signal_3169), .Q (new_AGEMA_signal_3170) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C (clk), .D (new_AGEMA_signal_3175), .Q (new_AGEMA_signal_3176) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C (clk), .D (new_AGEMA_signal_3181), .Q (new_AGEMA_signal_3182) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C (clk), .D (new_AGEMA_signal_3187), .Q (new_AGEMA_signal_3188) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C (clk), .D (new_AGEMA_signal_3193), .Q (new_AGEMA_signal_3194) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C (clk), .D (new_AGEMA_signal_3199), .Q (new_AGEMA_signal_3200) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C (clk), .D (new_AGEMA_signal_3205), .Q (new_AGEMA_signal_3206) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C (clk), .D (new_AGEMA_signal_3209), .Q (new_AGEMA_signal_3210) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C (clk), .D (new_AGEMA_signal_3211), .Q (new_AGEMA_signal_3212) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C (clk), .D (new_AGEMA_signal_3213), .Q (new_AGEMA_signal_3214) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C (clk), .D (new_AGEMA_signal_3215), .Q (new_AGEMA_signal_3216) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C (clk), .D (new_AGEMA_signal_3217), .Q (new_AGEMA_signal_3218) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C (clk), .D (new_AGEMA_signal_3219), .Q (new_AGEMA_signal_3220) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C (clk), .D (new_AGEMA_signal_3221), .Q (new_AGEMA_signal_3222) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C (clk), .D (new_AGEMA_signal_3223), .Q (new_AGEMA_signal_3224) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C (clk), .D (new_AGEMA_signal_3225), .Q (new_AGEMA_signal_3226) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C (clk), .D (new_AGEMA_signal_3227), .Q (new_AGEMA_signal_3228) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C (clk), .D (new_AGEMA_signal_3229), .Q (new_AGEMA_signal_3230) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C (clk), .D (new_AGEMA_signal_3231), .Q (new_AGEMA_signal_3232) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C (clk), .D (new_AGEMA_signal_3233), .Q (new_AGEMA_signal_3234) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C (clk), .D (new_AGEMA_signal_3235), .Q (new_AGEMA_signal_3236) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C (clk), .D (new_AGEMA_signal_3237), .Q (new_AGEMA_signal_3238) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C (clk), .D (new_AGEMA_signal_3239), .Q (new_AGEMA_signal_3240) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C (clk), .D (new_AGEMA_signal_3241), .Q (new_AGEMA_signal_3242) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C (clk), .D (new_AGEMA_signal_3243), .Q (new_AGEMA_signal_3244) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C (clk), .D (new_AGEMA_signal_3245), .Q (new_AGEMA_signal_3246) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C (clk), .D (new_AGEMA_signal_3247), .Q (new_AGEMA_signal_3248) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C (clk), .D (new_AGEMA_signal_3249), .Q (new_AGEMA_signal_3250) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C (clk), .D (new_AGEMA_signal_3251), .Q (new_AGEMA_signal_3252) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C (clk), .D (new_AGEMA_signal_3253), .Q (new_AGEMA_signal_3254) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C (clk), .D (new_AGEMA_signal_3255), .Q (new_AGEMA_signal_3256) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C (clk), .D (new_AGEMA_signal_3257), .Q (new_AGEMA_signal_3258) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C (clk), .D (new_AGEMA_signal_3259), .Q (new_AGEMA_signal_3260) ) ;
    buf_clk new_AGEMA_reg_buffer_1902 ( .C (clk), .D (new_AGEMA_signal_3261), .Q (new_AGEMA_signal_3262) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C (clk), .D (new_AGEMA_signal_3263), .Q (new_AGEMA_signal_3264) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C (clk), .D (new_AGEMA_signal_3265), .Q (new_AGEMA_signal_3266) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C (clk), .D (new_AGEMA_signal_3267), .Q (new_AGEMA_signal_3268) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C (clk), .D (new_AGEMA_signal_3269), .Q (new_AGEMA_signal_3270) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C (clk), .D (new_AGEMA_signal_3271), .Q (new_AGEMA_signal_3272) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C (clk), .D (new_AGEMA_signal_3273), .Q (new_AGEMA_signal_3274) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C (clk), .D (new_AGEMA_signal_3275), .Q (new_AGEMA_signal_3276) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C (clk), .D (new_AGEMA_signal_3277), .Q (new_AGEMA_signal_3278) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C (clk), .D (new_AGEMA_signal_3279), .Q (new_AGEMA_signal_3280) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C (clk), .D (new_AGEMA_signal_3281), .Q (new_AGEMA_signal_3282) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C (clk), .D (new_AGEMA_signal_3283), .Q (new_AGEMA_signal_3284) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C (clk), .D (new_AGEMA_signal_3285), .Q (new_AGEMA_signal_3286) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C (clk), .D (new_AGEMA_signal_3287), .Q (new_AGEMA_signal_3288) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C (clk), .D (new_AGEMA_signal_3289), .Q (new_AGEMA_signal_3290) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C (clk), .D (new_AGEMA_signal_3291), .Q (new_AGEMA_signal_3292) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C (clk), .D (new_AGEMA_signal_3293), .Q (new_AGEMA_signal_3294) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C (clk), .D (new_AGEMA_signal_3295), .Q (new_AGEMA_signal_3296) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C (clk), .D (new_AGEMA_signal_3297), .Q (new_AGEMA_signal_3298) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C (clk), .D (new_AGEMA_signal_3299), .Q (new_AGEMA_signal_3300) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C (clk), .D (new_AGEMA_signal_3301), .Q (new_AGEMA_signal_3302) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C (clk), .D (new_AGEMA_signal_3303), .Q (new_AGEMA_signal_3304) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C (clk), .D (new_AGEMA_signal_3305), .Q (new_AGEMA_signal_3306) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C (clk), .D (new_AGEMA_signal_3307), .Q (new_AGEMA_signal_3308) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C (clk), .D (new_AGEMA_signal_3309), .Q (new_AGEMA_signal_3310) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C (clk), .D (new_AGEMA_signal_3311), .Q (new_AGEMA_signal_3312) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C (clk), .D (new_AGEMA_signal_3313), .Q (new_AGEMA_signal_3314) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C (clk), .D (new_AGEMA_signal_3315), .Q (new_AGEMA_signal_3316) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C (clk), .D (new_AGEMA_signal_3317), .Q (new_AGEMA_signal_3318) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C (clk), .D (new_AGEMA_signal_3319), .Q (new_AGEMA_signal_3320) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C (clk), .D (new_AGEMA_signal_3321), .Q (new_AGEMA_signal_3322) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C (clk), .D (new_AGEMA_signal_3323), .Q (new_AGEMA_signal_3324) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C (clk), .D (new_AGEMA_signal_3325), .Q (new_AGEMA_signal_3326) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C (clk), .D (new_AGEMA_signal_3327), .Q (new_AGEMA_signal_3328) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C (clk), .D (new_AGEMA_signal_3329), .Q (new_AGEMA_signal_3330) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C (clk), .D (new_AGEMA_signal_3331), .Q (new_AGEMA_signal_3332) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C (clk), .D (new_AGEMA_signal_3333), .Q (new_AGEMA_signal_3334) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C (clk), .D (new_AGEMA_signal_3335), .Q (new_AGEMA_signal_3336) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C (clk), .D (new_AGEMA_signal_3337), .Q (new_AGEMA_signal_3338) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C (clk), .D (new_AGEMA_signal_3339), .Q (new_AGEMA_signal_3340) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C (clk), .D (new_AGEMA_signal_3341), .Q (new_AGEMA_signal_3342) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C (clk), .D (new_AGEMA_signal_3343), .Q (new_AGEMA_signal_3344) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C (clk), .D (new_AGEMA_signal_3345), .Q (new_AGEMA_signal_3346) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C (clk), .D (new_AGEMA_signal_3347), .Q (new_AGEMA_signal_3348) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C (clk), .D (new_AGEMA_signal_3349), .Q (new_AGEMA_signal_3350) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C (clk), .D (new_AGEMA_signal_3351), .Q (new_AGEMA_signal_3352) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C (clk), .D (new_AGEMA_signal_3353), .Q (new_AGEMA_signal_3354) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C (clk), .D (new_AGEMA_signal_3355), .Q (new_AGEMA_signal_3356) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C (clk), .D (new_AGEMA_signal_3357), .Q (new_AGEMA_signal_3358) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C (clk), .D (new_AGEMA_signal_3359), .Q (new_AGEMA_signal_3360) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C (clk), .D (new_AGEMA_signal_3361), .Q (new_AGEMA_signal_3362) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C (clk), .D (new_AGEMA_signal_3363), .Q (new_AGEMA_signal_3364) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C (clk), .D (new_AGEMA_signal_3365), .Q (new_AGEMA_signal_3366) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C (clk), .D (new_AGEMA_signal_3367), .Q (new_AGEMA_signal_3368) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C (clk), .D (new_AGEMA_signal_3369), .Q (new_AGEMA_signal_3370) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C (clk), .D (new_AGEMA_signal_3371), .Q (new_AGEMA_signal_3372) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C (clk), .D (new_AGEMA_signal_3373), .Q (new_AGEMA_signal_3374) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C (clk), .D (new_AGEMA_signal_3375), .Q (new_AGEMA_signal_3376) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C (clk), .D (new_AGEMA_signal_3377), .Q (new_AGEMA_signal_3378) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C (clk), .D (new_AGEMA_signal_3379), .Q (new_AGEMA_signal_3380) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C (clk), .D (new_AGEMA_signal_3381), .Q (new_AGEMA_signal_3382) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C (clk), .D (new_AGEMA_signal_3383), .Q (new_AGEMA_signal_3384) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C (clk), .D (new_AGEMA_signal_3385), .Q (new_AGEMA_signal_3386) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C (clk), .D (new_AGEMA_signal_3387), .Q (new_AGEMA_signal_3388) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C (clk), .D (new_AGEMA_signal_3389), .Q (new_AGEMA_signal_3390) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C (clk), .D (new_AGEMA_signal_3391), .Q (new_AGEMA_signal_3392) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C (clk), .D (new_AGEMA_signal_3393), .Q (new_AGEMA_signal_3394) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C (clk), .D (new_AGEMA_signal_3395), .Q (new_AGEMA_signal_3396) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C (clk), .D (new_AGEMA_signal_3397), .Q (new_AGEMA_signal_3398) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C (clk), .D (new_AGEMA_signal_3399), .Q (new_AGEMA_signal_3400) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C (clk), .D (new_AGEMA_signal_3405), .Q (new_AGEMA_signal_3406) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C (clk), .D (new_AGEMA_signal_3413), .Q (new_AGEMA_signal_3414) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C (clk), .D (new_AGEMA_signal_3421), .Q (new_AGEMA_signal_3422) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C (clk), .D (new_AGEMA_signal_3429), .Q (new_AGEMA_signal_3430) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C (clk), .D (new_AGEMA_signal_3437), .Q (new_AGEMA_signal_3438) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C (clk), .D (new_AGEMA_signal_3445), .Q (new_AGEMA_signal_3446) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C (clk), .D (new_AGEMA_signal_3453), .Q (new_AGEMA_signal_3454) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C (clk), .D (new_AGEMA_signal_3461), .Q (new_AGEMA_signal_3462) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C (clk), .D (new_AGEMA_signal_3469), .Q (new_AGEMA_signal_3470) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C (clk), .D (new_AGEMA_signal_3477), .Q (new_AGEMA_signal_3478) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C (clk), .D (new_AGEMA_signal_3485), .Q (new_AGEMA_signal_3486) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C (clk), .D (new_AGEMA_signal_3493), .Q (new_AGEMA_signal_3494) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C (clk), .D (new_AGEMA_signal_3501), .Q (new_AGEMA_signal_3502) ) ;
    buf_clk new_AGEMA_reg_buffer_2150 ( .C (clk), .D (new_AGEMA_signal_3509), .Q (new_AGEMA_signal_3510) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C (clk), .D (new_AGEMA_signal_3517), .Q (new_AGEMA_signal_3518) ) ;
    buf_clk new_AGEMA_reg_buffer_2166 ( .C (clk), .D (new_AGEMA_signal_3525), .Q (new_AGEMA_signal_3526) ) ;
    buf_clk new_AGEMA_reg_buffer_2174 ( .C (clk), .D (new_AGEMA_signal_3533), .Q (new_AGEMA_signal_3534) ) ;
    buf_clk new_AGEMA_reg_buffer_2182 ( .C (clk), .D (new_AGEMA_signal_3541), .Q (new_AGEMA_signal_3542) ) ;
    buf_clk new_AGEMA_reg_buffer_2190 ( .C (clk), .D (new_AGEMA_signal_3549), .Q (new_AGEMA_signal_3550) ) ;
    buf_clk new_AGEMA_reg_buffer_2198 ( .C (clk), .D (new_AGEMA_signal_3557), .Q (new_AGEMA_signal_3558) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C (clk), .D (new_AGEMA_signal_3565), .Q (new_AGEMA_signal_3566) ) ;
    buf_clk new_AGEMA_reg_buffer_2214 ( .C (clk), .D (new_AGEMA_signal_3573), .Q (new_AGEMA_signal_3574) ) ;
    buf_clk new_AGEMA_reg_buffer_2222 ( .C (clk), .D (new_AGEMA_signal_3581), .Q (new_AGEMA_signal_3582) ) ;
    buf_clk new_AGEMA_reg_buffer_2230 ( .C (clk), .D (new_AGEMA_signal_3589), .Q (new_AGEMA_signal_3590) ) ;
    buf_clk new_AGEMA_reg_buffer_2238 ( .C (clk), .D (new_AGEMA_signal_3597), .Q (new_AGEMA_signal_3598) ) ;
    buf_clk new_AGEMA_reg_buffer_2246 ( .C (clk), .D (new_AGEMA_signal_3605), .Q (new_AGEMA_signal_3606) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C (clk), .D (new_AGEMA_signal_3613), .Q (new_AGEMA_signal_3614) ) ;
    buf_clk new_AGEMA_reg_buffer_2262 ( .C (clk), .D (new_AGEMA_signal_3621), .Q (new_AGEMA_signal_3622) ) ;
    buf_clk new_AGEMA_reg_buffer_2270 ( .C (clk), .D (new_AGEMA_signal_3629), .Q (new_AGEMA_signal_3630) ) ;
    buf_clk new_AGEMA_reg_buffer_2278 ( .C (clk), .D (new_AGEMA_signal_3637), .Q (new_AGEMA_signal_3638) ) ;
    buf_clk new_AGEMA_reg_buffer_2286 ( .C (clk), .D (new_AGEMA_signal_3645), .Q (new_AGEMA_signal_3646) ) ;
    buf_clk new_AGEMA_reg_buffer_2294 ( .C (clk), .D (new_AGEMA_signal_3653), .Q (new_AGEMA_signal_3654) ) ;
    buf_clk new_AGEMA_reg_buffer_2302 ( .C (clk), .D (new_AGEMA_signal_3661), .Q (new_AGEMA_signal_3662) ) ;
    buf_clk new_AGEMA_reg_buffer_2310 ( .C (clk), .D (new_AGEMA_signal_3669), .Q (new_AGEMA_signal_3670) ) ;
    buf_clk new_AGEMA_reg_buffer_2318 ( .C (clk), .D (new_AGEMA_signal_3677), .Q (new_AGEMA_signal_3678) ) ;
    buf_clk new_AGEMA_reg_buffer_2326 ( .C (clk), .D (new_AGEMA_signal_3685), .Q (new_AGEMA_signal_3686) ) ;
    buf_clk new_AGEMA_reg_buffer_2334 ( .C (clk), .D (new_AGEMA_signal_3693), .Q (new_AGEMA_signal_3694) ) ;
    buf_clk new_AGEMA_reg_buffer_2342 ( .C (clk), .D (new_AGEMA_signal_3701), .Q (new_AGEMA_signal_3702) ) ;
    buf_clk new_AGEMA_reg_buffer_2350 ( .C (clk), .D (new_AGEMA_signal_3709), .Q (new_AGEMA_signal_3710) ) ;
    buf_clk new_AGEMA_reg_buffer_2358 ( .C (clk), .D (new_AGEMA_signal_3717), .Q (new_AGEMA_signal_3718) ) ;
    buf_clk new_AGEMA_reg_buffer_2366 ( .C (clk), .D (new_AGEMA_signal_3725), .Q (new_AGEMA_signal_3726) ) ;
    buf_clk new_AGEMA_reg_buffer_2374 ( .C (clk), .D (new_AGEMA_signal_3733), .Q (new_AGEMA_signal_3734) ) ;
    buf_clk new_AGEMA_reg_buffer_2382 ( .C (clk), .D (new_AGEMA_signal_3741), .Q (new_AGEMA_signal_3742) ) ;
    buf_clk new_AGEMA_reg_buffer_2390 ( .C (clk), .D (new_AGEMA_signal_3749), .Q (new_AGEMA_signal_3750) ) ;
    buf_clk new_AGEMA_reg_buffer_2398 ( .C (clk), .D (new_AGEMA_signal_3757), .Q (new_AGEMA_signal_3758) ) ;
    buf_clk new_AGEMA_reg_buffer_2406 ( .C (clk), .D (new_AGEMA_signal_3765), .Q (new_AGEMA_signal_3766) ) ;
    buf_clk new_AGEMA_reg_buffer_2414 ( .C (clk), .D (new_AGEMA_signal_3773), .Q (new_AGEMA_signal_3774) ) ;
    buf_clk new_AGEMA_reg_buffer_2422 ( .C (clk), .D (new_AGEMA_signal_3781), .Q (new_AGEMA_signal_3782) ) ;
    buf_clk new_AGEMA_reg_buffer_2430 ( .C (clk), .D (new_AGEMA_signal_3789), .Q (new_AGEMA_signal_3790) ) ;
    buf_clk new_AGEMA_reg_buffer_2438 ( .C (clk), .D (new_AGEMA_signal_3797), .Q (new_AGEMA_signal_3798) ) ;
    buf_clk new_AGEMA_reg_buffer_2446 ( .C (clk), .D (new_AGEMA_signal_3805), .Q (new_AGEMA_signal_3806) ) ;
    buf_clk new_AGEMA_reg_buffer_2454 ( .C (clk), .D (new_AGEMA_signal_3813), .Q (new_AGEMA_signal_3814) ) ;
    buf_clk new_AGEMA_reg_buffer_2462 ( .C (clk), .D (new_AGEMA_signal_3821), .Q (new_AGEMA_signal_3822) ) ;
    buf_clk new_AGEMA_reg_buffer_2470 ( .C (clk), .D (new_AGEMA_signal_3829), .Q (new_AGEMA_signal_3830) ) ;
    buf_clk new_AGEMA_reg_buffer_2478 ( .C (clk), .D (new_AGEMA_signal_3837), .Q (new_AGEMA_signal_3838) ) ;
    buf_clk new_AGEMA_reg_buffer_2486 ( .C (clk), .D (new_AGEMA_signal_3845), .Q (new_AGEMA_signal_3846) ) ;
    buf_clk new_AGEMA_reg_buffer_2494 ( .C (clk), .D (new_AGEMA_signal_3853), .Q (new_AGEMA_signal_3854) ) ;
    buf_clk new_AGEMA_reg_buffer_2502 ( .C (clk), .D (new_AGEMA_signal_3861), .Q (new_AGEMA_signal_3862) ) ;
    buf_clk new_AGEMA_reg_buffer_2510 ( .C (clk), .D (new_AGEMA_signal_3869), .Q (new_AGEMA_signal_3870) ) ;
    buf_clk new_AGEMA_reg_buffer_2518 ( .C (clk), .D (new_AGEMA_signal_3877), .Q (new_AGEMA_signal_3878) ) ;
    buf_clk new_AGEMA_reg_buffer_2526 ( .C (clk), .D (new_AGEMA_signal_3885), .Q (new_AGEMA_signal_3886) ) ;
    buf_clk new_AGEMA_reg_buffer_2534 ( .C (clk), .D (new_AGEMA_signal_3893), .Q (new_AGEMA_signal_3894) ) ;
    buf_clk new_AGEMA_reg_buffer_2542 ( .C (clk), .D (new_AGEMA_signal_3901), .Q (new_AGEMA_signal_3902) ) ;
    buf_clk new_AGEMA_reg_buffer_2550 ( .C (clk), .D (new_AGEMA_signal_3909), .Q (new_AGEMA_signal_3910) ) ;
    buf_clk new_AGEMA_reg_buffer_2558 ( .C (clk), .D (new_AGEMA_signal_3917), .Q (new_AGEMA_signal_3918) ) ;
    buf_clk new_AGEMA_reg_buffer_2566 ( .C (clk), .D (new_AGEMA_signal_3925), .Q (new_AGEMA_signal_3926) ) ;
    buf_clk new_AGEMA_reg_buffer_2574 ( .C (clk), .D (new_AGEMA_signal_3933), .Q (new_AGEMA_signal_3934) ) ;
    buf_clk new_AGEMA_reg_buffer_2582 ( .C (clk), .D (new_AGEMA_signal_3941), .Q (new_AGEMA_signal_3942) ) ;
    buf_clk new_AGEMA_reg_buffer_2590 ( .C (clk), .D (new_AGEMA_signal_3949), .Q (new_AGEMA_signal_3950) ) ;
    buf_clk new_AGEMA_reg_buffer_2598 ( .C (clk), .D (new_AGEMA_signal_3957), .Q (new_AGEMA_signal_3958) ) ;
    buf_clk new_AGEMA_reg_buffer_2606 ( .C (clk), .D (new_AGEMA_signal_3965), .Q (new_AGEMA_signal_3966) ) ;
    buf_clk new_AGEMA_reg_buffer_2614 ( .C (clk), .D (new_AGEMA_signal_3973), .Q (new_AGEMA_signal_3974) ) ;
    buf_clk new_AGEMA_reg_buffer_2622 ( .C (clk), .D (new_AGEMA_signal_3981), .Q (new_AGEMA_signal_3982) ) ;
    buf_clk new_AGEMA_reg_buffer_2630 ( .C (clk), .D (new_AGEMA_signal_3989), .Q (new_AGEMA_signal_3990) ) ;
    buf_clk new_AGEMA_reg_buffer_2638 ( .C (clk), .D (new_AGEMA_signal_3997), .Q (new_AGEMA_signal_3998) ) ;
    buf_clk new_AGEMA_reg_buffer_2646 ( .C (clk), .D (new_AGEMA_signal_4005), .Q (new_AGEMA_signal_4006) ) ;
    buf_clk new_AGEMA_reg_buffer_2654 ( .C (clk), .D (new_AGEMA_signal_4013), .Q (new_AGEMA_signal_4014) ) ;
    buf_clk new_AGEMA_reg_buffer_2662 ( .C (clk), .D (new_AGEMA_signal_4021), .Q (new_AGEMA_signal_4022) ) ;
    buf_clk new_AGEMA_reg_buffer_2670 ( .C (clk), .D (new_AGEMA_signal_4029), .Q (new_AGEMA_signal_4030) ) ;
    buf_clk new_AGEMA_reg_buffer_2678 ( .C (clk), .D (new_AGEMA_signal_4037), .Q (new_AGEMA_signal_4038) ) ;
    buf_clk new_AGEMA_reg_buffer_2686 ( .C (clk), .D (new_AGEMA_signal_4045), .Q (new_AGEMA_signal_4046) ) ;
    buf_clk new_AGEMA_reg_buffer_2694 ( .C (clk), .D (new_AGEMA_signal_4053), .Q (new_AGEMA_signal_4054) ) ;
    buf_clk new_AGEMA_reg_buffer_2702 ( .C (clk), .D (new_AGEMA_signal_4061), .Q (new_AGEMA_signal_4062) ) ;
    buf_clk new_AGEMA_reg_buffer_2710 ( .C (clk), .D (new_AGEMA_signal_4069), .Q (new_AGEMA_signal_4070) ) ;
    buf_clk new_AGEMA_reg_buffer_2718 ( .C (clk), .D (new_AGEMA_signal_4077), .Q (new_AGEMA_signal_4078) ) ;
    buf_clk new_AGEMA_reg_buffer_2726 ( .C (clk), .D (new_AGEMA_signal_4085), .Q (new_AGEMA_signal_4086) ) ;
    buf_clk new_AGEMA_reg_buffer_2734 ( .C (clk), .D (new_AGEMA_signal_4093), .Q (new_AGEMA_signal_4094) ) ;
    buf_clk new_AGEMA_reg_buffer_2742 ( .C (clk), .D (new_AGEMA_signal_4101), .Q (new_AGEMA_signal_4102) ) ;
    buf_clk new_AGEMA_reg_buffer_2750 ( .C (clk), .D (new_AGEMA_signal_4109), .Q (new_AGEMA_signal_4110) ) ;
    buf_clk new_AGEMA_reg_buffer_2758 ( .C (clk), .D (new_AGEMA_signal_4117), .Q (new_AGEMA_signal_4118) ) ;
    buf_clk new_AGEMA_reg_buffer_2766 ( .C (clk), .D (new_AGEMA_signal_4125), .Q (new_AGEMA_signal_4126) ) ;
    buf_clk new_AGEMA_reg_buffer_2774 ( .C (clk), .D (new_AGEMA_signal_4133), .Q (new_AGEMA_signal_4134) ) ;
    buf_clk new_AGEMA_reg_buffer_2782 ( .C (clk), .D (new_AGEMA_signal_4141), .Q (new_AGEMA_signal_4142) ) ;
    buf_clk new_AGEMA_reg_buffer_2790 ( .C (clk), .D (new_AGEMA_signal_4149), .Q (new_AGEMA_signal_4150) ) ;
    buf_clk new_AGEMA_reg_buffer_2798 ( .C (clk), .D (new_AGEMA_signal_4157), .Q (new_AGEMA_signal_4158) ) ;
    buf_clk new_AGEMA_reg_buffer_2806 ( .C (clk), .D (new_AGEMA_signal_4165), .Q (new_AGEMA_signal_4166) ) ;
    buf_clk new_AGEMA_reg_buffer_2814 ( .C (clk), .D (new_AGEMA_signal_4173), .Q (new_AGEMA_signal_4174) ) ;
    buf_clk new_AGEMA_reg_buffer_2822 ( .C (clk), .D (new_AGEMA_signal_4181), .Q (new_AGEMA_signal_4182) ) ;
    buf_clk new_AGEMA_reg_buffer_2830 ( .C (clk), .D (new_AGEMA_signal_4189), .Q (new_AGEMA_signal_4190) ) ;
    buf_clk new_AGEMA_reg_buffer_2838 ( .C (clk), .D (new_AGEMA_signal_4197), .Q (new_AGEMA_signal_4198) ) ;
    buf_clk new_AGEMA_reg_buffer_2846 ( .C (clk), .D (new_AGEMA_signal_4205), .Q (new_AGEMA_signal_4206) ) ;
    buf_clk new_AGEMA_reg_buffer_2854 ( .C (clk), .D (new_AGEMA_signal_4213), .Q (new_AGEMA_signal_4214) ) ;
    buf_clk new_AGEMA_reg_buffer_2862 ( .C (clk), .D (new_AGEMA_signal_4221), .Q (new_AGEMA_signal_4222) ) ;
    buf_clk new_AGEMA_reg_buffer_2870 ( .C (clk), .D (new_AGEMA_signal_4229), .Q (new_AGEMA_signal_4230) ) ;
    buf_clk new_AGEMA_reg_buffer_2878 ( .C (clk), .D (new_AGEMA_signal_4237), .Q (new_AGEMA_signal_4238) ) ;
    buf_clk new_AGEMA_reg_buffer_2886 ( .C (clk), .D (new_AGEMA_signal_4245), .Q (new_AGEMA_signal_4246) ) ;
    buf_clk new_AGEMA_reg_buffer_2894 ( .C (clk), .D (new_AGEMA_signal_4253), .Q (new_AGEMA_signal_4254) ) ;
    buf_clk new_AGEMA_reg_buffer_2902 ( .C (clk), .D (new_AGEMA_signal_4261), .Q (new_AGEMA_signal_4262) ) ;
    buf_clk new_AGEMA_reg_buffer_2910 ( .C (clk), .D (new_AGEMA_signal_4269), .Q (new_AGEMA_signal_4270) ) ;
    buf_clk new_AGEMA_reg_buffer_2918 ( .C (clk), .D (new_AGEMA_signal_4277), .Q (new_AGEMA_signal_4278) ) ;
    buf_clk new_AGEMA_reg_buffer_2926 ( .C (clk), .D (new_AGEMA_signal_4285), .Q (new_AGEMA_signal_4286) ) ;
    buf_clk new_AGEMA_reg_buffer_2934 ( .C (clk), .D (new_AGEMA_signal_4293), .Q (new_AGEMA_signal_4294) ) ;
    buf_clk new_AGEMA_reg_buffer_2942 ( .C (clk), .D (new_AGEMA_signal_4301), .Q (new_AGEMA_signal_4302) ) ;
    buf_clk new_AGEMA_reg_buffer_2950 ( .C (clk), .D (new_AGEMA_signal_4309), .Q (new_AGEMA_signal_4310) ) ;
    buf_clk new_AGEMA_reg_buffer_2958 ( .C (clk), .D (new_AGEMA_signal_4317), .Q (new_AGEMA_signal_4318) ) ;
    buf_clk new_AGEMA_reg_buffer_2966 ( .C (clk), .D (new_AGEMA_signal_4325), .Q (new_AGEMA_signal_4326) ) ;
    buf_clk new_AGEMA_reg_buffer_2974 ( .C (clk), .D (new_AGEMA_signal_4333), .Q (new_AGEMA_signal_4334) ) ;
    buf_clk new_AGEMA_reg_buffer_2982 ( .C (clk), .D (new_AGEMA_signal_4341), .Q (new_AGEMA_signal_4342) ) ;
    buf_clk new_AGEMA_reg_buffer_2990 ( .C (clk), .D (new_AGEMA_signal_4349), .Q (new_AGEMA_signal_4350) ) ;
    buf_clk new_AGEMA_reg_buffer_2998 ( .C (clk), .D (new_AGEMA_signal_4357), .Q (new_AGEMA_signal_4358) ) ;
    buf_clk new_AGEMA_reg_buffer_3006 ( .C (clk), .D (new_AGEMA_signal_4365), .Q (new_AGEMA_signal_4366) ) ;
    buf_clk new_AGEMA_reg_buffer_3014 ( .C (clk), .D (new_AGEMA_signal_4373), .Q (new_AGEMA_signal_4374) ) ;
    buf_clk new_AGEMA_reg_buffer_3022 ( .C (clk), .D (new_AGEMA_signal_4381), .Q (new_AGEMA_signal_4382) ) ;
    buf_clk new_AGEMA_reg_buffer_3030 ( .C (clk), .D (new_AGEMA_signal_4389), .Q (new_AGEMA_signal_4390) ) ;
    buf_clk new_AGEMA_reg_buffer_3038 ( .C (clk), .D (new_AGEMA_signal_4397), .Q (new_AGEMA_signal_4398) ) ;
    buf_clk new_AGEMA_reg_buffer_3046 ( .C (clk), .D (new_AGEMA_signal_4405), .Q (new_AGEMA_signal_4406) ) ;
    buf_clk new_AGEMA_reg_buffer_3054 ( .C (clk), .D (new_AGEMA_signal_4413), .Q (new_AGEMA_signal_4414) ) ;
    buf_clk new_AGEMA_reg_buffer_3062 ( .C (clk), .D (new_AGEMA_signal_4421), .Q (new_AGEMA_signal_4422) ) ;
    buf_clk new_AGEMA_reg_buffer_3072 ( .C (clk), .D (new_AGEMA_signal_4431), .Q (new_AGEMA_signal_4432) ) ;
    buf_clk new_AGEMA_reg_buffer_3076 ( .C (clk), .D (new_AGEMA_signal_4435), .Q (new_AGEMA_signal_4436) ) ;
    buf_clk new_AGEMA_reg_buffer_3084 ( .C (clk), .D (new_AGEMA_signal_4443), .Q (new_AGEMA_signal_4444) ) ;
    buf_clk new_AGEMA_reg_buffer_3088 ( .C (clk), .D (new_AGEMA_signal_4447), .Q (new_AGEMA_signal_4448) ) ;
    buf_clk new_AGEMA_reg_buffer_3096 ( .C (clk), .D (new_AGEMA_signal_4455), .Q (new_AGEMA_signal_4456) ) ;
    buf_clk new_AGEMA_reg_buffer_3100 ( .C (clk), .D (new_AGEMA_signal_4459), .Q (new_AGEMA_signal_4460) ) ;
    buf_clk new_AGEMA_reg_buffer_3108 ( .C (clk), .D (new_AGEMA_signal_4467), .Q (new_AGEMA_signal_4468) ) ;
    buf_clk new_AGEMA_reg_buffer_3112 ( .C (clk), .D (new_AGEMA_signal_4471), .Q (new_AGEMA_signal_4472) ) ;
    buf_clk new_AGEMA_reg_buffer_3120 ( .C (clk), .D (new_AGEMA_signal_4479), .Q (new_AGEMA_signal_4480) ) ;
    buf_clk new_AGEMA_reg_buffer_3124 ( .C (clk), .D (new_AGEMA_signal_4483), .Q (new_AGEMA_signal_4484) ) ;
    buf_clk new_AGEMA_reg_buffer_3132 ( .C (clk), .D (new_AGEMA_signal_4491), .Q (new_AGEMA_signal_4492) ) ;
    buf_clk new_AGEMA_reg_buffer_3136 ( .C (clk), .D (new_AGEMA_signal_4495), .Q (new_AGEMA_signal_4496) ) ;
    buf_clk new_AGEMA_reg_buffer_3144 ( .C (clk), .D (new_AGEMA_signal_4503), .Q (new_AGEMA_signal_4504) ) ;
    buf_clk new_AGEMA_reg_buffer_3148 ( .C (clk), .D (new_AGEMA_signal_4507), .Q (new_AGEMA_signal_4508) ) ;
    buf_clk new_AGEMA_reg_buffer_3156 ( .C (clk), .D (new_AGEMA_signal_4515), .Q (new_AGEMA_signal_4516) ) ;
    buf_clk new_AGEMA_reg_buffer_3160 ( .C (clk), .D (new_AGEMA_signal_4519), .Q (new_AGEMA_signal_4520) ) ;
    buf_clk new_AGEMA_reg_buffer_3168 ( .C (clk), .D (new_AGEMA_signal_4527), .Q (new_AGEMA_signal_4528) ) ;
    buf_clk new_AGEMA_reg_buffer_3172 ( .C (clk), .D (new_AGEMA_signal_4531), .Q (new_AGEMA_signal_4532) ) ;
    buf_clk new_AGEMA_reg_buffer_3180 ( .C (clk), .D (new_AGEMA_signal_4539), .Q (new_AGEMA_signal_4540) ) ;
    buf_clk new_AGEMA_reg_buffer_3184 ( .C (clk), .D (new_AGEMA_signal_4543), .Q (new_AGEMA_signal_4544) ) ;
    buf_clk new_AGEMA_reg_buffer_3192 ( .C (clk), .D (new_AGEMA_signal_4551), .Q (new_AGEMA_signal_4552) ) ;
    buf_clk new_AGEMA_reg_buffer_3196 ( .C (clk), .D (new_AGEMA_signal_4555), .Q (new_AGEMA_signal_4556) ) ;
    buf_clk new_AGEMA_reg_buffer_3204 ( .C (clk), .D (new_AGEMA_signal_4563), .Q (new_AGEMA_signal_4564) ) ;
    buf_clk new_AGEMA_reg_buffer_3208 ( .C (clk), .D (new_AGEMA_signal_4567), .Q (new_AGEMA_signal_4568) ) ;
    buf_clk new_AGEMA_reg_buffer_3216 ( .C (clk), .D (new_AGEMA_signal_4575), .Q (new_AGEMA_signal_4576) ) ;
    buf_clk new_AGEMA_reg_buffer_3220 ( .C (clk), .D (new_AGEMA_signal_4579), .Q (new_AGEMA_signal_4580) ) ;
    buf_clk new_AGEMA_reg_buffer_3228 ( .C (clk), .D (new_AGEMA_signal_4587), .Q (new_AGEMA_signal_4588) ) ;
    buf_clk new_AGEMA_reg_buffer_3232 ( .C (clk), .D (new_AGEMA_signal_4591), .Q (new_AGEMA_signal_4592) ) ;
    buf_clk new_AGEMA_reg_buffer_3240 ( .C (clk), .D (new_AGEMA_signal_4599), .Q (new_AGEMA_signal_4600) ) ;
    buf_clk new_AGEMA_reg_buffer_3244 ( .C (clk), .D (new_AGEMA_signal_4603), .Q (new_AGEMA_signal_4604) ) ;
    buf_clk new_AGEMA_reg_buffer_3252 ( .C (clk), .D (new_AGEMA_signal_4611), .Q (new_AGEMA_signal_4612) ) ;
    buf_clk new_AGEMA_reg_buffer_3256 ( .C (clk), .D (new_AGEMA_signal_4615), .Q (new_AGEMA_signal_4616) ) ;
    buf_clk new_AGEMA_reg_buffer_3390 ( .C (clk), .D (new_AGEMA_signal_4749), .Q (new_AGEMA_signal_4750) ) ;
    buf_clk new_AGEMA_reg_buffer_3398 ( .C (clk), .D (new_AGEMA_signal_4757), .Q (new_AGEMA_signal_4758) ) ;
    buf_clk new_AGEMA_reg_buffer_3406 ( .C (clk), .D (new_AGEMA_signal_4765), .Q (new_AGEMA_signal_4766) ) ;
    buf_clk new_AGEMA_reg_buffer_3414 ( .C (clk), .D (new_AGEMA_signal_4773), .Q (new_AGEMA_signal_4774) ) ;
    buf_clk new_AGEMA_reg_buffer_3422 ( .C (clk), .D (new_AGEMA_signal_4781), .Q (new_AGEMA_signal_4782) ) ;
    buf_clk new_AGEMA_reg_buffer_3430 ( .C (clk), .D (new_AGEMA_signal_4789), .Q (new_AGEMA_signal_4790) ) ;
    buf_clk new_AGEMA_reg_buffer_3438 ( .C (clk), .D (new_AGEMA_signal_4797), .Q (new_AGEMA_signal_4798) ) ;
    buf_clk new_AGEMA_reg_buffer_3446 ( .C (clk), .D (new_AGEMA_signal_4805), .Q (new_AGEMA_signal_4806) ) ;
    buf_clk new_AGEMA_reg_buffer_3454 ( .C (clk), .D (new_AGEMA_signal_4813), .Q (new_AGEMA_signal_4814) ) ;
    buf_clk new_AGEMA_reg_buffer_3462 ( .C (clk), .D (new_AGEMA_signal_4821), .Q (new_AGEMA_signal_4822) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_1079 ( .C (clk), .D (new_AGEMA_signal_2438), .Q (new_AGEMA_signal_2439) ) ;
    buf_clk new_AGEMA_reg_buffer_1085 ( .C (clk), .D (new_AGEMA_signal_2444), .Q (new_AGEMA_signal_2445) ) ;
    buf_clk new_AGEMA_reg_buffer_1091 ( .C (clk), .D (new_AGEMA_signal_2450), .Q (new_AGEMA_signal_2451) ) ;
    buf_clk new_AGEMA_reg_buffer_1097 ( .C (clk), .D (new_AGEMA_signal_2456), .Q (new_AGEMA_signal_2457) ) ;
    buf_clk new_AGEMA_reg_buffer_1103 ( .C (clk), .D (new_AGEMA_signal_2462), .Q (new_AGEMA_signal_2463) ) ;
    buf_clk new_AGEMA_reg_buffer_1109 ( .C (clk), .D (new_AGEMA_signal_2468), .Q (new_AGEMA_signal_2469) ) ;
    buf_clk new_AGEMA_reg_buffer_1115 ( .C (clk), .D (new_AGEMA_signal_2474), .Q (new_AGEMA_signal_2475) ) ;
    buf_clk new_AGEMA_reg_buffer_1121 ( .C (clk), .D (new_AGEMA_signal_2480), .Q (new_AGEMA_signal_2481) ) ;
    buf_clk new_AGEMA_reg_buffer_1127 ( .C (clk), .D (new_AGEMA_signal_2486), .Q (new_AGEMA_signal_2487) ) ;
    buf_clk new_AGEMA_reg_buffer_1133 ( .C (clk), .D (new_AGEMA_signal_2492), .Q (new_AGEMA_signal_2493) ) ;
    buf_clk new_AGEMA_reg_buffer_1139 ( .C (clk), .D (new_AGEMA_signal_2498), .Q (new_AGEMA_signal_2499) ) ;
    buf_clk new_AGEMA_reg_buffer_1145 ( .C (clk), .D (new_AGEMA_signal_2504), .Q (new_AGEMA_signal_2505) ) ;
    buf_clk new_AGEMA_reg_buffer_1151 ( .C (clk), .D (new_AGEMA_signal_2510), .Q (new_AGEMA_signal_2511) ) ;
    buf_clk new_AGEMA_reg_buffer_1157 ( .C (clk), .D (new_AGEMA_signal_2516), .Q (new_AGEMA_signal_2517) ) ;
    buf_clk new_AGEMA_reg_buffer_1163 ( .C (clk), .D (new_AGEMA_signal_2522), .Q (new_AGEMA_signal_2523) ) ;
    buf_clk new_AGEMA_reg_buffer_1169 ( .C (clk), .D (new_AGEMA_signal_2528), .Q (new_AGEMA_signal_2529) ) ;
    buf_clk new_AGEMA_reg_buffer_1175 ( .C (clk), .D (new_AGEMA_signal_2534), .Q (new_AGEMA_signal_2535) ) ;
    buf_clk new_AGEMA_reg_buffer_1181 ( .C (clk), .D (new_AGEMA_signal_2540), .Q (new_AGEMA_signal_2541) ) ;
    buf_clk new_AGEMA_reg_buffer_1187 ( .C (clk), .D (new_AGEMA_signal_2546), .Q (new_AGEMA_signal_2547) ) ;
    buf_clk new_AGEMA_reg_buffer_1193 ( .C (clk), .D (new_AGEMA_signal_2552), .Q (new_AGEMA_signal_2553) ) ;
    buf_clk new_AGEMA_reg_buffer_1199 ( .C (clk), .D (new_AGEMA_signal_2558), .Q (new_AGEMA_signal_2559) ) ;
    buf_clk new_AGEMA_reg_buffer_1205 ( .C (clk), .D (new_AGEMA_signal_2564), .Q (new_AGEMA_signal_2565) ) ;
    buf_clk new_AGEMA_reg_buffer_1211 ( .C (clk), .D (new_AGEMA_signal_2570), .Q (new_AGEMA_signal_2571) ) ;
    buf_clk new_AGEMA_reg_buffer_1217 ( .C (clk), .D (new_AGEMA_signal_2576), .Q (new_AGEMA_signal_2577) ) ;
    buf_clk new_AGEMA_reg_buffer_1223 ( .C (clk), .D (new_AGEMA_signal_2582), .Q (new_AGEMA_signal_2583) ) ;
    buf_clk new_AGEMA_reg_buffer_1229 ( .C (clk), .D (new_AGEMA_signal_2588), .Q (new_AGEMA_signal_2589) ) ;
    buf_clk new_AGEMA_reg_buffer_1235 ( .C (clk), .D (new_AGEMA_signal_2594), .Q (new_AGEMA_signal_2595) ) ;
    buf_clk new_AGEMA_reg_buffer_1241 ( .C (clk), .D (new_AGEMA_signal_2600), .Q (new_AGEMA_signal_2601) ) ;
    buf_clk new_AGEMA_reg_buffer_1247 ( .C (clk), .D (new_AGEMA_signal_2606), .Q (new_AGEMA_signal_2607) ) ;
    buf_clk new_AGEMA_reg_buffer_1253 ( .C (clk), .D (new_AGEMA_signal_2612), .Q (new_AGEMA_signal_2613) ) ;
    buf_clk new_AGEMA_reg_buffer_1259 ( .C (clk), .D (new_AGEMA_signal_2618), .Q (new_AGEMA_signal_2619) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C (clk), .D (new_AGEMA_signal_2624), .Q (new_AGEMA_signal_2625) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C (clk), .D (new_AGEMA_signal_2630), .Q (new_AGEMA_signal_2631) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C (clk), .D (new_AGEMA_signal_2636), .Q (new_AGEMA_signal_2637) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C (clk), .D (new_AGEMA_signal_2642), .Q (new_AGEMA_signal_2643) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C (clk), .D (new_AGEMA_signal_2648), .Q (new_AGEMA_signal_2649) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C (clk), .D (new_AGEMA_signal_2654), .Q (new_AGEMA_signal_2655) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C (clk), .D (new_AGEMA_signal_2660), .Q (new_AGEMA_signal_2661) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C (clk), .D (new_AGEMA_signal_2666), .Q (new_AGEMA_signal_2667) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C (clk), .D (new_AGEMA_signal_2672), .Q (new_AGEMA_signal_2673) ) ;
    buf_clk new_AGEMA_reg_buffer_1319 ( .C (clk), .D (new_AGEMA_signal_2678), .Q (new_AGEMA_signal_2679) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C (clk), .D (new_AGEMA_signal_2684), .Q (new_AGEMA_signal_2685) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C (clk), .D (new_AGEMA_signal_2690), .Q (new_AGEMA_signal_2691) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C (clk), .D (new_AGEMA_signal_2696), .Q (new_AGEMA_signal_2697) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C (clk), .D (new_AGEMA_signal_2702), .Q (new_AGEMA_signal_2703) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C (clk), .D (new_AGEMA_signal_2708), .Q (new_AGEMA_signal_2709) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C (clk), .D (new_AGEMA_signal_2714), .Q (new_AGEMA_signal_2715) ) ;
    buf_clk new_AGEMA_reg_buffer_1361 ( .C (clk), .D (new_AGEMA_signal_2720), .Q (new_AGEMA_signal_2721) ) ;
    buf_clk new_AGEMA_reg_buffer_1367 ( .C (clk), .D (new_AGEMA_signal_2726), .Q (new_AGEMA_signal_2727) ) ;
    buf_clk new_AGEMA_reg_buffer_1373 ( .C (clk), .D (new_AGEMA_signal_2732), .Q (new_AGEMA_signal_2733) ) ;
    buf_clk new_AGEMA_reg_buffer_1379 ( .C (clk), .D (new_AGEMA_signal_2738), .Q (new_AGEMA_signal_2739) ) ;
    buf_clk new_AGEMA_reg_buffer_1385 ( .C (clk), .D (new_AGEMA_signal_2744), .Q (new_AGEMA_signal_2745) ) ;
    buf_clk new_AGEMA_reg_buffer_1391 ( .C (clk), .D (new_AGEMA_signal_2750), .Q (new_AGEMA_signal_2751) ) ;
    buf_clk new_AGEMA_reg_buffer_1397 ( .C (clk), .D (new_AGEMA_signal_2756), .Q (new_AGEMA_signal_2757) ) ;
    buf_clk new_AGEMA_reg_buffer_1403 ( .C (clk), .D (new_AGEMA_signal_2762), .Q (new_AGEMA_signal_2763) ) ;
    buf_clk new_AGEMA_reg_buffer_1409 ( .C (clk), .D (new_AGEMA_signal_2768), .Q (new_AGEMA_signal_2769) ) ;
    buf_clk new_AGEMA_reg_buffer_1415 ( .C (clk), .D (new_AGEMA_signal_2774), .Q (new_AGEMA_signal_2775) ) ;
    buf_clk new_AGEMA_reg_buffer_1421 ( .C (clk), .D (new_AGEMA_signal_2780), .Q (new_AGEMA_signal_2781) ) ;
    buf_clk new_AGEMA_reg_buffer_1427 ( .C (clk), .D (new_AGEMA_signal_2786), .Q (new_AGEMA_signal_2787) ) ;
    buf_clk new_AGEMA_reg_buffer_1433 ( .C (clk), .D (new_AGEMA_signal_2792), .Q (new_AGEMA_signal_2793) ) ;
    buf_clk new_AGEMA_reg_buffer_1439 ( .C (clk), .D (new_AGEMA_signal_2798), .Q (new_AGEMA_signal_2799) ) ;
    buf_clk new_AGEMA_reg_buffer_1445 ( .C (clk), .D (new_AGEMA_signal_2804), .Q (new_AGEMA_signal_2805) ) ;
    buf_clk new_AGEMA_reg_buffer_1451 ( .C (clk), .D (new_AGEMA_signal_2810), .Q (new_AGEMA_signal_2811) ) ;
    buf_clk new_AGEMA_reg_buffer_1457 ( .C (clk), .D (new_AGEMA_signal_2816), .Q (new_AGEMA_signal_2817) ) ;
    buf_clk new_AGEMA_reg_buffer_1463 ( .C (clk), .D (new_AGEMA_signal_2822), .Q (new_AGEMA_signal_2823) ) ;
    buf_clk new_AGEMA_reg_buffer_1469 ( .C (clk), .D (new_AGEMA_signal_2828), .Q (new_AGEMA_signal_2829) ) ;
    buf_clk new_AGEMA_reg_buffer_1475 ( .C (clk), .D (new_AGEMA_signal_2834), .Q (new_AGEMA_signal_2835) ) ;
    buf_clk new_AGEMA_reg_buffer_1481 ( .C (clk), .D (new_AGEMA_signal_2840), .Q (new_AGEMA_signal_2841) ) ;
    buf_clk new_AGEMA_reg_buffer_1487 ( .C (clk), .D (new_AGEMA_signal_2846), .Q (new_AGEMA_signal_2847) ) ;
    buf_clk new_AGEMA_reg_buffer_1493 ( .C (clk), .D (new_AGEMA_signal_2852), .Q (new_AGEMA_signal_2853) ) ;
    buf_clk new_AGEMA_reg_buffer_1499 ( .C (clk), .D (new_AGEMA_signal_2858), .Q (new_AGEMA_signal_2859) ) ;
    buf_clk new_AGEMA_reg_buffer_1505 ( .C (clk), .D (new_AGEMA_signal_2864), .Q (new_AGEMA_signal_2865) ) ;
    buf_clk new_AGEMA_reg_buffer_1511 ( .C (clk), .D (new_AGEMA_signal_2870), .Q (new_AGEMA_signal_2871) ) ;
    buf_clk new_AGEMA_reg_buffer_1517 ( .C (clk), .D (new_AGEMA_signal_2876), .Q (new_AGEMA_signal_2877) ) ;
    buf_clk new_AGEMA_reg_buffer_1523 ( .C (clk), .D (new_AGEMA_signal_2882), .Q (new_AGEMA_signal_2883) ) ;
    buf_clk new_AGEMA_reg_buffer_1529 ( .C (clk), .D (new_AGEMA_signal_2888), .Q (new_AGEMA_signal_2889) ) ;
    buf_clk new_AGEMA_reg_buffer_1535 ( .C (clk), .D (new_AGEMA_signal_2894), .Q (new_AGEMA_signal_2895) ) ;
    buf_clk new_AGEMA_reg_buffer_1541 ( .C (clk), .D (new_AGEMA_signal_2900), .Q (new_AGEMA_signal_2901) ) ;
    buf_clk new_AGEMA_reg_buffer_1547 ( .C (clk), .D (new_AGEMA_signal_2906), .Q (new_AGEMA_signal_2907) ) ;
    buf_clk new_AGEMA_reg_buffer_1553 ( .C (clk), .D (new_AGEMA_signal_2912), .Q (new_AGEMA_signal_2913) ) ;
    buf_clk new_AGEMA_reg_buffer_1559 ( .C (clk), .D (new_AGEMA_signal_2918), .Q (new_AGEMA_signal_2919) ) ;
    buf_clk new_AGEMA_reg_buffer_1565 ( .C (clk), .D (new_AGEMA_signal_2924), .Q (new_AGEMA_signal_2925) ) ;
    buf_clk new_AGEMA_reg_buffer_1571 ( .C (clk), .D (new_AGEMA_signal_2930), .Q (new_AGEMA_signal_2931) ) ;
    buf_clk new_AGEMA_reg_buffer_1577 ( .C (clk), .D (new_AGEMA_signal_2936), .Q (new_AGEMA_signal_2937) ) ;
    buf_clk new_AGEMA_reg_buffer_1583 ( .C (clk), .D (new_AGEMA_signal_2942), .Q (new_AGEMA_signal_2943) ) ;
    buf_clk new_AGEMA_reg_buffer_1589 ( .C (clk), .D (new_AGEMA_signal_2948), .Q (new_AGEMA_signal_2949) ) ;
    buf_clk new_AGEMA_reg_buffer_1595 ( .C (clk), .D (new_AGEMA_signal_2954), .Q (new_AGEMA_signal_2955) ) ;
    buf_clk new_AGEMA_reg_buffer_1601 ( .C (clk), .D (new_AGEMA_signal_2960), .Q (new_AGEMA_signal_2961) ) ;
    buf_clk new_AGEMA_reg_buffer_1607 ( .C (clk), .D (new_AGEMA_signal_2966), .Q (new_AGEMA_signal_2967) ) ;
    buf_clk new_AGEMA_reg_buffer_1613 ( .C (clk), .D (new_AGEMA_signal_2972), .Q (new_AGEMA_signal_2973) ) ;
    buf_clk new_AGEMA_reg_buffer_1619 ( .C (clk), .D (new_AGEMA_signal_2978), .Q (new_AGEMA_signal_2979) ) ;
    buf_clk new_AGEMA_reg_buffer_1625 ( .C (clk), .D (new_AGEMA_signal_2984), .Q (new_AGEMA_signal_2985) ) ;
    buf_clk new_AGEMA_reg_buffer_1631 ( .C (clk), .D (new_AGEMA_signal_2990), .Q (new_AGEMA_signal_2991) ) ;
    buf_clk new_AGEMA_reg_buffer_1637 ( .C (clk), .D (new_AGEMA_signal_2996), .Q (new_AGEMA_signal_2997) ) ;
    buf_clk new_AGEMA_reg_buffer_1643 ( .C (clk), .D (new_AGEMA_signal_3002), .Q (new_AGEMA_signal_3003) ) ;
    buf_clk new_AGEMA_reg_buffer_1649 ( .C (clk), .D (new_AGEMA_signal_3008), .Q (new_AGEMA_signal_3009) ) ;
    buf_clk new_AGEMA_reg_buffer_1655 ( .C (clk), .D (new_AGEMA_signal_3014), .Q (new_AGEMA_signal_3015) ) ;
    buf_clk new_AGEMA_reg_buffer_1661 ( .C (clk), .D (new_AGEMA_signal_3020), .Q (new_AGEMA_signal_3021) ) ;
    buf_clk new_AGEMA_reg_buffer_1667 ( .C (clk), .D (new_AGEMA_signal_3026), .Q (new_AGEMA_signal_3027) ) ;
    buf_clk new_AGEMA_reg_buffer_1673 ( .C (clk), .D (new_AGEMA_signal_3032), .Q (new_AGEMA_signal_3033) ) ;
    buf_clk new_AGEMA_reg_buffer_1679 ( .C (clk), .D (new_AGEMA_signal_3038), .Q (new_AGEMA_signal_3039) ) ;
    buf_clk new_AGEMA_reg_buffer_1685 ( .C (clk), .D (new_AGEMA_signal_3044), .Q (new_AGEMA_signal_3045) ) ;
    buf_clk new_AGEMA_reg_buffer_1691 ( .C (clk), .D (new_AGEMA_signal_3050), .Q (new_AGEMA_signal_3051) ) ;
    buf_clk new_AGEMA_reg_buffer_1697 ( .C (clk), .D (new_AGEMA_signal_3056), .Q (new_AGEMA_signal_3057) ) ;
    buf_clk new_AGEMA_reg_buffer_1703 ( .C (clk), .D (new_AGEMA_signal_3062), .Q (new_AGEMA_signal_3063) ) ;
    buf_clk new_AGEMA_reg_buffer_1709 ( .C (clk), .D (new_AGEMA_signal_3068), .Q (new_AGEMA_signal_3069) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C (clk), .D (new_AGEMA_signal_3074), .Q (new_AGEMA_signal_3075) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C (clk), .D (new_AGEMA_signal_3080), .Q (new_AGEMA_signal_3081) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C (clk), .D (new_AGEMA_signal_3086), .Q (new_AGEMA_signal_3087) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C (clk), .D (new_AGEMA_signal_3092), .Q (new_AGEMA_signal_3093) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C (clk), .D (new_AGEMA_signal_3098), .Q (new_AGEMA_signal_3099) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C (clk), .D (new_AGEMA_signal_3104), .Q (new_AGEMA_signal_3105) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C (clk), .D (new_AGEMA_signal_3110), .Q (new_AGEMA_signal_3111) ) ;
    buf_clk new_AGEMA_reg_buffer_1757 ( .C (clk), .D (new_AGEMA_signal_3116), .Q (new_AGEMA_signal_3117) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C (clk), .D (new_AGEMA_signal_3122), .Q (new_AGEMA_signal_3123) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C (clk), .D (new_AGEMA_signal_3128), .Q (new_AGEMA_signal_3129) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C (clk), .D (new_AGEMA_signal_3134), .Q (new_AGEMA_signal_3135) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C (clk), .D (new_AGEMA_signal_3140), .Q (new_AGEMA_signal_3141) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C (clk), .D (new_AGEMA_signal_3146), .Q (new_AGEMA_signal_3147) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C (clk), .D (new_AGEMA_signal_3152), .Q (new_AGEMA_signal_3153) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C (clk), .D (new_AGEMA_signal_3158), .Q (new_AGEMA_signal_3159) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C (clk), .D (new_AGEMA_signal_3164), .Q (new_AGEMA_signal_3165) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C (clk), .D (new_AGEMA_signal_3170), .Q (new_AGEMA_signal_3171) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C (clk), .D (new_AGEMA_signal_3176), .Q (new_AGEMA_signal_3177) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C (clk), .D (new_AGEMA_signal_3182), .Q (new_AGEMA_signal_3183) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C (clk), .D (new_AGEMA_signal_3188), .Q (new_AGEMA_signal_3189) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C (clk), .D (new_AGEMA_signal_3194), .Q (new_AGEMA_signal_3195) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C (clk), .D (new_AGEMA_signal_3200), .Q (new_AGEMA_signal_3201) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C (clk), .D (new_AGEMA_signal_3206), .Q (new_AGEMA_signal_3207) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C (clk), .D (new_AGEMA_signal_3406), .Q (new_AGEMA_signal_3407) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C (clk), .D (new_AGEMA_signal_3414), .Q (new_AGEMA_signal_3415) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C (clk), .D (new_AGEMA_signal_3422), .Q (new_AGEMA_signal_3423) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C (clk), .D (new_AGEMA_signal_3430), .Q (new_AGEMA_signal_3431) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C (clk), .D (new_AGEMA_signal_3438), .Q (new_AGEMA_signal_3439) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C (clk), .D (new_AGEMA_signal_3446), .Q (new_AGEMA_signal_3447) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C (clk), .D (new_AGEMA_signal_3454), .Q (new_AGEMA_signal_3455) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C (clk), .D (new_AGEMA_signal_3462), .Q (new_AGEMA_signal_3463) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C (clk), .D (new_AGEMA_signal_3470), .Q (new_AGEMA_signal_3471) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C (clk), .D (new_AGEMA_signal_3478), .Q (new_AGEMA_signal_3479) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C (clk), .D (new_AGEMA_signal_3486), .Q (new_AGEMA_signal_3487) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C (clk), .D (new_AGEMA_signal_3494), .Q (new_AGEMA_signal_3495) ) ;
    buf_clk new_AGEMA_reg_buffer_2143 ( .C (clk), .D (new_AGEMA_signal_3502), .Q (new_AGEMA_signal_3503) ) ;
    buf_clk new_AGEMA_reg_buffer_2151 ( .C (clk), .D (new_AGEMA_signal_3510), .Q (new_AGEMA_signal_3511) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C (clk), .D (new_AGEMA_signal_3518), .Q (new_AGEMA_signal_3519) ) ;
    buf_clk new_AGEMA_reg_buffer_2167 ( .C (clk), .D (new_AGEMA_signal_3526), .Q (new_AGEMA_signal_3527) ) ;
    buf_clk new_AGEMA_reg_buffer_2175 ( .C (clk), .D (new_AGEMA_signal_3534), .Q (new_AGEMA_signal_3535) ) ;
    buf_clk new_AGEMA_reg_buffer_2183 ( .C (clk), .D (new_AGEMA_signal_3542), .Q (new_AGEMA_signal_3543) ) ;
    buf_clk new_AGEMA_reg_buffer_2191 ( .C (clk), .D (new_AGEMA_signal_3550), .Q (new_AGEMA_signal_3551) ) ;
    buf_clk new_AGEMA_reg_buffer_2199 ( .C (clk), .D (new_AGEMA_signal_3558), .Q (new_AGEMA_signal_3559) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C (clk), .D (new_AGEMA_signal_3566), .Q (new_AGEMA_signal_3567) ) ;
    buf_clk new_AGEMA_reg_buffer_2215 ( .C (clk), .D (new_AGEMA_signal_3574), .Q (new_AGEMA_signal_3575) ) ;
    buf_clk new_AGEMA_reg_buffer_2223 ( .C (clk), .D (new_AGEMA_signal_3582), .Q (new_AGEMA_signal_3583) ) ;
    buf_clk new_AGEMA_reg_buffer_2231 ( .C (clk), .D (new_AGEMA_signal_3590), .Q (new_AGEMA_signal_3591) ) ;
    buf_clk new_AGEMA_reg_buffer_2239 ( .C (clk), .D (new_AGEMA_signal_3598), .Q (new_AGEMA_signal_3599) ) ;
    buf_clk new_AGEMA_reg_buffer_2247 ( .C (clk), .D (new_AGEMA_signal_3606), .Q (new_AGEMA_signal_3607) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C (clk), .D (new_AGEMA_signal_3614), .Q (new_AGEMA_signal_3615) ) ;
    buf_clk new_AGEMA_reg_buffer_2263 ( .C (clk), .D (new_AGEMA_signal_3622), .Q (new_AGEMA_signal_3623) ) ;
    buf_clk new_AGEMA_reg_buffer_2271 ( .C (clk), .D (new_AGEMA_signal_3630), .Q (new_AGEMA_signal_3631) ) ;
    buf_clk new_AGEMA_reg_buffer_2279 ( .C (clk), .D (new_AGEMA_signal_3638), .Q (new_AGEMA_signal_3639) ) ;
    buf_clk new_AGEMA_reg_buffer_2287 ( .C (clk), .D (new_AGEMA_signal_3646), .Q (new_AGEMA_signal_3647) ) ;
    buf_clk new_AGEMA_reg_buffer_2295 ( .C (clk), .D (new_AGEMA_signal_3654), .Q (new_AGEMA_signal_3655) ) ;
    buf_clk new_AGEMA_reg_buffer_2303 ( .C (clk), .D (new_AGEMA_signal_3662), .Q (new_AGEMA_signal_3663) ) ;
    buf_clk new_AGEMA_reg_buffer_2311 ( .C (clk), .D (new_AGEMA_signal_3670), .Q (new_AGEMA_signal_3671) ) ;
    buf_clk new_AGEMA_reg_buffer_2319 ( .C (clk), .D (new_AGEMA_signal_3678), .Q (new_AGEMA_signal_3679) ) ;
    buf_clk new_AGEMA_reg_buffer_2327 ( .C (clk), .D (new_AGEMA_signal_3686), .Q (new_AGEMA_signal_3687) ) ;
    buf_clk new_AGEMA_reg_buffer_2335 ( .C (clk), .D (new_AGEMA_signal_3694), .Q (new_AGEMA_signal_3695) ) ;
    buf_clk new_AGEMA_reg_buffer_2343 ( .C (clk), .D (new_AGEMA_signal_3702), .Q (new_AGEMA_signal_3703) ) ;
    buf_clk new_AGEMA_reg_buffer_2351 ( .C (clk), .D (new_AGEMA_signal_3710), .Q (new_AGEMA_signal_3711) ) ;
    buf_clk new_AGEMA_reg_buffer_2359 ( .C (clk), .D (new_AGEMA_signal_3718), .Q (new_AGEMA_signal_3719) ) ;
    buf_clk new_AGEMA_reg_buffer_2367 ( .C (clk), .D (new_AGEMA_signal_3726), .Q (new_AGEMA_signal_3727) ) ;
    buf_clk new_AGEMA_reg_buffer_2375 ( .C (clk), .D (new_AGEMA_signal_3734), .Q (new_AGEMA_signal_3735) ) ;
    buf_clk new_AGEMA_reg_buffer_2383 ( .C (clk), .D (new_AGEMA_signal_3742), .Q (new_AGEMA_signal_3743) ) ;
    buf_clk new_AGEMA_reg_buffer_2391 ( .C (clk), .D (new_AGEMA_signal_3750), .Q (new_AGEMA_signal_3751) ) ;
    buf_clk new_AGEMA_reg_buffer_2399 ( .C (clk), .D (new_AGEMA_signal_3758), .Q (new_AGEMA_signal_3759) ) ;
    buf_clk new_AGEMA_reg_buffer_2407 ( .C (clk), .D (new_AGEMA_signal_3766), .Q (new_AGEMA_signal_3767) ) ;
    buf_clk new_AGEMA_reg_buffer_2415 ( .C (clk), .D (new_AGEMA_signal_3774), .Q (new_AGEMA_signal_3775) ) ;
    buf_clk new_AGEMA_reg_buffer_2423 ( .C (clk), .D (new_AGEMA_signal_3782), .Q (new_AGEMA_signal_3783) ) ;
    buf_clk new_AGEMA_reg_buffer_2431 ( .C (clk), .D (new_AGEMA_signal_3790), .Q (new_AGEMA_signal_3791) ) ;
    buf_clk new_AGEMA_reg_buffer_2439 ( .C (clk), .D (new_AGEMA_signal_3798), .Q (new_AGEMA_signal_3799) ) ;
    buf_clk new_AGEMA_reg_buffer_2447 ( .C (clk), .D (new_AGEMA_signal_3806), .Q (new_AGEMA_signal_3807) ) ;
    buf_clk new_AGEMA_reg_buffer_2455 ( .C (clk), .D (new_AGEMA_signal_3814), .Q (new_AGEMA_signal_3815) ) ;
    buf_clk new_AGEMA_reg_buffer_2463 ( .C (clk), .D (new_AGEMA_signal_3822), .Q (new_AGEMA_signal_3823) ) ;
    buf_clk new_AGEMA_reg_buffer_2471 ( .C (clk), .D (new_AGEMA_signal_3830), .Q (new_AGEMA_signal_3831) ) ;
    buf_clk new_AGEMA_reg_buffer_2479 ( .C (clk), .D (new_AGEMA_signal_3838), .Q (new_AGEMA_signal_3839) ) ;
    buf_clk new_AGEMA_reg_buffer_2487 ( .C (clk), .D (new_AGEMA_signal_3846), .Q (new_AGEMA_signal_3847) ) ;
    buf_clk new_AGEMA_reg_buffer_2495 ( .C (clk), .D (new_AGEMA_signal_3854), .Q (new_AGEMA_signal_3855) ) ;
    buf_clk new_AGEMA_reg_buffer_2503 ( .C (clk), .D (new_AGEMA_signal_3862), .Q (new_AGEMA_signal_3863) ) ;
    buf_clk new_AGEMA_reg_buffer_2511 ( .C (clk), .D (new_AGEMA_signal_3870), .Q (new_AGEMA_signal_3871) ) ;
    buf_clk new_AGEMA_reg_buffer_2519 ( .C (clk), .D (new_AGEMA_signal_3878), .Q (new_AGEMA_signal_3879) ) ;
    buf_clk new_AGEMA_reg_buffer_2527 ( .C (clk), .D (new_AGEMA_signal_3886), .Q (new_AGEMA_signal_3887) ) ;
    buf_clk new_AGEMA_reg_buffer_2535 ( .C (clk), .D (new_AGEMA_signal_3894), .Q (new_AGEMA_signal_3895) ) ;
    buf_clk new_AGEMA_reg_buffer_2543 ( .C (clk), .D (new_AGEMA_signal_3902), .Q (new_AGEMA_signal_3903) ) ;
    buf_clk new_AGEMA_reg_buffer_2551 ( .C (clk), .D (new_AGEMA_signal_3910), .Q (new_AGEMA_signal_3911) ) ;
    buf_clk new_AGEMA_reg_buffer_2559 ( .C (clk), .D (new_AGEMA_signal_3918), .Q (new_AGEMA_signal_3919) ) ;
    buf_clk new_AGEMA_reg_buffer_2567 ( .C (clk), .D (new_AGEMA_signal_3926), .Q (new_AGEMA_signal_3927) ) ;
    buf_clk new_AGEMA_reg_buffer_2575 ( .C (clk), .D (new_AGEMA_signal_3934), .Q (new_AGEMA_signal_3935) ) ;
    buf_clk new_AGEMA_reg_buffer_2583 ( .C (clk), .D (new_AGEMA_signal_3942), .Q (new_AGEMA_signal_3943) ) ;
    buf_clk new_AGEMA_reg_buffer_2591 ( .C (clk), .D (new_AGEMA_signal_3950), .Q (new_AGEMA_signal_3951) ) ;
    buf_clk new_AGEMA_reg_buffer_2599 ( .C (clk), .D (new_AGEMA_signal_3958), .Q (new_AGEMA_signal_3959) ) ;
    buf_clk new_AGEMA_reg_buffer_2607 ( .C (clk), .D (new_AGEMA_signal_3966), .Q (new_AGEMA_signal_3967) ) ;
    buf_clk new_AGEMA_reg_buffer_2615 ( .C (clk), .D (new_AGEMA_signal_3974), .Q (new_AGEMA_signal_3975) ) ;
    buf_clk new_AGEMA_reg_buffer_2623 ( .C (clk), .D (new_AGEMA_signal_3982), .Q (new_AGEMA_signal_3983) ) ;
    buf_clk new_AGEMA_reg_buffer_2631 ( .C (clk), .D (new_AGEMA_signal_3990), .Q (new_AGEMA_signal_3991) ) ;
    buf_clk new_AGEMA_reg_buffer_2639 ( .C (clk), .D (new_AGEMA_signal_3998), .Q (new_AGEMA_signal_3999) ) ;
    buf_clk new_AGEMA_reg_buffer_2647 ( .C (clk), .D (new_AGEMA_signal_4006), .Q (new_AGEMA_signal_4007) ) ;
    buf_clk new_AGEMA_reg_buffer_2655 ( .C (clk), .D (new_AGEMA_signal_4014), .Q (new_AGEMA_signal_4015) ) ;
    buf_clk new_AGEMA_reg_buffer_2663 ( .C (clk), .D (new_AGEMA_signal_4022), .Q (new_AGEMA_signal_4023) ) ;
    buf_clk new_AGEMA_reg_buffer_2671 ( .C (clk), .D (new_AGEMA_signal_4030), .Q (new_AGEMA_signal_4031) ) ;
    buf_clk new_AGEMA_reg_buffer_2679 ( .C (clk), .D (new_AGEMA_signal_4038), .Q (new_AGEMA_signal_4039) ) ;
    buf_clk new_AGEMA_reg_buffer_2687 ( .C (clk), .D (new_AGEMA_signal_4046), .Q (new_AGEMA_signal_4047) ) ;
    buf_clk new_AGEMA_reg_buffer_2695 ( .C (clk), .D (new_AGEMA_signal_4054), .Q (new_AGEMA_signal_4055) ) ;
    buf_clk new_AGEMA_reg_buffer_2703 ( .C (clk), .D (new_AGEMA_signal_4062), .Q (new_AGEMA_signal_4063) ) ;
    buf_clk new_AGEMA_reg_buffer_2711 ( .C (clk), .D (new_AGEMA_signal_4070), .Q (new_AGEMA_signal_4071) ) ;
    buf_clk new_AGEMA_reg_buffer_2719 ( .C (clk), .D (new_AGEMA_signal_4078), .Q (new_AGEMA_signal_4079) ) ;
    buf_clk new_AGEMA_reg_buffer_2727 ( .C (clk), .D (new_AGEMA_signal_4086), .Q (new_AGEMA_signal_4087) ) ;
    buf_clk new_AGEMA_reg_buffer_2735 ( .C (clk), .D (new_AGEMA_signal_4094), .Q (new_AGEMA_signal_4095) ) ;
    buf_clk new_AGEMA_reg_buffer_2743 ( .C (clk), .D (new_AGEMA_signal_4102), .Q (new_AGEMA_signal_4103) ) ;
    buf_clk new_AGEMA_reg_buffer_2751 ( .C (clk), .D (new_AGEMA_signal_4110), .Q (new_AGEMA_signal_4111) ) ;
    buf_clk new_AGEMA_reg_buffer_2759 ( .C (clk), .D (new_AGEMA_signal_4118), .Q (new_AGEMA_signal_4119) ) ;
    buf_clk new_AGEMA_reg_buffer_2767 ( .C (clk), .D (new_AGEMA_signal_4126), .Q (new_AGEMA_signal_4127) ) ;
    buf_clk new_AGEMA_reg_buffer_2775 ( .C (clk), .D (new_AGEMA_signal_4134), .Q (new_AGEMA_signal_4135) ) ;
    buf_clk new_AGEMA_reg_buffer_2783 ( .C (clk), .D (new_AGEMA_signal_4142), .Q (new_AGEMA_signal_4143) ) ;
    buf_clk new_AGEMA_reg_buffer_2791 ( .C (clk), .D (new_AGEMA_signal_4150), .Q (new_AGEMA_signal_4151) ) ;
    buf_clk new_AGEMA_reg_buffer_2799 ( .C (clk), .D (new_AGEMA_signal_4158), .Q (new_AGEMA_signal_4159) ) ;
    buf_clk new_AGEMA_reg_buffer_2807 ( .C (clk), .D (new_AGEMA_signal_4166), .Q (new_AGEMA_signal_4167) ) ;
    buf_clk new_AGEMA_reg_buffer_2815 ( .C (clk), .D (new_AGEMA_signal_4174), .Q (new_AGEMA_signal_4175) ) ;
    buf_clk new_AGEMA_reg_buffer_2823 ( .C (clk), .D (new_AGEMA_signal_4182), .Q (new_AGEMA_signal_4183) ) ;
    buf_clk new_AGEMA_reg_buffer_2831 ( .C (clk), .D (new_AGEMA_signal_4190), .Q (new_AGEMA_signal_4191) ) ;
    buf_clk new_AGEMA_reg_buffer_2839 ( .C (clk), .D (new_AGEMA_signal_4198), .Q (new_AGEMA_signal_4199) ) ;
    buf_clk new_AGEMA_reg_buffer_2847 ( .C (clk), .D (new_AGEMA_signal_4206), .Q (new_AGEMA_signal_4207) ) ;
    buf_clk new_AGEMA_reg_buffer_2855 ( .C (clk), .D (new_AGEMA_signal_4214), .Q (new_AGEMA_signal_4215) ) ;
    buf_clk new_AGEMA_reg_buffer_2863 ( .C (clk), .D (new_AGEMA_signal_4222), .Q (new_AGEMA_signal_4223) ) ;
    buf_clk new_AGEMA_reg_buffer_2871 ( .C (clk), .D (new_AGEMA_signal_4230), .Q (new_AGEMA_signal_4231) ) ;
    buf_clk new_AGEMA_reg_buffer_2879 ( .C (clk), .D (new_AGEMA_signal_4238), .Q (new_AGEMA_signal_4239) ) ;
    buf_clk new_AGEMA_reg_buffer_2887 ( .C (clk), .D (new_AGEMA_signal_4246), .Q (new_AGEMA_signal_4247) ) ;
    buf_clk new_AGEMA_reg_buffer_2895 ( .C (clk), .D (new_AGEMA_signal_4254), .Q (new_AGEMA_signal_4255) ) ;
    buf_clk new_AGEMA_reg_buffer_2903 ( .C (clk), .D (new_AGEMA_signal_4262), .Q (new_AGEMA_signal_4263) ) ;
    buf_clk new_AGEMA_reg_buffer_2911 ( .C (clk), .D (new_AGEMA_signal_4270), .Q (new_AGEMA_signal_4271) ) ;
    buf_clk new_AGEMA_reg_buffer_2919 ( .C (clk), .D (new_AGEMA_signal_4278), .Q (new_AGEMA_signal_4279) ) ;
    buf_clk new_AGEMA_reg_buffer_2927 ( .C (clk), .D (new_AGEMA_signal_4286), .Q (new_AGEMA_signal_4287) ) ;
    buf_clk new_AGEMA_reg_buffer_2935 ( .C (clk), .D (new_AGEMA_signal_4294), .Q (new_AGEMA_signal_4295) ) ;
    buf_clk new_AGEMA_reg_buffer_2943 ( .C (clk), .D (new_AGEMA_signal_4302), .Q (new_AGEMA_signal_4303) ) ;
    buf_clk new_AGEMA_reg_buffer_2951 ( .C (clk), .D (new_AGEMA_signal_4310), .Q (new_AGEMA_signal_4311) ) ;
    buf_clk new_AGEMA_reg_buffer_2959 ( .C (clk), .D (new_AGEMA_signal_4318), .Q (new_AGEMA_signal_4319) ) ;
    buf_clk new_AGEMA_reg_buffer_2967 ( .C (clk), .D (new_AGEMA_signal_4326), .Q (new_AGEMA_signal_4327) ) ;
    buf_clk new_AGEMA_reg_buffer_2975 ( .C (clk), .D (new_AGEMA_signal_4334), .Q (new_AGEMA_signal_4335) ) ;
    buf_clk new_AGEMA_reg_buffer_2983 ( .C (clk), .D (new_AGEMA_signal_4342), .Q (new_AGEMA_signal_4343) ) ;
    buf_clk new_AGEMA_reg_buffer_2991 ( .C (clk), .D (new_AGEMA_signal_4350), .Q (new_AGEMA_signal_4351) ) ;
    buf_clk new_AGEMA_reg_buffer_2999 ( .C (clk), .D (new_AGEMA_signal_4358), .Q (new_AGEMA_signal_4359) ) ;
    buf_clk new_AGEMA_reg_buffer_3007 ( .C (clk), .D (new_AGEMA_signal_4366), .Q (new_AGEMA_signal_4367) ) ;
    buf_clk new_AGEMA_reg_buffer_3015 ( .C (clk), .D (new_AGEMA_signal_4374), .Q (new_AGEMA_signal_4375) ) ;
    buf_clk new_AGEMA_reg_buffer_3023 ( .C (clk), .D (new_AGEMA_signal_4382), .Q (new_AGEMA_signal_4383) ) ;
    buf_clk new_AGEMA_reg_buffer_3031 ( .C (clk), .D (new_AGEMA_signal_4390), .Q (new_AGEMA_signal_4391) ) ;
    buf_clk new_AGEMA_reg_buffer_3039 ( .C (clk), .D (new_AGEMA_signal_4398), .Q (new_AGEMA_signal_4399) ) ;
    buf_clk new_AGEMA_reg_buffer_3047 ( .C (clk), .D (new_AGEMA_signal_4406), .Q (new_AGEMA_signal_4407) ) ;
    buf_clk new_AGEMA_reg_buffer_3055 ( .C (clk), .D (new_AGEMA_signal_4414), .Q (new_AGEMA_signal_4415) ) ;
    buf_clk new_AGEMA_reg_buffer_3063 ( .C (clk), .D (new_AGEMA_signal_4422), .Q (new_AGEMA_signal_4423) ) ;
    buf_clk new_AGEMA_reg_buffer_3067 ( .C (clk), .D (new_AGEMA_signal_3210), .Q (new_AGEMA_signal_4427) ) ;
    buf_clk new_AGEMA_reg_buffer_3069 ( .C (clk), .D (new_AGEMA_signal_3212), .Q (new_AGEMA_signal_4429) ) ;
    buf_clk new_AGEMA_reg_buffer_3073 ( .C (clk), .D (new_AGEMA_signal_4432), .Q (new_AGEMA_signal_4433) ) ;
    buf_clk new_AGEMA_reg_buffer_3077 ( .C (clk), .D (new_AGEMA_signal_4436), .Q (new_AGEMA_signal_4437) ) ;
    buf_clk new_AGEMA_reg_buffer_3079 ( .C (clk), .D (new_AGEMA_signal_3222), .Q (new_AGEMA_signal_4439) ) ;
    buf_clk new_AGEMA_reg_buffer_3081 ( .C (clk), .D (new_AGEMA_signal_3224), .Q (new_AGEMA_signal_4441) ) ;
    buf_clk new_AGEMA_reg_buffer_3085 ( .C (clk), .D (new_AGEMA_signal_4444), .Q (new_AGEMA_signal_4445) ) ;
    buf_clk new_AGEMA_reg_buffer_3089 ( .C (clk), .D (new_AGEMA_signal_4448), .Q (new_AGEMA_signal_4449) ) ;
    buf_clk new_AGEMA_reg_buffer_3091 ( .C (clk), .D (new_AGEMA_signal_3234), .Q (new_AGEMA_signal_4451) ) ;
    buf_clk new_AGEMA_reg_buffer_3093 ( .C (clk), .D (new_AGEMA_signal_3236), .Q (new_AGEMA_signal_4453) ) ;
    buf_clk new_AGEMA_reg_buffer_3097 ( .C (clk), .D (new_AGEMA_signal_4456), .Q (new_AGEMA_signal_4457) ) ;
    buf_clk new_AGEMA_reg_buffer_3101 ( .C (clk), .D (new_AGEMA_signal_4460), .Q (new_AGEMA_signal_4461) ) ;
    buf_clk new_AGEMA_reg_buffer_3103 ( .C (clk), .D (new_AGEMA_signal_3246), .Q (new_AGEMA_signal_4463) ) ;
    buf_clk new_AGEMA_reg_buffer_3105 ( .C (clk), .D (new_AGEMA_signal_3248), .Q (new_AGEMA_signal_4465) ) ;
    buf_clk new_AGEMA_reg_buffer_3109 ( .C (clk), .D (new_AGEMA_signal_4468), .Q (new_AGEMA_signal_4469) ) ;
    buf_clk new_AGEMA_reg_buffer_3113 ( .C (clk), .D (new_AGEMA_signal_4472), .Q (new_AGEMA_signal_4473) ) ;
    buf_clk new_AGEMA_reg_buffer_3115 ( .C (clk), .D (new_AGEMA_signal_3258), .Q (new_AGEMA_signal_4475) ) ;
    buf_clk new_AGEMA_reg_buffer_3117 ( .C (clk), .D (new_AGEMA_signal_3260), .Q (new_AGEMA_signal_4477) ) ;
    buf_clk new_AGEMA_reg_buffer_3121 ( .C (clk), .D (new_AGEMA_signal_4480), .Q (new_AGEMA_signal_4481) ) ;
    buf_clk new_AGEMA_reg_buffer_3125 ( .C (clk), .D (new_AGEMA_signal_4484), .Q (new_AGEMA_signal_4485) ) ;
    buf_clk new_AGEMA_reg_buffer_3127 ( .C (clk), .D (new_AGEMA_signal_3270), .Q (new_AGEMA_signal_4487) ) ;
    buf_clk new_AGEMA_reg_buffer_3129 ( .C (clk), .D (new_AGEMA_signal_3272), .Q (new_AGEMA_signal_4489) ) ;
    buf_clk new_AGEMA_reg_buffer_3133 ( .C (clk), .D (new_AGEMA_signal_4492), .Q (new_AGEMA_signal_4493) ) ;
    buf_clk new_AGEMA_reg_buffer_3137 ( .C (clk), .D (new_AGEMA_signal_4496), .Q (new_AGEMA_signal_4497) ) ;
    buf_clk new_AGEMA_reg_buffer_3139 ( .C (clk), .D (new_AGEMA_signal_3282), .Q (new_AGEMA_signal_4499) ) ;
    buf_clk new_AGEMA_reg_buffer_3141 ( .C (clk), .D (new_AGEMA_signal_3284), .Q (new_AGEMA_signal_4501) ) ;
    buf_clk new_AGEMA_reg_buffer_3145 ( .C (clk), .D (new_AGEMA_signal_4504), .Q (new_AGEMA_signal_4505) ) ;
    buf_clk new_AGEMA_reg_buffer_3149 ( .C (clk), .D (new_AGEMA_signal_4508), .Q (new_AGEMA_signal_4509) ) ;
    buf_clk new_AGEMA_reg_buffer_3151 ( .C (clk), .D (new_AGEMA_signal_3294), .Q (new_AGEMA_signal_4511) ) ;
    buf_clk new_AGEMA_reg_buffer_3153 ( .C (clk), .D (new_AGEMA_signal_3296), .Q (new_AGEMA_signal_4513) ) ;
    buf_clk new_AGEMA_reg_buffer_3157 ( .C (clk), .D (new_AGEMA_signal_4516), .Q (new_AGEMA_signal_4517) ) ;
    buf_clk new_AGEMA_reg_buffer_3161 ( .C (clk), .D (new_AGEMA_signal_4520), .Q (new_AGEMA_signal_4521) ) ;
    buf_clk new_AGEMA_reg_buffer_3163 ( .C (clk), .D (new_AGEMA_signal_3306), .Q (new_AGEMA_signal_4523) ) ;
    buf_clk new_AGEMA_reg_buffer_3165 ( .C (clk), .D (new_AGEMA_signal_3308), .Q (new_AGEMA_signal_4525) ) ;
    buf_clk new_AGEMA_reg_buffer_3169 ( .C (clk), .D (new_AGEMA_signal_4528), .Q (new_AGEMA_signal_4529) ) ;
    buf_clk new_AGEMA_reg_buffer_3173 ( .C (clk), .D (new_AGEMA_signal_4532), .Q (new_AGEMA_signal_4533) ) ;
    buf_clk new_AGEMA_reg_buffer_3175 ( .C (clk), .D (new_AGEMA_signal_3318), .Q (new_AGEMA_signal_4535) ) ;
    buf_clk new_AGEMA_reg_buffer_3177 ( .C (clk), .D (new_AGEMA_signal_3320), .Q (new_AGEMA_signal_4537) ) ;
    buf_clk new_AGEMA_reg_buffer_3181 ( .C (clk), .D (new_AGEMA_signal_4540), .Q (new_AGEMA_signal_4541) ) ;
    buf_clk new_AGEMA_reg_buffer_3185 ( .C (clk), .D (new_AGEMA_signal_4544), .Q (new_AGEMA_signal_4545) ) ;
    buf_clk new_AGEMA_reg_buffer_3187 ( .C (clk), .D (new_AGEMA_signal_3330), .Q (new_AGEMA_signal_4547) ) ;
    buf_clk new_AGEMA_reg_buffer_3189 ( .C (clk), .D (new_AGEMA_signal_3332), .Q (new_AGEMA_signal_4549) ) ;
    buf_clk new_AGEMA_reg_buffer_3193 ( .C (clk), .D (new_AGEMA_signal_4552), .Q (new_AGEMA_signal_4553) ) ;
    buf_clk new_AGEMA_reg_buffer_3197 ( .C (clk), .D (new_AGEMA_signal_4556), .Q (new_AGEMA_signal_4557) ) ;
    buf_clk new_AGEMA_reg_buffer_3199 ( .C (clk), .D (new_AGEMA_signal_3342), .Q (new_AGEMA_signal_4559) ) ;
    buf_clk new_AGEMA_reg_buffer_3201 ( .C (clk), .D (new_AGEMA_signal_3344), .Q (new_AGEMA_signal_4561) ) ;
    buf_clk new_AGEMA_reg_buffer_3205 ( .C (clk), .D (new_AGEMA_signal_4564), .Q (new_AGEMA_signal_4565) ) ;
    buf_clk new_AGEMA_reg_buffer_3209 ( .C (clk), .D (new_AGEMA_signal_4568), .Q (new_AGEMA_signal_4569) ) ;
    buf_clk new_AGEMA_reg_buffer_3211 ( .C (clk), .D (new_AGEMA_signal_3354), .Q (new_AGEMA_signal_4571) ) ;
    buf_clk new_AGEMA_reg_buffer_3213 ( .C (clk), .D (new_AGEMA_signal_3356), .Q (new_AGEMA_signal_4573) ) ;
    buf_clk new_AGEMA_reg_buffer_3217 ( .C (clk), .D (new_AGEMA_signal_4576), .Q (new_AGEMA_signal_4577) ) ;
    buf_clk new_AGEMA_reg_buffer_3221 ( .C (clk), .D (new_AGEMA_signal_4580), .Q (new_AGEMA_signal_4581) ) ;
    buf_clk new_AGEMA_reg_buffer_3223 ( .C (clk), .D (new_AGEMA_signal_3366), .Q (new_AGEMA_signal_4583) ) ;
    buf_clk new_AGEMA_reg_buffer_3225 ( .C (clk), .D (new_AGEMA_signal_3368), .Q (new_AGEMA_signal_4585) ) ;
    buf_clk new_AGEMA_reg_buffer_3229 ( .C (clk), .D (new_AGEMA_signal_4588), .Q (new_AGEMA_signal_4589) ) ;
    buf_clk new_AGEMA_reg_buffer_3233 ( .C (clk), .D (new_AGEMA_signal_4592), .Q (new_AGEMA_signal_4593) ) ;
    buf_clk new_AGEMA_reg_buffer_3235 ( .C (clk), .D (new_AGEMA_signal_3378), .Q (new_AGEMA_signal_4595) ) ;
    buf_clk new_AGEMA_reg_buffer_3237 ( .C (clk), .D (new_AGEMA_signal_3380), .Q (new_AGEMA_signal_4597) ) ;
    buf_clk new_AGEMA_reg_buffer_3241 ( .C (clk), .D (new_AGEMA_signal_4600), .Q (new_AGEMA_signal_4601) ) ;
    buf_clk new_AGEMA_reg_buffer_3245 ( .C (clk), .D (new_AGEMA_signal_4604), .Q (new_AGEMA_signal_4605) ) ;
    buf_clk new_AGEMA_reg_buffer_3247 ( .C (clk), .D (new_AGEMA_signal_3390), .Q (new_AGEMA_signal_4607) ) ;
    buf_clk new_AGEMA_reg_buffer_3249 ( .C (clk), .D (new_AGEMA_signal_3392), .Q (new_AGEMA_signal_4609) ) ;
    buf_clk new_AGEMA_reg_buffer_3253 ( .C (clk), .D (new_AGEMA_signal_4612), .Q (new_AGEMA_signal_4613) ) ;
    buf_clk new_AGEMA_reg_buffer_3257 ( .C (clk), .D (new_AGEMA_signal_4616), .Q (new_AGEMA_signal_4617) ) ;
    buf_clk new_AGEMA_reg_buffer_3391 ( .C (clk), .D (new_AGEMA_signal_4750), .Q (new_AGEMA_signal_4751) ) ;
    buf_clk new_AGEMA_reg_buffer_3399 ( .C (clk), .D (new_AGEMA_signal_4758), .Q (new_AGEMA_signal_4759) ) ;
    buf_clk new_AGEMA_reg_buffer_3407 ( .C (clk), .D (new_AGEMA_signal_4766), .Q (new_AGEMA_signal_4767) ) ;
    buf_clk new_AGEMA_reg_buffer_3415 ( .C (clk), .D (new_AGEMA_signal_4774), .Q (new_AGEMA_signal_4775) ) ;
    buf_clk new_AGEMA_reg_buffer_3423 ( .C (clk), .D (new_AGEMA_signal_4782), .Q (new_AGEMA_signal_4783) ) ;
    buf_clk new_AGEMA_reg_buffer_3431 ( .C (clk), .D (new_AGEMA_signal_4790), .Q (new_AGEMA_signal_4791) ) ;
    buf_clk new_AGEMA_reg_buffer_3439 ( .C (clk), .D (new_AGEMA_signal_4798), .Q (new_AGEMA_signal_4799) ) ;
    buf_clk new_AGEMA_reg_buffer_3447 ( .C (clk), .D (new_AGEMA_signal_4806), .Q (new_AGEMA_signal_4807) ) ;
    buf_clk new_AGEMA_reg_buffer_3455 ( .C (clk), .D (new_AGEMA_signal_4814), .Q (new_AGEMA_signal_4815) ) ;
    buf_clk new_AGEMA_reg_buffer_3463 ( .C (clk), .D (new_AGEMA_signal_4822), .Q (new_AGEMA_signal_4823) ) ;

    /* cells in depth 6 */
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_1_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1373, Feedback[1]}), .a ({new_AGEMA_signal_2452, new_AGEMA_signal_2446}), .c ({new_AGEMA_signal_1582, MCOutput[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_3_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1371, Feedback[3]}), .a ({new_AGEMA_signal_2464, new_AGEMA_signal_2458}), .c ({new_AGEMA_signal_1586, MCOutput[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_5_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1377, Feedback[5]}), .a ({new_AGEMA_signal_2476, new_AGEMA_signal_2470}), .c ({new_AGEMA_signal_1590, MCOutput[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_7_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1375, Feedback[7]}), .a ({new_AGEMA_signal_2488, new_AGEMA_signal_2482}), .c ({new_AGEMA_signal_1594, MCOutput[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_9_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1381, Feedback[9]}), .a ({new_AGEMA_signal_2500, new_AGEMA_signal_2494}), .c ({new_AGEMA_signal_1598, MCOutput[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_11_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1379, Feedback[11]}), .a ({new_AGEMA_signal_2512, new_AGEMA_signal_2506}), .c ({new_AGEMA_signal_1602, MCOutput[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_13_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1385, Feedback[13]}), .a ({new_AGEMA_signal_2524, new_AGEMA_signal_2518}), .c ({new_AGEMA_signal_1606, MCOutput[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_15_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1383, Feedback[15]}), .a ({new_AGEMA_signal_2536, new_AGEMA_signal_2530}), .c ({new_AGEMA_signal_1610, MCOutput[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_17_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1389, Feedback[17]}), .a ({new_AGEMA_signal_2548, new_AGEMA_signal_2542}), .c ({new_AGEMA_signal_1614, MCOutput[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_19_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1387, Feedback[19]}), .a ({new_AGEMA_signal_2560, new_AGEMA_signal_2554}), .c ({new_AGEMA_signal_1618, MCOutput[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_21_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1393, Feedback[21]}), .a ({new_AGEMA_signal_2572, new_AGEMA_signal_2566}), .c ({new_AGEMA_signal_1622, MCOutput[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_23_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1391, Feedback[23]}), .a ({new_AGEMA_signal_2584, new_AGEMA_signal_2578}), .c ({new_AGEMA_signal_1626, MCOutput[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_25_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1397, Feedback[25]}), .a ({new_AGEMA_signal_2596, new_AGEMA_signal_2590}), .c ({new_AGEMA_signal_1630, MCOutput[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_27_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1395, Feedback[27]}), .a ({new_AGEMA_signal_2608, new_AGEMA_signal_2602}), .c ({new_AGEMA_signal_1634, MCOutput[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_29_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1401, Feedback[29]}), .a ({new_AGEMA_signal_2620, new_AGEMA_signal_2614}), .c ({new_AGEMA_signal_1638, MCOutput[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_31_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1399, Feedback[31]}), .a ({new_AGEMA_signal_2632, new_AGEMA_signal_2626}), .c ({new_AGEMA_signal_1642, MCOutput[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_33_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1405, Feedback[33]}), .a ({new_AGEMA_signal_2644, new_AGEMA_signal_2638}), .c ({new_AGEMA_signal_1646, MCInput[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_35_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1403, Feedback[35]}), .a ({new_AGEMA_signal_2656, new_AGEMA_signal_2650}), .c ({new_AGEMA_signal_1650, MCInput[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_37_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1409, Feedback[37]}), .a ({new_AGEMA_signal_2668, new_AGEMA_signal_2662}), .c ({new_AGEMA_signal_1654, MCInput[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_39_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1407, Feedback[39]}), .a ({new_AGEMA_signal_2680, new_AGEMA_signal_2674}), .c ({new_AGEMA_signal_1658, MCInput[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_41_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1413, Feedback[41]}), .a ({new_AGEMA_signal_2692, new_AGEMA_signal_2686}), .c ({new_AGEMA_signal_1662, MCInput[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_43_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1411, Feedback[43]}), .a ({new_AGEMA_signal_2704, new_AGEMA_signal_2698}), .c ({new_AGEMA_signal_1666, MCInput[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_45_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1417, Feedback[45]}), .a ({new_AGEMA_signal_2716, new_AGEMA_signal_2710}), .c ({new_AGEMA_signal_1670, MCInput[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_47_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1415, Feedback[47]}), .a ({new_AGEMA_signal_2728, new_AGEMA_signal_2722}), .c ({new_AGEMA_signal_1674, MCInput[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_49_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1421, Feedback[49]}), .a ({new_AGEMA_signal_2740, new_AGEMA_signal_2734}), .c ({new_AGEMA_signal_1678, MCInput[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_51_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1419, Feedback[51]}), .a ({new_AGEMA_signal_2752, new_AGEMA_signal_2746}), .c ({new_AGEMA_signal_1682, MCInput[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_53_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1425, Feedback[53]}), .a ({new_AGEMA_signal_2764, new_AGEMA_signal_2758}), .c ({new_AGEMA_signal_1686, MCInput[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_55_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1423, Feedback[55]}), .a ({new_AGEMA_signal_2776, new_AGEMA_signal_2770}), .c ({new_AGEMA_signal_1690, MCInput[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_57_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1429, Feedback[57]}), .a ({new_AGEMA_signal_2788, new_AGEMA_signal_2782}), .c ({new_AGEMA_signal_1694, MCInput[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_59_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1427, Feedback[59]}), .a ({new_AGEMA_signal_2800, new_AGEMA_signal_2794}), .c ({new_AGEMA_signal_1698, MCInput[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_61_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1433, Feedback[61]}), .a ({new_AGEMA_signal_2812, new_AGEMA_signal_2806}), .c ({new_AGEMA_signal_1702, MCInput[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_63_U1 ( .s (new_AGEMA_signal_2440), .b ({new_AGEMA_signal_1431, Feedback[63]}), .a ({new_AGEMA_signal_2824, new_AGEMA_signal_2818}), .c ({new_AGEMA_signal_1706, MCInput[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_1_U3 ( .a ({new_AGEMA_signal_1719, MCInst_XOR_r0_Inst_1_n2}), .b ({new_AGEMA_signal_1718, MCInst_XOR_r0_Inst_1_n1}), .c ({new_AGEMA_signal_1797, MCOutput[49]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_1_U2 ( .a ({new_AGEMA_signal_1614, MCOutput[17]}), .b ({new_AGEMA_signal_1582, MCOutput[1]}), .c ({new_AGEMA_signal_1718, MCInst_XOR_r0_Inst_1_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1678, MCInput[49]}), .c ({new_AGEMA_signal_1719, MCInst_XOR_r0_Inst_1_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_1_U2 ( .a ({new_AGEMA_signal_1720, MCInst_XOR_r1_Inst_1_n1}), .b ({new_AGEMA_signal_1582, MCOutput[1]}), .c ({new_AGEMA_signal_1798, MCOutput[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1646, MCInput[33]}), .c ({new_AGEMA_signal_1720, MCInst_XOR_r1_Inst_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_3_U3 ( .a ({new_AGEMA_signal_1725, MCInst_XOR_r0_Inst_3_n2}), .b ({new_AGEMA_signal_1724, MCInst_XOR_r0_Inst_3_n1}), .c ({new_AGEMA_signal_1801, MCOutput[51]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_3_U2 ( .a ({new_AGEMA_signal_1618, MCOutput[19]}), .b ({new_AGEMA_signal_1586, MCOutput[3]}), .c ({new_AGEMA_signal_1724, MCInst_XOR_r0_Inst_3_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1682, MCInput[51]}), .c ({new_AGEMA_signal_1725, MCInst_XOR_r0_Inst_3_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_3_U2 ( .a ({new_AGEMA_signal_1726, MCInst_XOR_r1_Inst_3_n1}), .b ({new_AGEMA_signal_1586, MCOutput[3]}), .c ({new_AGEMA_signal_1802, MCOutput[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1650, MCInput[35]}), .c ({new_AGEMA_signal_1726, MCInst_XOR_r1_Inst_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_5_U3 ( .a ({new_AGEMA_signal_1731, MCInst_XOR_r0_Inst_5_n2}), .b ({new_AGEMA_signal_1730, MCInst_XOR_r0_Inst_5_n1}), .c ({new_AGEMA_signal_1805, MCOutput[53]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_5_U2 ( .a ({new_AGEMA_signal_1622, MCOutput[21]}), .b ({new_AGEMA_signal_1590, MCOutput[5]}), .c ({new_AGEMA_signal_1730, MCInst_XOR_r0_Inst_5_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_5_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1686, MCInput[53]}), .c ({new_AGEMA_signal_1731, MCInst_XOR_r0_Inst_5_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_5_U2 ( .a ({new_AGEMA_signal_1732, MCInst_XOR_r1_Inst_5_n1}), .b ({new_AGEMA_signal_1590, MCOutput[5]}), .c ({new_AGEMA_signal_1806, MCOutput[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_5_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1654, MCInput[37]}), .c ({new_AGEMA_signal_1732, MCInst_XOR_r1_Inst_5_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_7_U3 ( .a ({new_AGEMA_signal_1737, MCInst_XOR_r0_Inst_7_n2}), .b ({new_AGEMA_signal_1736, MCInst_XOR_r0_Inst_7_n1}), .c ({new_AGEMA_signal_1809, MCOutput[55]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_7_U2 ( .a ({new_AGEMA_signal_1626, MCOutput[23]}), .b ({new_AGEMA_signal_1594, MCOutput[7]}), .c ({new_AGEMA_signal_1736, MCInst_XOR_r0_Inst_7_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_7_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1690, MCInput[55]}), .c ({new_AGEMA_signal_1737, MCInst_XOR_r0_Inst_7_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_7_U2 ( .a ({new_AGEMA_signal_1738, MCInst_XOR_r1_Inst_7_n1}), .b ({new_AGEMA_signal_1594, MCOutput[7]}), .c ({new_AGEMA_signal_1810, MCOutput[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_7_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1658, MCInput[39]}), .c ({new_AGEMA_signal_1738, MCInst_XOR_r1_Inst_7_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_9_U3 ( .a ({new_AGEMA_signal_1743, MCInst_XOR_r0_Inst_9_n2}), .b ({new_AGEMA_signal_1742, MCInst_XOR_r0_Inst_9_n1}), .c ({new_AGEMA_signal_1813, MCOutput[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_9_U2 ( .a ({new_AGEMA_signal_1630, MCOutput[25]}), .b ({new_AGEMA_signal_1598, MCOutput[9]}), .c ({new_AGEMA_signal_1742, MCInst_XOR_r0_Inst_9_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_9_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1694, MCInput[57]}), .c ({new_AGEMA_signal_1743, MCInst_XOR_r0_Inst_9_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_9_U2 ( .a ({new_AGEMA_signal_1744, MCInst_XOR_r1_Inst_9_n1}), .b ({new_AGEMA_signal_1598, MCOutput[9]}), .c ({new_AGEMA_signal_1814, MCOutput[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_9_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1662, MCInput[41]}), .c ({new_AGEMA_signal_1744, MCInst_XOR_r1_Inst_9_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_11_U3 ( .a ({new_AGEMA_signal_1749, MCInst_XOR_r0_Inst_11_n2}), .b ({new_AGEMA_signal_1748, MCInst_XOR_r0_Inst_11_n1}), .c ({new_AGEMA_signal_1817, MCOutput[59]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_11_U2 ( .a ({new_AGEMA_signal_1634, MCOutput[27]}), .b ({new_AGEMA_signal_1602, MCOutput[11]}), .c ({new_AGEMA_signal_1748, MCInst_XOR_r0_Inst_11_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_11_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1698, MCInput[59]}), .c ({new_AGEMA_signal_1749, MCInst_XOR_r0_Inst_11_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_11_U2 ( .a ({new_AGEMA_signal_1750, MCInst_XOR_r1_Inst_11_n1}), .b ({new_AGEMA_signal_1602, MCOutput[11]}), .c ({new_AGEMA_signal_1818, MCOutput[43]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_11_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1666, MCInput[43]}), .c ({new_AGEMA_signal_1750, MCInst_XOR_r1_Inst_11_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_13_U3 ( .a ({new_AGEMA_signal_1755, MCInst_XOR_r0_Inst_13_n2}), .b ({new_AGEMA_signal_1754, MCInst_XOR_r0_Inst_13_n1}), .c ({new_AGEMA_signal_1821, MCOutput[61]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_13_U2 ( .a ({new_AGEMA_signal_1638, MCOutput[29]}), .b ({new_AGEMA_signal_1606, MCOutput[13]}), .c ({new_AGEMA_signal_1754, MCInst_XOR_r0_Inst_13_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_13_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1702, MCInput[61]}), .c ({new_AGEMA_signal_1755, MCInst_XOR_r0_Inst_13_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_13_U2 ( .a ({new_AGEMA_signal_1756, MCInst_XOR_r1_Inst_13_n1}), .b ({new_AGEMA_signal_1606, MCOutput[13]}), .c ({new_AGEMA_signal_1822, MCOutput[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_13_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1670, MCInput[45]}), .c ({new_AGEMA_signal_1756, MCInst_XOR_r1_Inst_13_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_15_U3 ( .a ({new_AGEMA_signal_1761, MCInst_XOR_r0_Inst_15_n2}), .b ({new_AGEMA_signal_1760, MCInst_XOR_r0_Inst_15_n1}), .c ({new_AGEMA_signal_1825, MCOutput[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_15_U2 ( .a ({new_AGEMA_signal_1642, MCOutput[31]}), .b ({new_AGEMA_signal_1610, MCOutput[15]}), .c ({new_AGEMA_signal_1760, MCInst_XOR_r0_Inst_15_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_15_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1706, MCInput[63]}), .c ({new_AGEMA_signal_1761, MCInst_XOR_r0_Inst_15_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_15_U2 ( .a ({new_AGEMA_signal_1762, MCInst_XOR_r1_Inst_15_n1}), .b ({new_AGEMA_signal_1610, MCOutput[15]}), .c ({new_AGEMA_signal_1826, MCOutput[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_15_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1674, MCInput[47]}), .c ({new_AGEMA_signal_1762, MCInst_XOR_r1_Inst_15_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_1860, AddKeyXOR1_XORInst_0_1_n1}), .b ({new_AGEMA_signal_2836, new_AGEMA_signal_2830}), .c ({new_AGEMA_signal_1892, AddRoundKeyOutput[49]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_0_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1797, MCOutput[49]}), .c ({new_AGEMA_signal_1860, AddKeyXOR1_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_1862, AddKeyXOR1_XORInst_0_3_n1}), .b ({new_AGEMA_signal_2848, new_AGEMA_signal_2842}), .c ({new_AGEMA_signal_1894, AddRoundKeyOutput[51]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_0_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1801, MCOutput[51]}), .c ({new_AGEMA_signal_1862, AddKeyXOR1_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_1864, AddKeyXOR1_XORInst_1_1_n1}), .b ({new_AGEMA_signal_2860, new_AGEMA_signal_2854}), .c ({new_AGEMA_signal_1896, AddRoundKeyOutput[53]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_1_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1805, MCOutput[53]}), .c ({new_AGEMA_signal_1864, AddKeyXOR1_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_1866, AddKeyXOR1_XORInst_1_3_n1}), .b ({new_AGEMA_signal_2872, new_AGEMA_signal_2866}), .c ({new_AGEMA_signal_1898, AddRoundKeyOutput[55]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_1_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1809, MCOutput[55]}), .c ({new_AGEMA_signal_1866, AddKeyXOR1_XORInst_1_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_1868, AddKeyXOR1_XORInst_2_1_n1}), .b ({new_AGEMA_signal_2884, new_AGEMA_signal_2878}), .c ({new_AGEMA_signal_1900, AddRoundKeyOutput[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_2_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1813, MCOutput[57]}), .c ({new_AGEMA_signal_1868, AddKeyXOR1_XORInst_2_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_1870, AddKeyXOR1_XORInst_2_3_n1}), .b ({new_AGEMA_signal_2896, new_AGEMA_signal_2890}), .c ({new_AGEMA_signal_1902, AddRoundKeyOutput[59]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_2_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1817, MCOutput[59]}), .c ({new_AGEMA_signal_1870, AddKeyXOR1_XORInst_2_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_1872, AddKeyXOR1_XORInst_3_1_n1}), .b ({new_AGEMA_signal_2908, new_AGEMA_signal_2902}), .c ({new_AGEMA_signal_1904, AddRoundKeyOutput[61]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_3_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1821, MCOutput[61]}), .c ({new_AGEMA_signal_1872, AddKeyXOR1_XORInst_3_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_1874, AddKeyXOR1_XORInst_3_3_n1}), .b ({new_AGEMA_signal_2920, new_AGEMA_signal_2914}), .c ({new_AGEMA_signal_1906, AddRoundKeyOutput[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_3_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1825, MCOutput[63]}), .c ({new_AGEMA_signal_1874, AddKeyXOR1_XORInst_3_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_1_U3 ( .a ({new_AGEMA_signal_1876, AddKeyConstXOR_XORInst_0_1_n2}), .b ({new_AGEMA_signal_2932, new_AGEMA_signal_2926}), .c ({new_AGEMA_signal_1908, AddRoundKeyOutput[41]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1814, MCOutput[41]}), .c ({new_AGEMA_signal_1876, AddKeyConstXOR_XORInst_0_1_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_3_U3 ( .a ({new_AGEMA_signal_1878, AddKeyConstXOR_XORInst_0_3_n2}), .b ({new_AGEMA_signal_2944, new_AGEMA_signal_2938}), .c ({new_AGEMA_signal_1910, AddRoundKeyOutput[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1818, MCOutput[43]}), .c ({new_AGEMA_signal_1878, AddKeyConstXOR_XORInst_0_3_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_1_U3 ( .a ({new_AGEMA_signal_1880, AddKeyConstXOR_XORInst_1_1_n2}), .b ({new_AGEMA_signal_2956, new_AGEMA_signal_2950}), .c ({new_AGEMA_signal_1912, AddRoundKeyOutput[45]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1822, MCOutput[45]}), .c ({new_AGEMA_signal_1880, AddKeyConstXOR_XORInst_1_1_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_3_U3 ( .a ({new_AGEMA_signal_1882, AddKeyConstXOR_XORInst_1_3_n2}), .b ({new_AGEMA_signal_2968, new_AGEMA_signal_2962}), .c ({new_AGEMA_signal_1914, AddRoundKeyOutput[47]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1826, MCOutput[47]}), .c ({new_AGEMA_signal_1882, AddKeyConstXOR_XORInst_1_3_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_1764, AddKeyXOR2_XORInst_0_1_n1}), .b ({new_AGEMA_signal_2980, new_AGEMA_signal_2974}), .c ({new_AGEMA_signal_1828, AddRoundKeyOutput[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_0_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1582, MCOutput[1]}), .c ({new_AGEMA_signal_1764, AddKeyXOR2_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_1766, AddKeyXOR2_XORInst_0_3_n1}), .b ({new_AGEMA_signal_2992, new_AGEMA_signal_2986}), .c ({new_AGEMA_signal_1830, AddRoundKeyOutput[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_0_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1586, MCOutput[3]}), .c ({new_AGEMA_signal_1766, AddKeyXOR2_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_1768, AddKeyXOR2_XORInst_1_1_n1}), .b ({new_AGEMA_signal_3004, new_AGEMA_signal_2998}), .c ({new_AGEMA_signal_1832, AddRoundKeyOutput[5]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_1_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1590, MCOutput[5]}), .c ({new_AGEMA_signal_1768, AddKeyXOR2_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_1770, AddKeyXOR2_XORInst_1_3_n1}), .b ({new_AGEMA_signal_3016, new_AGEMA_signal_3010}), .c ({new_AGEMA_signal_1834, AddRoundKeyOutput[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_1_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1594, MCOutput[7]}), .c ({new_AGEMA_signal_1770, AddKeyXOR2_XORInst_1_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_1772, AddKeyXOR2_XORInst_2_1_n1}), .b ({new_AGEMA_signal_3028, new_AGEMA_signal_3022}), .c ({new_AGEMA_signal_1836, AddRoundKeyOutput[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_2_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1598, MCOutput[9]}), .c ({new_AGEMA_signal_1772, AddKeyXOR2_XORInst_2_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_1774, AddKeyXOR2_XORInst_2_3_n1}), .b ({new_AGEMA_signal_3040, new_AGEMA_signal_3034}), .c ({new_AGEMA_signal_1838, AddRoundKeyOutput[11]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_2_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1602, MCOutput[11]}), .c ({new_AGEMA_signal_1774, AddKeyXOR2_XORInst_2_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_1776, AddKeyXOR2_XORInst_3_1_n1}), .b ({new_AGEMA_signal_3052, new_AGEMA_signal_3046}), .c ({new_AGEMA_signal_1840, AddRoundKeyOutput[13]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_3_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1606, MCOutput[13]}), .c ({new_AGEMA_signal_1776, AddKeyXOR2_XORInst_3_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_1778, AddKeyXOR2_XORInst_3_3_n1}), .b ({new_AGEMA_signal_3064, new_AGEMA_signal_3058}), .c ({new_AGEMA_signal_1842, AddRoundKeyOutput[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_3_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1610, MCOutput[15]}), .c ({new_AGEMA_signal_1778, AddKeyXOR2_XORInst_3_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_4_1_U2 ( .a ({new_AGEMA_signal_1780, AddKeyXOR2_XORInst_4_1_n1}), .b ({new_AGEMA_signal_3076, new_AGEMA_signal_3070}), .c ({new_AGEMA_signal_1844, AddRoundKeyOutput[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_4_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1614, MCOutput[17]}), .c ({new_AGEMA_signal_1780, AddKeyXOR2_XORInst_4_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_4_3_U2 ( .a ({new_AGEMA_signal_1782, AddKeyXOR2_XORInst_4_3_n1}), .b ({new_AGEMA_signal_3088, new_AGEMA_signal_3082}), .c ({new_AGEMA_signal_1846, AddRoundKeyOutput[19]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_4_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1618, MCOutput[19]}), .c ({new_AGEMA_signal_1782, AddKeyXOR2_XORInst_4_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_5_1_U2 ( .a ({new_AGEMA_signal_1784, AddKeyXOR2_XORInst_5_1_n1}), .b ({new_AGEMA_signal_3100, new_AGEMA_signal_3094}), .c ({new_AGEMA_signal_1848, AddRoundKeyOutput[21]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_5_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1622, MCOutput[21]}), .c ({new_AGEMA_signal_1784, AddKeyXOR2_XORInst_5_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_5_3_U2 ( .a ({new_AGEMA_signal_1786, AddKeyXOR2_XORInst_5_3_n1}), .b ({new_AGEMA_signal_3112, new_AGEMA_signal_3106}), .c ({new_AGEMA_signal_1850, AddRoundKeyOutput[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_5_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1626, MCOutput[23]}), .c ({new_AGEMA_signal_1786, AddKeyXOR2_XORInst_5_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_6_1_U2 ( .a ({new_AGEMA_signal_1788, AddKeyXOR2_XORInst_6_1_n1}), .b ({new_AGEMA_signal_3124, new_AGEMA_signal_3118}), .c ({new_AGEMA_signal_1852, AddRoundKeyOutput[25]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_6_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1630, MCOutput[25]}), .c ({new_AGEMA_signal_1788, AddKeyXOR2_XORInst_6_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_6_3_U2 ( .a ({new_AGEMA_signal_1790, AddKeyXOR2_XORInst_6_3_n1}), .b ({new_AGEMA_signal_3136, new_AGEMA_signal_3130}), .c ({new_AGEMA_signal_1854, AddRoundKeyOutput[27]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_6_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1634, MCOutput[27]}), .c ({new_AGEMA_signal_1790, AddKeyXOR2_XORInst_6_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_7_1_U2 ( .a ({new_AGEMA_signal_1792, AddKeyXOR2_XORInst_7_1_n1}), .b ({new_AGEMA_signal_3148, new_AGEMA_signal_3142}), .c ({new_AGEMA_signal_1856, AddRoundKeyOutput[29]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_7_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1638, MCOutput[29]}), .c ({new_AGEMA_signal_1792, AddKeyXOR2_XORInst_7_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_7_3_U2 ( .a ({new_AGEMA_signal_1794, AddKeyXOR2_XORInst_7_3_n1}), .b ({new_AGEMA_signal_3160, new_AGEMA_signal_3154}), .c ({new_AGEMA_signal_1858, AddRoundKeyOutput[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_7_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1642, MCOutput[31]}), .c ({new_AGEMA_signal_1794, AddKeyXOR2_XORInst_7_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_8_1_U2 ( .a ({new_AGEMA_signal_1884, AddKeyXOR2_XORInst_8_1_n1}), .b ({new_AGEMA_signal_3172, new_AGEMA_signal_3166}), .c ({new_AGEMA_signal_1916, AddRoundKeyOutput[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_8_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1798, MCOutput[33]}), .c ({new_AGEMA_signal_1884, AddKeyXOR2_XORInst_8_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_8_3_U2 ( .a ({new_AGEMA_signal_1886, AddKeyXOR2_XORInst_8_3_n1}), .b ({new_AGEMA_signal_3184, new_AGEMA_signal_3178}), .c ({new_AGEMA_signal_1918, AddRoundKeyOutput[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_8_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1802, MCOutput[35]}), .c ({new_AGEMA_signal_1886, AddKeyXOR2_XORInst_8_3_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_9_1_U2 ( .a ({new_AGEMA_signal_1888, AddKeyXOR2_XORInst_9_1_n1}), .b ({new_AGEMA_signal_3196, new_AGEMA_signal_3190}), .c ({new_AGEMA_signal_1920, AddRoundKeyOutput[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_9_1_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1806, MCOutput[37]}), .c ({new_AGEMA_signal_1888, AddKeyXOR2_XORInst_9_1_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_9_3_U2 ( .a ({new_AGEMA_signal_1890, AddKeyXOR2_XORInst_9_3_n1}), .b ({new_AGEMA_signal_3208, new_AGEMA_signal_3202}), .c ({new_AGEMA_signal_1922, AddRoundKeyOutput[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_9_3_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1810, MCOutput[39]}), .c ({new_AGEMA_signal_1890, AddKeyXOR2_XORInst_9_3_n1}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U19 ( .a ({new_AGEMA_signal_3212, new_AGEMA_signal_3210}), .b ({new_AGEMA_signal_1292, SubCellInst_SboxInst_0_n14}), .clk (clk), .r (Fresh[160]), .c ({new_AGEMA_signal_1371, Feedback[3]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U16 ( .a ({new_AGEMA_signal_1147, SubCellInst_SboxInst_0_n11}), .b ({new_AGEMA_signal_3216, new_AGEMA_signal_3214}), .clk (clk), .r (Fresh[161]), .c ({new_AGEMA_signal_1293, SubCellInst_SboxInst_0_n12}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U12 ( .a ({new_AGEMA_signal_3220, new_AGEMA_signal_3218}), .b ({new_AGEMA_signal_1294, SubCellInst_SboxInst_0_n5}), .clk (clk), .r (Fresh[162]), .c ({new_AGEMA_signal_1373, Feedback[1]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U7 ( .a ({new_AGEMA_signal_3216, new_AGEMA_signal_3214}), .b ({new_AGEMA_signal_1151, SubCellInst_SboxInst_0_n2}), .clk (clk), .r (Fresh[163]), .c ({new_AGEMA_signal_1295, SubCellInst_SboxInst_0_n3}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U19 ( .a ({new_AGEMA_signal_3224, new_AGEMA_signal_3222}), .b ({new_AGEMA_signal_1297, SubCellInst_SboxInst_1_n14}), .clk (clk), .r (Fresh[164]), .c ({new_AGEMA_signal_1375, Feedback[7]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U16 ( .a ({new_AGEMA_signal_1153, SubCellInst_SboxInst_1_n11}), .b ({new_AGEMA_signal_3228, new_AGEMA_signal_3226}), .clk (clk), .r (Fresh[165]), .c ({new_AGEMA_signal_1298, SubCellInst_SboxInst_1_n12}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U12 ( .a ({new_AGEMA_signal_3232, new_AGEMA_signal_3230}), .b ({new_AGEMA_signal_1299, SubCellInst_SboxInst_1_n5}), .clk (clk), .r (Fresh[166]), .c ({new_AGEMA_signal_1377, Feedback[5]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U7 ( .a ({new_AGEMA_signal_3228, new_AGEMA_signal_3226}), .b ({new_AGEMA_signal_1157, SubCellInst_SboxInst_1_n2}), .clk (clk), .r (Fresh[167]), .c ({new_AGEMA_signal_1300, SubCellInst_SboxInst_1_n3}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U19 ( .a ({new_AGEMA_signal_3236, new_AGEMA_signal_3234}), .b ({new_AGEMA_signal_1302, SubCellInst_SboxInst_2_n14}), .clk (clk), .r (Fresh[168]), .c ({new_AGEMA_signal_1379, Feedback[11]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U16 ( .a ({new_AGEMA_signal_1159, SubCellInst_SboxInst_2_n11}), .b ({new_AGEMA_signal_3240, new_AGEMA_signal_3238}), .clk (clk), .r (Fresh[169]), .c ({new_AGEMA_signal_1303, SubCellInst_SboxInst_2_n12}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U12 ( .a ({new_AGEMA_signal_3244, new_AGEMA_signal_3242}), .b ({new_AGEMA_signal_1304, SubCellInst_SboxInst_2_n5}), .clk (clk), .r (Fresh[170]), .c ({new_AGEMA_signal_1381, Feedback[9]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U7 ( .a ({new_AGEMA_signal_3240, new_AGEMA_signal_3238}), .b ({new_AGEMA_signal_1163, SubCellInst_SboxInst_2_n2}), .clk (clk), .r (Fresh[171]), .c ({new_AGEMA_signal_1305, SubCellInst_SboxInst_2_n3}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U19 ( .a ({new_AGEMA_signal_3248, new_AGEMA_signal_3246}), .b ({new_AGEMA_signal_1307, SubCellInst_SboxInst_3_n14}), .clk (clk), .r (Fresh[172]), .c ({new_AGEMA_signal_1383, Feedback[15]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U16 ( .a ({new_AGEMA_signal_1165, SubCellInst_SboxInst_3_n11}), .b ({new_AGEMA_signal_3252, new_AGEMA_signal_3250}), .clk (clk), .r (Fresh[173]), .c ({new_AGEMA_signal_1308, SubCellInst_SboxInst_3_n12}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U12 ( .a ({new_AGEMA_signal_3256, new_AGEMA_signal_3254}), .b ({new_AGEMA_signal_1309, SubCellInst_SboxInst_3_n5}), .clk (clk), .r (Fresh[174]), .c ({new_AGEMA_signal_1385, Feedback[13]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U7 ( .a ({new_AGEMA_signal_3252, new_AGEMA_signal_3250}), .b ({new_AGEMA_signal_1169, SubCellInst_SboxInst_3_n2}), .clk (clk), .r (Fresh[175]), .c ({new_AGEMA_signal_1310, SubCellInst_SboxInst_3_n3}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U19 ( .a ({new_AGEMA_signal_3260, new_AGEMA_signal_3258}), .b ({new_AGEMA_signal_1312, SubCellInst_SboxInst_4_n14}), .clk (clk), .r (Fresh[176]), .c ({new_AGEMA_signal_1387, Feedback[19]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U16 ( .a ({new_AGEMA_signal_1171, SubCellInst_SboxInst_4_n11}), .b ({new_AGEMA_signal_3264, new_AGEMA_signal_3262}), .clk (clk), .r (Fresh[177]), .c ({new_AGEMA_signal_1313, SubCellInst_SboxInst_4_n12}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U12 ( .a ({new_AGEMA_signal_3268, new_AGEMA_signal_3266}), .b ({new_AGEMA_signal_1314, SubCellInst_SboxInst_4_n5}), .clk (clk), .r (Fresh[178]), .c ({new_AGEMA_signal_1389, Feedback[17]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U7 ( .a ({new_AGEMA_signal_3264, new_AGEMA_signal_3262}), .b ({new_AGEMA_signal_1175, SubCellInst_SboxInst_4_n2}), .clk (clk), .r (Fresh[179]), .c ({new_AGEMA_signal_1315, SubCellInst_SboxInst_4_n3}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U19 ( .a ({new_AGEMA_signal_3272, new_AGEMA_signal_3270}), .b ({new_AGEMA_signal_1317, SubCellInst_SboxInst_5_n14}), .clk (clk), .r (Fresh[180]), .c ({new_AGEMA_signal_1391, Feedback[23]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U16 ( .a ({new_AGEMA_signal_1177, SubCellInst_SboxInst_5_n11}), .b ({new_AGEMA_signal_3276, new_AGEMA_signal_3274}), .clk (clk), .r (Fresh[181]), .c ({new_AGEMA_signal_1318, SubCellInst_SboxInst_5_n12}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U12 ( .a ({new_AGEMA_signal_3280, new_AGEMA_signal_3278}), .b ({new_AGEMA_signal_1319, SubCellInst_SboxInst_5_n5}), .clk (clk), .r (Fresh[182]), .c ({new_AGEMA_signal_1393, Feedback[21]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U7 ( .a ({new_AGEMA_signal_3276, new_AGEMA_signal_3274}), .b ({new_AGEMA_signal_1181, SubCellInst_SboxInst_5_n2}), .clk (clk), .r (Fresh[183]), .c ({new_AGEMA_signal_1320, SubCellInst_SboxInst_5_n3}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U19 ( .a ({new_AGEMA_signal_3284, new_AGEMA_signal_3282}), .b ({new_AGEMA_signal_1322, SubCellInst_SboxInst_6_n14}), .clk (clk), .r (Fresh[184]), .c ({new_AGEMA_signal_1395, Feedback[27]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U16 ( .a ({new_AGEMA_signal_1183, SubCellInst_SboxInst_6_n11}), .b ({new_AGEMA_signal_3288, new_AGEMA_signal_3286}), .clk (clk), .r (Fresh[185]), .c ({new_AGEMA_signal_1323, SubCellInst_SboxInst_6_n12}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U12 ( .a ({new_AGEMA_signal_3292, new_AGEMA_signal_3290}), .b ({new_AGEMA_signal_1324, SubCellInst_SboxInst_6_n5}), .clk (clk), .r (Fresh[186]), .c ({new_AGEMA_signal_1397, Feedback[25]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U7 ( .a ({new_AGEMA_signal_3288, new_AGEMA_signal_3286}), .b ({new_AGEMA_signal_1187, SubCellInst_SboxInst_6_n2}), .clk (clk), .r (Fresh[187]), .c ({new_AGEMA_signal_1325, SubCellInst_SboxInst_6_n3}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U19 ( .a ({new_AGEMA_signal_3296, new_AGEMA_signal_3294}), .b ({new_AGEMA_signal_1327, SubCellInst_SboxInst_7_n14}), .clk (clk), .r (Fresh[188]), .c ({new_AGEMA_signal_1399, Feedback[31]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U16 ( .a ({new_AGEMA_signal_1189, SubCellInst_SboxInst_7_n11}), .b ({new_AGEMA_signal_3300, new_AGEMA_signal_3298}), .clk (clk), .r (Fresh[189]), .c ({new_AGEMA_signal_1328, SubCellInst_SboxInst_7_n12}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U12 ( .a ({new_AGEMA_signal_3304, new_AGEMA_signal_3302}), .b ({new_AGEMA_signal_1329, SubCellInst_SboxInst_7_n5}), .clk (clk), .r (Fresh[190]), .c ({new_AGEMA_signal_1401, Feedback[29]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U7 ( .a ({new_AGEMA_signal_3300, new_AGEMA_signal_3298}), .b ({new_AGEMA_signal_1193, SubCellInst_SboxInst_7_n2}), .clk (clk), .r (Fresh[191]), .c ({new_AGEMA_signal_1330, SubCellInst_SboxInst_7_n3}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U19 ( .a ({new_AGEMA_signal_3308, new_AGEMA_signal_3306}), .b ({new_AGEMA_signal_1332, SubCellInst_SboxInst_8_n14}), .clk (clk), .r (Fresh[192]), .c ({new_AGEMA_signal_1403, Feedback[35]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U16 ( .a ({new_AGEMA_signal_1195, SubCellInst_SboxInst_8_n11}), .b ({new_AGEMA_signal_3312, new_AGEMA_signal_3310}), .clk (clk), .r (Fresh[193]), .c ({new_AGEMA_signal_1333, SubCellInst_SboxInst_8_n12}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U12 ( .a ({new_AGEMA_signal_3316, new_AGEMA_signal_3314}), .b ({new_AGEMA_signal_1334, SubCellInst_SboxInst_8_n5}), .clk (clk), .r (Fresh[194]), .c ({new_AGEMA_signal_1405, Feedback[33]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U7 ( .a ({new_AGEMA_signal_3312, new_AGEMA_signal_3310}), .b ({new_AGEMA_signal_1199, SubCellInst_SboxInst_8_n2}), .clk (clk), .r (Fresh[195]), .c ({new_AGEMA_signal_1335, SubCellInst_SboxInst_8_n3}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U19 ( .a ({new_AGEMA_signal_3320, new_AGEMA_signal_3318}), .b ({new_AGEMA_signal_1337, SubCellInst_SboxInst_9_n14}), .clk (clk), .r (Fresh[196]), .c ({new_AGEMA_signal_1407, Feedback[39]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U16 ( .a ({new_AGEMA_signal_1201, SubCellInst_SboxInst_9_n11}), .b ({new_AGEMA_signal_3324, new_AGEMA_signal_3322}), .clk (clk), .r (Fresh[197]), .c ({new_AGEMA_signal_1338, SubCellInst_SboxInst_9_n12}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U12 ( .a ({new_AGEMA_signal_3328, new_AGEMA_signal_3326}), .b ({new_AGEMA_signal_1339, SubCellInst_SboxInst_9_n5}), .clk (clk), .r (Fresh[198]), .c ({new_AGEMA_signal_1409, Feedback[37]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U7 ( .a ({new_AGEMA_signal_3324, new_AGEMA_signal_3322}), .b ({new_AGEMA_signal_1205, SubCellInst_SboxInst_9_n2}), .clk (clk), .r (Fresh[199]), .c ({new_AGEMA_signal_1340, SubCellInst_SboxInst_9_n3}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U19 ( .a ({new_AGEMA_signal_3332, new_AGEMA_signal_3330}), .b ({new_AGEMA_signal_1342, SubCellInst_SboxInst_10_n14}), .clk (clk), .r (Fresh[200]), .c ({new_AGEMA_signal_1411, Feedback[43]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U16 ( .a ({new_AGEMA_signal_1207, SubCellInst_SboxInst_10_n11}), .b ({new_AGEMA_signal_3336, new_AGEMA_signal_3334}), .clk (clk), .r (Fresh[201]), .c ({new_AGEMA_signal_1343, SubCellInst_SboxInst_10_n12}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U12 ( .a ({new_AGEMA_signal_3340, new_AGEMA_signal_3338}), .b ({new_AGEMA_signal_1344, SubCellInst_SboxInst_10_n5}), .clk (clk), .r (Fresh[202]), .c ({new_AGEMA_signal_1413, Feedback[41]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U7 ( .a ({new_AGEMA_signal_3336, new_AGEMA_signal_3334}), .b ({new_AGEMA_signal_1211, SubCellInst_SboxInst_10_n2}), .clk (clk), .r (Fresh[203]), .c ({new_AGEMA_signal_1345, SubCellInst_SboxInst_10_n3}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U19 ( .a ({new_AGEMA_signal_3344, new_AGEMA_signal_3342}), .b ({new_AGEMA_signal_1347, SubCellInst_SboxInst_11_n14}), .clk (clk), .r (Fresh[204]), .c ({new_AGEMA_signal_1415, Feedback[47]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U16 ( .a ({new_AGEMA_signal_1213, SubCellInst_SboxInst_11_n11}), .b ({new_AGEMA_signal_3348, new_AGEMA_signal_3346}), .clk (clk), .r (Fresh[205]), .c ({new_AGEMA_signal_1348, SubCellInst_SboxInst_11_n12}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U12 ( .a ({new_AGEMA_signal_3352, new_AGEMA_signal_3350}), .b ({new_AGEMA_signal_1349, SubCellInst_SboxInst_11_n5}), .clk (clk), .r (Fresh[206]), .c ({new_AGEMA_signal_1417, Feedback[45]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U7 ( .a ({new_AGEMA_signal_3348, new_AGEMA_signal_3346}), .b ({new_AGEMA_signal_1217, SubCellInst_SboxInst_11_n2}), .clk (clk), .r (Fresh[207]), .c ({new_AGEMA_signal_1350, SubCellInst_SboxInst_11_n3}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U19 ( .a ({new_AGEMA_signal_3356, new_AGEMA_signal_3354}), .b ({new_AGEMA_signal_1352, SubCellInst_SboxInst_12_n14}), .clk (clk), .r (Fresh[208]), .c ({new_AGEMA_signal_1419, Feedback[51]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U16 ( .a ({new_AGEMA_signal_1219, SubCellInst_SboxInst_12_n11}), .b ({new_AGEMA_signal_3360, new_AGEMA_signal_3358}), .clk (clk), .r (Fresh[209]), .c ({new_AGEMA_signal_1353, SubCellInst_SboxInst_12_n12}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U12 ( .a ({new_AGEMA_signal_3364, new_AGEMA_signal_3362}), .b ({new_AGEMA_signal_1354, SubCellInst_SboxInst_12_n5}), .clk (clk), .r (Fresh[210]), .c ({new_AGEMA_signal_1421, Feedback[49]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U7 ( .a ({new_AGEMA_signal_3360, new_AGEMA_signal_3358}), .b ({new_AGEMA_signal_1223, SubCellInst_SboxInst_12_n2}), .clk (clk), .r (Fresh[211]), .c ({new_AGEMA_signal_1355, SubCellInst_SboxInst_12_n3}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U19 ( .a ({new_AGEMA_signal_3368, new_AGEMA_signal_3366}), .b ({new_AGEMA_signal_1357, SubCellInst_SboxInst_13_n14}), .clk (clk), .r (Fresh[212]), .c ({new_AGEMA_signal_1423, Feedback[55]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U16 ( .a ({new_AGEMA_signal_1225, SubCellInst_SboxInst_13_n11}), .b ({new_AGEMA_signal_3372, new_AGEMA_signal_3370}), .clk (clk), .r (Fresh[213]), .c ({new_AGEMA_signal_1358, SubCellInst_SboxInst_13_n12}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U12 ( .a ({new_AGEMA_signal_3376, new_AGEMA_signal_3374}), .b ({new_AGEMA_signal_1359, SubCellInst_SboxInst_13_n5}), .clk (clk), .r (Fresh[214]), .c ({new_AGEMA_signal_1425, Feedback[53]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U7 ( .a ({new_AGEMA_signal_3372, new_AGEMA_signal_3370}), .b ({new_AGEMA_signal_1229, SubCellInst_SboxInst_13_n2}), .clk (clk), .r (Fresh[215]), .c ({new_AGEMA_signal_1360, SubCellInst_SboxInst_13_n3}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U19 ( .a ({new_AGEMA_signal_3380, new_AGEMA_signal_3378}), .b ({new_AGEMA_signal_1362, SubCellInst_SboxInst_14_n14}), .clk (clk), .r (Fresh[216]), .c ({new_AGEMA_signal_1427, Feedback[59]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U16 ( .a ({new_AGEMA_signal_1231, SubCellInst_SboxInst_14_n11}), .b ({new_AGEMA_signal_3384, new_AGEMA_signal_3382}), .clk (clk), .r (Fresh[217]), .c ({new_AGEMA_signal_1363, SubCellInst_SboxInst_14_n12}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U12 ( .a ({new_AGEMA_signal_3388, new_AGEMA_signal_3386}), .b ({new_AGEMA_signal_1364, SubCellInst_SboxInst_14_n5}), .clk (clk), .r (Fresh[218]), .c ({new_AGEMA_signal_1429, Feedback[57]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U7 ( .a ({new_AGEMA_signal_3384, new_AGEMA_signal_3382}), .b ({new_AGEMA_signal_1235, SubCellInst_SboxInst_14_n2}), .clk (clk), .r (Fresh[219]), .c ({new_AGEMA_signal_1365, SubCellInst_SboxInst_14_n3}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U19 ( .a ({new_AGEMA_signal_3392, new_AGEMA_signal_3390}), .b ({new_AGEMA_signal_1367, SubCellInst_SboxInst_15_n14}), .clk (clk), .r (Fresh[220]), .c ({new_AGEMA_signal_1431, Feedback[63]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U16 ( .a ({new_AGEMA_signal_1237, SubCellInst_SboxInst_15_n11}), .b ({new_AGEMA_signal_3396, new_AGEMA_signal_3394}), .clk (clk), .r (Fresh[221]), .c ({new_AGEMA_signal_1368, SubCellInst_SboxInst_15_n12}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U12 ( .a ({new_AGEMA_signal_3400, new_AGEMA_signal_3398}), .b ({new_AGEMA_signal_1369, SubCellInst_SboxInst_15_n5}), .clk (clk), .r (Fresh[222]), .c ({new_AGEMA_signal_1433, Feedback[61]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U7 ( .a ({new_AGEMA_signal_3396, new_AGEMA_signal_3394}), .b ({new_AGEMA_signal_1241, SubCellInst_SboxInst_15_n2}), .clk (clk), .r (Fresh[223]), .c ({new_AGEMA_signal_1370, SubCellInst_SboxInst_15_n3}) ) ;
    buf_clk new_AGEMA_reg_buffer_1080 ( .C (clk), .D (new_AGEMA_signal_2439), .Q (new_AGEMA_signal_2440) ) ;
    buf_clk new_AGEMA_reg_buffer_1086 ( .C (clk), .D (new_AGEMA_signal_2445), .Q (new_AGEMA_signal_2446) ) ;
    buf_clk new_AGEMA_reg_buffer_1092 ( .C (clk), .D (new_AGEMA_signal_2451), .Q (new_AGEMA_signal_2452) ) ;
    buf_clk new_AGEMA_reg_buffer_1098 ( .C (clk), .D (new_AGEMA_signal_2457), .Q (new_AGEMA_signal_2458) ) ;
    buf_clk new_AGEMA_reg_buffer_1104 ( .C (clk), .D (new_AGEMA_signal_2463), .Q (new_AGEMA_signal_2464) ) ;
    buf_clk new_AGEMA_reg_buffer_1110 ( .C (clk), .D (new_AGEMA_signal_2469), .Q (new_AGEMA_signal_2470) ) ;
    buf_clk new_AGEMA_reg_buffer_1116 ( .C (clk), .D (new_AGEMA_signal_2475), .Q (new_AGEMA_signal_2476) ) ;
    buf_clk new_AGEMA_reg_buffer_1122 ( .C (clk), .D (new_AGEMA_signal_2481), .Q (new_AGEMA_signal_2482) ) ;
    buf_clk new_AGEMA_reg_buffer_1128 ( .C (clk), .D (new_AGEMA_signal_2487), .Q (new_AGEMA_signal_2488) ) ;
    buf_clk new_AGEMA_reg_buffer_1134 ( .C (clk), .D (new_AGEMA_signal_2493), .Q (new_AGEMA_signal_2494) ) ;
    buf_clk new_AGEMA_reg_buffer_1140 ( .C (clk), .D (new_AGEMA_signal_2499), .Q (new_AGEMA_signal_2500) ) ;
    buf_clk new_AGEMA_reg_buffer_1146 ( .C (clk), .D (new_AGEMA_signal_2505), .Q (new_AGEMA_signal_2506) ) ;
    buf_clk new_AGEMA_reg_buffer_1152 ( .C (clk), .D (new_AGEMA_signal_2511), .Q (new_AGEMA_signal_2512) ) ;
    buf_clk new_AGEMA_reg_buffer_1158 ( .C (clk), .D (new_AGEMA_signal_2517), .Q (new_AGEMA_signal_2518) ) ;
    buf_clk new_AGEMA_reg_buffer_1164 ( .C (clk), .D (new_AGEMA_signal_2523), .Q (new_AGEMA_signal_2524) ) ;
    buf_clk new_AGEMA_reg_buffer_1170 ( .C (clk), .D (new_AGEMA_signal_2529), .Q (new_AGEMA_signal_2530) ) ;
    buf_clk new_AGEMA_reg_buffer_1176 ( .C (clk), .D (new_AGEMA_signal_2535), .Q (new_AGEMA_signal_2536) ) ;
    buf_clk new_AGEMA_reg_buffer_1182 ( .C (clk), .D (new_AGEMA_signal_2541), .Q (new_AGEMA_signal_2542) ) ;
    buf_clk new_AGEMA_reg_buffer_1188 ( .C (clk), .D (new_AGEMA_signal_2547), .Q (new_AGEMA_signal_2548) ) ;
    buf_clk new_AGEMA_reg_buffer_1194 ( .C (clk), .D (new_AGEMA_signal_2553), .Q (new_AGEMA_signal_2554) ) ;
    buf_clk new_AGEMA_reg_buffer_1200 ( .C (clk), .D (new_AGEMA_signal_2559), .Q (new_AGEMA_signal_2560) ) ;
    buf_clk new_AGEMA_reg_buffer_1206 ( .C (clk), .D (new_AGEMA_signal_2565), .Q (new_AGEMA_signal_2566) ) ;
    buf_clk new_AGEMA_reg_buffer_1212 ( .C (clk), .D (new_AGEMA_signal_2571), .Q (new_AGEMA_signal_2572) ) ;
    buf_clk new_AGEMA_reg_buffer_1218 ( .C (clk), .D (new_AGEMA_signal_2577), .Q (new_AGEMA_signal_2578) ) ;
    buf_clk new_AGEMA_reg_buffer_1224 ( .C (clk), .D (new_AGEMA_signal_2583), .Q (new_AGEMA_signal_2584) ) ;
    buf_clk new_AGEMA_reg_buffer_1230 ( .C (clk), .D (new_AGEMA_signal_2589), .Q (new_AGEMA_signal_2590) ) ;
    buf_clk new_AGEMA_reg_buffer_1236 ( .C (clk), .D (new_AGEMA_signal_2595), .Q (new_AGEMA_signal_2596) ) ;
    buf_clk new_AGEMA_reg_buffer_1242 ( .C (clk), .D (new_AGEMA_signal_2601), .Q (new_AGEMA_signal_2602) ) ;
    buf_clk new_AGEMA_reg_buffer_1248 ( .C (clk), .D (new_AGEMA_signal_2607), .Q (new_AGEMA_signal_2608) ) ;
    buf_clk new_AGEMA_reg_buffer_1254 ( .C (clk), .D (new_AGEMA_signal_2613), .Q (new_AGEMA_signal_2614) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C (clk), .D (new_AGEMA_signal_2619), .Q (new_AGEMA_signal_2620) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C (clk), .D (new_AGEMA_signal_2625), .Q (new_AGEMA_signal_2626) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C (clk), .D (new_AGEMA_signal_2631), .Q (new_AGEMA_signal_2632) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C (clk), .D (new_AGEMA_signal_2637), .Q (new_AGEMA_signal_2638) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C (clk), .D (new_AGEMA_signal_2643), .Q (new_AGEMA_signal_2644) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C (clk), .D (new_AGEMA_signal_2649), .Q (new_AGEMA_signal_2650) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C (clk), .D (new_AGEMA_signal_2655), .Q (new_AGEMA_signal_2656) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C (clk), .D (new_AGEMA_signal_2661), .Q (new_AGEMA_signal_2662) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C (clk), .D (new_AGEMA_signal_2667), .Q (new_AGEMA_signal_2668) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C (clk), .D (new_AGEMA_signal_2673), .Q (new_AGEMA_signal_2674) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C (clk), .D (new_AGEMA_signal_2679), .Q (new_AGEMA_signal_2680) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C (clk), .D (new_AGEMA_signal_2685), .Q (new_AGEMA_signal_2686) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C (clk), .D (new_AGEMA_signal_2691), .Q (new_AGEMA_signal_2692) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C (clk), .D (new_AGEMA_signal_2697), .Q (new_AGEMA_signal_2698) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C (clk), .D (new_AGEMA_signal_2703), .Q (new_AGEMA_signal_2704) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C (clk), .D (new_AGEMA_signal_2709), .Q (new_AGEMA_signal_2710) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C (clk), .D (new_AGEMA_signal_2715), .Q (new_AGEMA_signal_2716) ) ;
    buf_clk new_AGEMA_reg_buffer_1362 ( .C (clk), .D (new_AGEMA_signal_2721), .Q (new_AGEMA_signal_2722) ) ;
    buf_clk new_AGEMA_reg_buffer_1368 ( .C (clk), .D (new_AGEMA_signal_2727), .Q (new_AGEMA_signal_2728) ) ;
    buf_clk new_AGEMA_reg_buffer_1374 ( .C (clk), .D (new_AGEMA_signal_2733), .Q (new_AGEMA_signal_2734) ) ;
    buf_clk new_AGEMA_reg_buffer_1380 ( .C (clk), .D (new_AGEMA_signal_2739), .Q (new_AGEMA_signal_2740) ) ;
    buf_clk new_AGEMA_reg_buffer_1386 ( .C (clk), .D (new_AGEMA_signal_2745), .Q (new_AGEMA_signal_2746) ) ;
    buf_clk new_AGEMA_reg_buffer_1392 ( .C (clk), .D (new_AGEMA_signal_2751), .Q (new_AGEMA_signal_2752) ) ;
    buf_clk new_AGEMA_reg_buffer_1398 ( .C (clk), .D (new_AGEMA_signal_2757), .Q (new_AGEMA_signal_2758) ) ;
    buf_clk new_AGEMA_reg_buffer_1404 ( .C (clk), .D (new_AGEMA_signal_2763), .Q (new_AGEMA_signal_2764) ) ;
    buf_clk new_AGEMA_reg_buffer_1410 ( .C (clk), .D (new_AGEMA_signal_2769), .Q (new_AGEMA_signal_2770) ) ;
    buf_clk new_AGEMA_reg_buffer_1416 ( .C (clk), .D (new_AGEMA_signal_2775), .Q (new_AGEMA_signal_2776) ) ;
    buf_clk new_AGEMA_reg_buffer_1422 ( .C (clk), .D (new_AGEMA_signal_2781), .Q (new_AGEMA_signal_2782) ) ;
    buf_clk new_AGEMA_reg_buffer_1428 ( .C (clk), .D (new_AGEMA_signal_2787), .Q (new_AGEMA_signal_2788) ) ;
    buf_clk new_AGEMA_reg_buffer_1434 ( .C (clk), .D (new_AGEMA_signal_2793), .Q (new_AGEMA_signal_2794) ) ;
    buf_clk new_AGEMA_reg_buffer_1440 ( .C (clk), .D (new_AGEMA_signal_2799), .Q (new_AGEMA_signal_2800) ) ;
    buf_clk new_AGEMA_reg_buffer_1446 ( .C (clk), .D (new_AGEMA_signal_2805), .Q (new_AGEMA_signal_2806) ) ;
    buf_clk new_AGEMA_reg_buffer_1452 ( .C (clk), .D (new_AGEMA_signal_2811), .Q (new_AGEMA_signal_2812) ) ;
    buf_clk new_AGEMA_reg_buffer_1458 ( .C (clk), .D (new_AGEMA_signal_2817), .Q (new_AGEMA_signal_2818) ) ;
    buf_clk new_AGEMA_reg_buffer_1464 ( .C (clk), .D (new_AGEMA_signal_2823), .Q (new_AGEMA_signal_2824) ) ;
    buf_clk new_AGEMA_reg_buffer_1470 ( .C (clk), .D (new_AGEMA_signal_2829), .Q (new_AGEMA_signal_2830) ) ;
    buf_clk new_AGEMA_reg_buffer_1476 ( .C (clk), .D (new_AGEMA_signal_2835), .Q (new_AGEMA_signal_2836) ) ;
    buf_clk new_AGEMA_reg_buffer_1482 ( .C (clk), .D (new_AGEMA_signal_2841), .Q (new_AGEMA_signal_2842) ) ;
    buf_clk new_AGEMA_reg_buffer_1488 ( .C (clk), .D (new_AGEMA_signal_2847), .Q (new_AGEMA_signal_2848) ) ;
    buf_clk new_AGEMA_reg_buffer_1494 ( .C (clk), .D (new_AGEMA_signal_2853), .Q (new_AGEMA_signal_2854) ) ;
    buf_clk new_AGEMA_reg_buffer_1500 ( .C (clk), .D (new_AGEMA_signal_2859), .Q (new_AGEMA_signal_2860) ) ;
    buf_clk new_AGEMA_reg_buffer_1506 ( .C (clk), .D (new_AGEMA_signal_2865), .Q (new_AGEMA_signal_2866) ) ;
    buf_clk new_AGEMA_reg_buffer_1512 ( .C (clk), .D (new_AGEMA_signal_2871), .Q (new_AGEMA_signal_2872) ) ;
    buf_clk new_AGEMA_reg_buffer_1518 ( .C (clk), .D (new_AGEMA_signal_2877), .Q (new_AGEMA_signal_2878) ) ;
    buf_clk new_AGEMA_reg_buffer_1524 ( .C (clk), .D (new_AGEMA_signal_2883), .Q (new_AGEMA_signal_2884) ) ;
    buf_clk new_AGEMA_reg_buffer_1530 ( .C (clk), .D (new_AGEMA_signal_2889), .Q (new_AGEMA_signal_2890) ) ;
    buf_clk new_AGEMA_reg_buffer_1536 ( .C (clk), .D (new_AGEMA_signal_2895), .Q (new_AGEMA_signal_2896) ) ;
    buf_clk new_AGEMA_reg_buffer_1542 ( .C (clk), .D (new_AGEMA_signal_2901), .Q (new_AGEMA_signal_2902) ) ;
    buf_clk new_AGEMA_reg_buffer_1548 ( .C (clk), .D (new_AGEMA_signal_2907), .Q (new_AGEMA_signal_2908) ) ;
    buf_clk new_AGEMA_reg_buffer_1554 ( .C (clk), .D (new_AGEMA_signal_2913), .Q (new_AGEMA_signal_2914) ) ;
    buf_clk new_AGEMA_reg_buffer_1560 ( .C (clk), .D (new_AGEMA_signal_2919), .Q (new_AGEMA_signal_2920) ) ;
    buf_clk new_AGEMA_reg_buffer_1566 ( .C (clk), .D (new_AGEMA_signal_2925), .Q (new_AGEMA_signal_2926) ) ;
    buf_clk new_AGEMA_reg_buffer_1572 ( .C (clk), .D (new_AGEMA_signal_2931), .Q (new_AGEMA_signal_2932) ) ;
    buf_clk new_AGEMA_reg_buffer_1578 ( .C (clk), .D (new_AGEMA_signal_2937), .Q (new_AGEMA_signal_2938) ) ;
    buf_clk new_AGEMA_reg_buffer_1584 ( .C (clk), .D (new_AGEMA_signal_2943), .Q (new_AGEMA_signal_2944) ) ;
    buf_clk new_AGEMA_reg_buffer_1590 ( .C (clk), .D (new_AGEMA_signal_2949), .Q (new_AGEMA_signal_2950) ) ;
    buf_clk new_AGEMA_reg_buffer_1596 ( .C (clk), .D (new_AGEMA_signal_2955), .Q (new_AGEMA_signal_2956) ) ;
    buf_clk new_AGEMA_reg_buffer_1602 ( .C (clk), .D (new_AGEMA_signal_2961), .Q (new_AGEMA_signal_2962) ) ;
    buf_clk new_AGEMA_reg_buffer_1608 ( .C (clk), .D (new_AGEMA_signal_2967), .Q (new_AGEMA_signal_2968) ) ;
    buf_clk new_AGEMA_reg_buffer_1614 ( .C (clk), .D (new_AGEMA_signal_2973), .Q (new_AGEMA_signal_2974) ) ;
    buf_clk new_AGEMA_reg_buffer_1620 ( .C (clk), .D (new_AGEMA_signal_2979), .Q (new_AGEMA_signal_2980) ) ;
    buf_clk new_AGEMA_reg_buffer_1626 ( .C (clk), .D (new_AGEMA_signal_2985), .Q (new_AGEMA_signal_2986) ) ;
    buf_clk new_AGEMA_reg_buffer_1632 ( .C (clk), .D (new_AGEMA_signal_2991), .Q (new_AGEMA_signal_2992) ) ;
    buf_clk new_AGEMA_reg_buffer_1638 ( .C (clk), .D (new_AGEMA_signal_2997), .Q (new_AGEMA_signal_2998) ) ;
    buf_clk new_AGEMA_reg_buffer_1644 ( .C (clk), .D (new_AGEMA_signal_3003), .Q (new_AGEMA_signal_3004) ) ;
    buf_clk new_AGEMA_reg_buffer_1650 ( .C (clk), .D (new_AGEMA_signal_3009), .Q (new_AGEMA_signal_3010) ) ;
    buf_clk new_AGEMA_reg_buffer_1656 ( .C (clk), .D (new_AGEMA_signal_3015), .Q (new_AGEMA_signal_3016) ) ;
    buf_clk new_AGEMA_reg_buffer_1662 ( .C (clk), .D (new_AGEMA_signal_3021), .Q (new_AGEMA_signal_3022) ) ;
    buf_clk new_AGEMA_reg_buffer_1668 ( .C (clk), .D (new_AGEMA_signal_3027), .Q (new_AGEMA_signal_3028) ) ;
    buf_clk new_AGEMA_reg_buffer_1674 ( .C (clk), .D (new_AGEMA_signal_3033), .Q (new_AGEMA_signal_3034) ) ;
    buf_clk new_AGEMA_reg_buffer_1680 ( .C (clk), .D (new_AGEMA_signal_3039), .Q (new_AGEMA_signal_3040) ) ;
    buf_clk new_AGEMA_reg_buffer_1686 ( .C (clk), .D (new_AGEMA_signal_3045), .Q (new_AGEMA_signal_3046) ) ;
    buf_clk new_AGEMA_reg_buffer_1692 ( .C (clk), .D (new_AGEMA_signal_3051), .Q (new_AGEMA_signal_3052) ) ;
    buf_clk new_AGEMA_reg_buffer_1698 ( .C (clk), .D (new_AGEMA_signal_3057), .Q (new_AGEMA_signal_3058) ) ;
    buf_clk new_AGEMA_reg_buffer_1704 ( .C (clk), .D (new_AGEMA_signal_3063), .Q (new_AGEMA_signal_3064) ) ;
    buf_clk new_AGEMA_reg_buffer_1710 ( .C (clk), .D (new_AGEMA_signal_3069), .Q (new_AGEMA_signal_3070) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C (clk), .D (new_AGEMA_signal_3075), .Q (new_AGEMA_signal_3076) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C (clk), .D (new_AGEMA_signal_3081), .Q (new_AGEMA_signal_3082) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C (clk), .D (new_AGEMA_signal_3087), .Q (new_AGEMA_signal_3088) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C (clk), .D (new_AGEMA_signal_3093), .Q (new_AGEMA_signal_3094) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C (clk), .D (new_AGEMA_signal_3099), .Q (new_AGEMA_signal_3100) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C (clk), .D (new_AGEMA_signal_3105), .Q (new_AGEMA_signal_3106) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C (clk), .D (new_AGEMA_signal_3111), .Q (new_AGEMA_signal_3112) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C (clk), .D (new_AGEMA_signal_3117), .Q (new_AGEMA_signal_3118) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C (clk), .D (new_AGEMA_signal_3123), .Q (new_AGEMA_signal_3124) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C (clk), .D (new_AGEMA_signal_3129), .Q (new_AGEMA_signal_3130) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C (clk), .D (new_AGEMA_signal_3135), .Q (new_AGEMA_signal_3136) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C (clk), .D (new_AGEMA_signal_3141), .Q (new_AGEMA_signal_3142) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C (clk), .D (new_AGEMA_signal_3147), .Q (new_AGEMA_signal_3148) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C (clk), .D (new_AGEMA_signal_3153), .Q (new_AGEMA_signal_3154) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C (clk), .D (new_AGEMA_signal_3159), .Q (new_AGEMA_signal_3160) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C (clk), .D (new_AGEMA_signal_3165), .Q (new_AGEMA_signal_3166) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C (clk), .D (new_AGEMA_signal_3171), .Q (new_AGEMA_signal_3172) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C (clk), .D (new_AGEMA_signal_3177), .Q (new_AGEMA_signal_3178) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C (clk), .D (new_AGEMA_signal_3183), .Q (new_AGEMA_signal_3184) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C (clk), .D (new_AGEMA_signal_3189), .Q (new_AGEMA_signal_3190) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C (clk), .D (new_AGEMA_signal_3195), .Q (new_AGEMA_signal_3196) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C (clk), .D (new_AGEMA_signal_3201), .Q (new_AGEMA_signal_3202) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C (clk), .D (new_AGEMA_signal_3207), .Q (new_AGEMA_signal_3208) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C (clk), .D (new_AGEMA_signal_3407), .Q (new_AGEMA_signal_3408) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C (clk), .D (new_AGEMA_signal_3415), .Q (new_AGEMA_signal_3416) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C (clk), .D (new_AGEMA_signal_3423), .Q (new_AGEMA_signal_3424) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C (clk), .D (new_AGEMA_signal_3431), .Q (new_AGEMA_signal_3432) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C (clk), .D (new_AGEMA_signal_3439), .Q (new_AGEMA_signal_3440) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C (clk), .D (new_AGEMA_signal_3447), .Q (new_AGEMA_signal_3448) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C (clk), .D (new_AGEMA_signal_3455), .Q (new_AGEMA_signal_3456) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C (clk), .D (new_AGEMA_signal_3463), .Q (new_AGEMA_signal_3464) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C (clk), .D (new_AGEMA_signal_3471), .Q (new_AGEMA_signal_3472) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C (clk), .D (new_AGEMA_signal_3479), .Q (new_AGEMA_signal_3480) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C (clk), .D (new_AGEMA_signal_3487), .Q (new_AGEMA_signal_3488) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C (clk), .D (new_AGEMA_signal_3495), .Q (new_AGEMA_signal_3496) ) ;
    buf_clk new_AGEMA_reg_buffer_2144 ( .C (clk), .D (new_AGEMA_signal_3503), .Q (new_AGEMA_signal_3504) ) ;
    buf_clk new_AGEMA_reg_buffer_2152 ( .C (clk), .D (new_AGEMA_signal_3511), .Q (new_AGEMA_signal_3512) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C (clk), .D (new_AGEMA_signal_3519), .Q (new_AGEMA_signal_3520) ) ;
    buf_clk new_AGEMA_reg_buffer_2168 ( .C (clk), .D (new_AGEMA_signal_3527), .Q (new_AGEMA_signal_3528) ) ;
    buf_clk new_AGEMA_reg_buffer_2176 ( .C (clk), .D (new_AGEMA_signal_3535), .Q (new_AGEMA_signal_3536) ) ;
    buf_clk new_AGEMA_reg_buffer_2184 ( .C (clk), .D (new_AGEMA_signal_3543), .Q (new_AGEMA_signal_3544) ) ;
    buf_clk new_AGEMA_reg_buffer_2192 ( .C (clk), .D (new_AGEMA_signal_3551), .Q (new_AGEMA_signal_3552) ) ;
    buf_clk new_AGEMA_reg_buffer_2200 ( .C (clk), .D (new_AGEMA_signal_3559), .Q (new_AGEMA_signal_3560) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C (clk), .D (new_AGEMA_signal_3567), .Q (new_AGEMA_signal_3568) ) ;
    buf_clk new_AGEMA_reg_buffer_2216 ( .C (clk), .D (new_AGEMA_signal_3575), .Q (new_AGEMA_signal_3576) ) ;
    buf_clk new_AGEMA_reg_buffer_2224 ( .C (clk), .D (new_AGEMA_signal_3583), .Q (new_AGEMA_signal_3584) ) ;
    buf_clk new_AGEMA_reg_buffer_2232 ( .C (clk), .D (new_AGEMA_signal_3591), .Q (new_AGEMA_signal_3592) ) ;
    buf_clk new_AGEMA_reg_buffer_2240 ( .C (clk), .D (new_AGEMA_signal_3599), .Q (new_AGEMA_signal_3600) ) ;
    buf_clk new_AGEMA_reg_buffer_2248 ( .C (clk), .D (new_AGEMA_signal_3607), .Q (new_AGEMA_signal_3608) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C (clk), .D (new_AGEMA_signal_3615), .Q (new_AGEMA_signal_3616) ) ;
    buf_clk new_AGEMA_reg_buffer_2264 ( .C (clk), .D (new_AGEMA_signal_3623), .Q (new_AGEMA_signal_3624) ) ;
    buf_clk new_AGEMA_reg_buffer_2272 ( .C (clk), .D (new_AGEMA_signal_3631), .Q (new_AGEMA_signal_3632) ) ;
    buf_clk new_AGEMA_reg_buffer_2280 ( .C (clk), .D (new_AGEMA_signal_3639), .Q (new_AGEMA_signal_3640) ) ;
    buf_clk new_AGEMA_reg_buffer_2288 ( .C (clk), .D (new_AGEMA_signal_3647), .Q (new_AGEMA_signal_3648) ) ;
    buf_clk new_AGEMA_reg_buffer_2296 ( .C (clk), .D (new_AGEMA_signal_3655), .Q (new_AGEMA_signal_3656) ) ;
    buf_clk new_AGEMA_reg_buffer_2304 ( .C (clk), .D (new_AGEMA_signal_3663), .Q (new_AGEMA_signal_3664) ) ;
    buf_clk new_AGEMA_reg_buffer_2312 ( .C (clk), .D (new_AGEMA_signal_3671), .Q (new_AGEMA_signal_3672) ) ;
    buf_clk new_AGEMA_reg_buffer_2320 ( .C (clk), .D (new_AGEMA_signal_3679), .Q (new_AGEMA_signal_3680) ) ;
    buf_clk new_AGEMA_reg_buffer_2328 ( .C (clk), .D (new_AGEMA_signal_3687), .Q (new_AGEMA_signal_3688) ) ;
    buf_clk new_AGEMA_reg_buffer_2336 ( .C (clk), .D (new_AGEMA_signal_3695), .Q (new_AGEMA_signal_3696) ) ;
    buf_clk new_AGEMA_reg_buffer_2344 ( .C (clk), .D (new_AGEMA_signal_3703), .Q (new_AGEMA_signal_3704) ) ;
    buf_clk new_AGEMA_reg_buffer_2352 ( .C (clk), .D (new_AGEMA_signal_3711), .Q (new_AGEMA_signal_3712) ) ;
    buf_clk new_AGEMA_reg_buffer_2360 ( .C (clk), .D (new_AGEMA_signal_3719), .Q (new_AGEMA_signal_3720) ) ;
    buf_clk new_AGEMA_reg_buffer_2368 ( .C (clk), .D (new_AGEMA_signal_3727), .Q (new_AGEMA_signal_3728) ) ;
    buf_clk new_AGEMA_reg_buffer_2376 ( .C (clk), .D (new_AGEMA_signal_3735), .Q (new_AGEMA_signal_3736) ) ;
    buf_clk new_AGEMA_reg_buffer_2384 ( .C (clk), .D (new_AGEMA_signal_3743), .Q (new_AGEMA_signal_3744) ) ;
    buf_clk new_AGEMA_reg_buffer_2392 ( .C (clk), .D (new_AGEMA_signal_3751), .Q (new_AGEMA_signal_3752) ) ;
    buf_clk new_AGEMA_reg_buffer_2400 ( .C (clk), .D (new_AGEMA_signal_3759), .Q (new_AGEMA_signal_3760) ) ;
    buf_clk new_AGEMA_reg_buffer_2408 ( .C (clk), .D (new_AGEMA_signal_3767), .Q (new_AGEMA_signal_3768) ) ;
    buf_clk new_AGEMA_reg_buffer_2416 ( .C (clk), .D (new_AGEMA_signal_3775), .Q (new_AGEMA_signal_3776) ) ;
    buf_clk new_AGEMA_reg_buffer_2424 ( .C (clk), .D (new_AGEMA_signal_3783), .Q (new_AGEMA_signal_3784) ) ;
    buf_clk new_AGEMA_reg_buffer_2432 ( .C (clk), .D (new_AGEMA_signal_3791), .Q (new_AGEMA_signal_3792) ) ;
    buf_clk new_AGEMA_reg_buffer_2440 ( .C (clk), .D (new_AGEMA_signal_3799), .Q (new_AGEMA_signal_3800) ) ;
    buf_clk new_AGEMA_reg_buffer_2448 ( .C (clk), .D (new_AGEMA_signal_3807), .Q (new_AGEMA_signal_3808) ) ;
    buf_clk new_AGEMA_reg_buffer_2456 ( .C (clk), .D (new_AGEMA_signal_3815), .Q (new_AGEMA_signal_3816) ) ;
    buf_clk new_AGEMA_reg_buffer_2464 ( .C (clk), .D (new_AGEMA_signal_3823), .Q (new_AGEMA_signal_3824) ) ;
    buf_clk new_AGEMA_reg_buffer_2472 ( .C (clk), .D (new_AGEMA_signal_3831), .Q (new_AGEMA_signal_3832) ) ;
    buf_clk new_AGEMA_reg_buffer_2480 ( .C (clk), .D (new_AGEMA_signal_3839), .Q (new_AGEMA_signal_3840) ) ;
    buf_clk new_AGEMA_reg_buffer_2488 ( .C (clk), .D (new_AGEMA_signal_3847), .Q (new_AGEMA_signal_3848) ) ;
    buf_clk new_AGEMA_reg_buffer_2496 ( .C (clk), .D (new_AGEMA_signal_3855), .Q (new_AGEMA_signal_3856) ) ;
    buf_clk new_AGEMA_reg_buffer_2504 ( .C (clk), .D (new_AGEMA_signal_3863), .Q (new_AGEMA_signal_3864) ) ;
    buf_clk new_AGEMA_reg_buffer_2512 ( .C (clk), .D (new_AGEMA_signal_3871), .Q (new_AGEMA_signal_3872) ) ;
    buf_clk new_AGEMA_reg_buffer_2520 ( .C (clk), .D (new_AGEMA_signal_3879), .Q (new_AGEMA_signal_3880) ) ;
    buf_clk new_AGEMA_reg_buffer_2528 ( .C (clk), .D (new_AGEMA_signal_3887), .Q (new_AGEMA_signal_3888) ) ;
    buf_clk new_AGEMA_reg_buffer_2536 ( .C (clk), .D (new_AGEMA_signal_3895), .Q (new_AGEMA_signal_3896) ) ;
    buf_clk new_AGEMA_reg_buffer_2544 ( .C (clk), .D (new_AGEMA_signal_3903), .Q (new_AGEMA_signal_3904) ) ;
    buf_clk new_AGEMA_reg_buffer_2552 ( .C (clk), .D (new_AGEMA_signal_3911), .Q (new_AGEMA_signal_3912) ) ;
    buf_clk new_AGEMA_reg_buffer_2560 ( .C (clk), .D (new_AGEMA_signal_3919), .Q (new_AGEMA_signal_3920) ) ;
    buf_clk new_AGEMA_reg_buffer_2568 ( .C (clk), .D (new_AGEMA_signal_3927), .Q (new_AGEMA_signal_3928) ) ;
    buf_clk new_AGEMA_reg_buffer_2576 ( .C (clk), .D (new_AGEMA_signal_3935), .Q (new_AGEMA_signal_3936) ) ;
    buf_clk new_AGEMA_reg_buffer_2584 ( .C (clk), .D (new_AGEMA_signal_3943), .Q (new_AGEMA_signal_3944) ) ;
    buf_clk new_AGEMA_reg_buffer_2592 ( .C (clk), .D (new_AGEMA_signal_3951), .Q (new_AGEMA_signal_3952) ) ;
    buf_clk new_AGEMA_reg_buffer_2600 ( .C (clk), .D (new_AGEMA_signal_3959), .Q (new_AGEMA_signal_3960) ) ;
    buf_clk new_AGEMA_reg_buffer_2608 ( .C (clk), .D (new_AGEMA_signal_3967), .Q (new_AGEMA_signal_3968) ) ;
    buf_clk new_AGEMA_reg_buffer_2616 ( .C (clk), .D (new_AGEMA_signal_3975), .Q (new_AGEMA_signal_3976) ) ;
    buf_clk new_AGEMA_reg_buffer_2624 ( .C (clk), .D (new_AGEMA_signal_3983), .Q (new_AGEMA_signal_3984) ) ;
    buf_clk new_AGEMA_reg_buffer_2632 ( .C (clk), .D (new_AGEMA_signal_3991), .Q (new_AGEMA_signal_3992) ) ;
    buf_clk new_AGEMA_reg_buffer_2640 ( .C (clk), .D (new_AGEMA_signal_3999), .Q (new_AGEMA_signal_4000) ) ;
    buf_clk new_AGEMA_reg_buffer_2648 ( .C (clk), .D (new_AGEMA_signal_4007), .Q (new_AGEMA_signal_4008) ) ;
    buf_clk new_AGEMA_reg_buffer_2656 ( .C (clk), .D (new_AGEMA_signal_4015), .Q (new_AGEMA_signal_4016) ) ;
    buf_clk new_AGEMA_reg_buffer_2664 ( .C (clk), .D (new_AGEMA_signal_4023), .Q (new_AGEMA_signal_4024) ) ;
    buf_clk new_AGEMA_reg_buffer_2672 ( .C (clk), .D (new_AGEMA_signal_4031), .Q (new_AGEMA_signal_4032) ) ;
    buf_clk new_AGEMA_reg_buffer_2680 ( .C (clk), .D (new_AGEMA_signal_4039), .Q (new_AGEMA_signal_4040) ) ;
    buf_clk new_AGEMA_reg_buffer_2688 ( .C (clk), .D (new_AGEMA_signal_4047), .Q (new_AGEMA_signal_4048) ) ;
    buf_clk new_AGEMA_reg_buffer_2696 ( .C (clk), .D (new_AGEMA_signal_4055), .Q (new_AGEMA_signal_4056) ) ;
    buf_clk new_AGEMA_reg_buffer_2704 ( .C (clk), .D (new_AGEMA_signal_4063), .Q (new_AGEMA_signal_4064) ) ;
    buf_clk new_AGEMA_reg_buffer_2712 ( .C (clk), .D (new_AGEMA_signal_4071), .Q (new_AGEMA_signal_4072) ) ;
    buf_clk new_AGEMA_reg_buffer_2720 ( .C (clk), .D (new_AGEMA_signal_4079), .Q (new_AGEMA_signal_4080) ) ;
    buf_clk new_AGEMA_reg_buffer_2728 ( .C (clk), .D (new_AGEMA_signal_4087), .Q (new_AGEMA_signal_4088) ) ;
    buf_clk new_AGEMA_reg_buffer_2736 ( .C (clk), .D (new_AGEMA_signal_4095), .Q (new_AGEMA_signal_4096) ) ;
    buf_clk new_AGEMA_reg_buffer_2744 ( .C (clk), .D (new_AGEMA_signal_4103), .Q (new_AGEMA_signal_4104) ) ;
    buf_clk new_AGEMA_reg_buffer_2752 ( .C (clk), .D (new_AGEMA_signal_4111), .Q (new_AGEMA_signal_4112) ) ;
    buf_clk new_AGEMA_reg_buffer_2760 ( .C (clk), .D (new_AGEMA_signal_4119), .Q (new_AGEMA_signal_4120) ) ;
    buf_clk new_AGEMA_reg_buffer_2768 ( .C (clk), .D (new_AGEMA_signal_4127), .Q (new_AGEMA_signal_4128) ) ;
    buf_clk new_AGEMA_reg_buffer_2776 ( .C (clk), .D (new_AGEMA_signal_4135), .Q (new_AGEMA_signal_4136) ) ;
    buf_clk new_AGEMA_reg_buffer_2784 ( .C (clk), .D (new_AGEMA_signal_4143), .Q (new_AGEMA_signal_4144) ) ;
    buf_clk new_AGEMA_reg_buffer_2792 ( .C (clk), .D (new_AGEMA_signal_4151), .Q (new_AGEMA_signal_4152) ) ;
    buf_clk new_AGEMA_reg_buffer_2800 ( .C (clk), .D (new_AGEMA_signal_4159), .Q (new_AGEMA_signal_4160) ) ;
    buf_clk new_AGEMA_reg_buffer_2808 ( .C (clk), .D (new_AGEMA_signal_4167), .Q (new_AGEMA_signal_4168) ) ;
    buf_clk new_AGEMA_reg_buffer_2816 ( .C (clk), .D (new_AGEMA_signal_4175), .Q (new_AGEMA_signal_4176) ) ;
    buf_clk new_AGEMA_reg_buffer_2824 ( .C (clk), .D (new_AGEMA_signal_4183), .Q (new_AGEMA_signal_4184) ) ;
    buf_clk new_AGEMA_reg_buffer_2832 ( .C (clk), .D (new_AGEMA_signal_4191), .Q (new_AGEMA_signal_4192) ) ;
    buf_clk new_AGEMA_reg_buffer_2840 ( .C (clk), .D (new_AGEMA_signal_4199), .Q (new_AGEMA_signal_4200) ) ;
    buf_clk new_AGEMA_reg_buffer_2848 ( .C (clk), .D (new_AGEMA_signal_4207), .Q (new_AGEMA_signal_4208) ) ;
    buf_clk new_AGEMA_reg_buffer_2856 ( .C (clk), .D (new_AGEMA_signal_4215), .Q (new_AGEMA_signal_4216) ) ;
    buf_clk new_AGEMA_reg_buffer_2864 ( .C (clk), .D (new_AGEMA_signal_4223), .Q (new_AGEMA_signal_4224) ) ;
    buf_clk new_AGEMA_reg_buffer_2872 ( .C (clk), .D (new_AGEMA_signal_4231), .Q (new_AGEMA_signal_4232) ) ;
    buf_clk new_AGEMA_reg_buffer_2880 ( .C (clk), .D (new_AGEMA_signal_4239), .Q (new_AGEMA_signal_4240) ) ;
    buf_clk new_AGEMA_reg_buffer_2888 ( .C (clk), .D (new_AGEMA_signal_4247), .Q (new_AGEMA_signal_4248) ) ;
    buf_clk new_AGEMA_reg_buffer_2896 ( .C (clk), .D (new_AGEMA_signal_4255), .Q (new_AGEMA_signal_4256) ) ;
    buf_clk new_AGEMA_reg_buffer_2904 ( .C (clk), .D (new_AGEMA_signal_4263), .Q (new_AGEMA_signal_4264) ) ;
    buf_clk new_AGEMA_reg_buffer_2912 ( .C (clk), .D (new_AGEMA_signal_4271), .Q (new_AGEMA_signal_4272) ) ;
    buf_clk new_AGEMA_reg_buffer_2920 ( .C (clk), .D (new_AGEMA_signal_4279), .Q (new_AGEMA_signal_4280) ) ;
    buf_clk new_AGEMA_reg_buffer_2928 ( .C (clk), .D (new_AGEMA_signal_4287), .Q (new_AGEMA_signal_4288) ) ;
    buf_clk new_AGEMA_reg_buffer_2936 ( .C (clk), .D (new_AGEMA_signal_4295), .Q (new_AGEMA_signal_4296) ) ;
    buf_clk new_AGEMA_reg_buffer_2944 ( .C (clk), .D (new_AGEMA_signal_4303), .Q (new_AGEMA_signal_4304) ) ;
    buf_clk new_AGEMA_reg_buffer_2952 ( .C (clk), .D (new_AGEMA_signal_4311), .Q (new_AGEMA_signal_4312) ) ;
    buf_clk new_AGEMA_reg_buffer_2960 ( .C (clk), .D (new_AGEMA_signal_4319), .Q (new_AGEMA_signal_4320) ) ;
    buf_clk new_AGEMA_reg_buffer_2968 ( .C (clk), .D (new_AGEMA_signal_4327), .Q (new_AGEMA_signal_4328) ) ;
    buf_clk new_AGEMA_reg_buffer_2976 ( .C (clk), .D (new_AGEMA_signal_4335), .Q (new_AGEMA_signal_4336) ) ;
    buf_clk new_AGEMA_reg_buffer_2984 ( .C (clk), .D (new_AGEMA_signal_4343), .Q (new_AGEMA_signal_4344) ) ;
    buf_clk new_AGEMA_reg_buffer_2992 ( .C (clk), .D (new_AGEMA_signal_4351), .Q (new_AGEMA_signal_4352) ) ;
    buf_clk new_AGEMA_reg_buffer_3000 ( .C (clk), .D (new_AGEMA_signal_4359), .Q (new_AGEMA_signal_4360) ) ;
    buf_clk new_AGEMA_reg_buffer_3008 ( .C (clk), .D (new_AGEMA_signal_4367), .Q (new_AGEMA_signal_4368) ) ;
    buf_clk new_AGEMA_reg_buffer_3016 ( .C (clk), .D (new_AGEMA_signal_4375), .Q (new_AGEMA_signal_4376) ) ;
    buf_clk new_AGEMA_reg_buffer_3024 ( .C (clk), .D (new_AGEMA_signal_4383), .Q (new_AGEMA_signal_4384) ) ;
    buf_clk new_AGEMA_reg_buffer_3032 ( .C (clk), .D (new_AGEMA_signal_4391), .Q (new_AGEMA_signal_4392) ) ;
    buf_clk new_AGEMA_reg_buffer_3040 ( .C (clk), .D (new_AGEMA_signal_4399), .Q (new_AGEMA_signal_4400) ) ;
    buf_clk new_AGEMA_reg_buffer_3048 ( .C (clk), .D (new_AGEMA_signal_4407), .Q (new_AGEMA_signal_4408) ) ;
    buf_clk new_AGEMA_reg_buffer_3056 ( .C (clk), .D (new_AGEMA_signal_4415), .Q (new_AGEMA_signal_4416) ) ;
    buf_clk new_AGEMA_reg_buffer_3064 ( .C (clk), .D (new_AGEMA_signal_4423), .Q (new_AGEMA_signal_4424) ) ;
    buf_clk new_AGEMA_reg_buffer_3068 ( .C (clk), .D (new_AGEMA_signal_4427), .Q (new_AGEMA_signal_4428) ) ;
    buf_clk new_AGEMA_reg_buffer_3070 ( .C (clk), .D (new_AGEMA_signal_4429), .Q (new_AGEMA_signal_4430) ) ;
    buf_clk new_AGEMA_reg_buffer_3074 ( .C (clk), .D (new_AGEMA_signal_4433), .Q (new_AGEMA_signal_4434) ) ;
    buf_clk new_AGEMA_reg_buffer_3078 ( .C (clk), .D (new_AGEMA_signal_4437), .Q (new_AGEMA_signal_4438) ) ;
    buf_clk new_AGEMA_reg_buffer_3080 ( .C (clk), .D (new_AGEMA_signal_4439), .Q (new_AGEMA_signal_4440) ) ;
    buf_clk new_AGEMA_reg_buffer_3082 ( .C (clk), .D (new_AGEMA_signal_4441), .Q (new_AGEMA_signal_4442) ) ;
    buf_clk new_AGEMA_reg_buffer_3086 ( .C (clk), .D (new_AGEMA_signal_4445), .Q (new_AGEMA_signal_4446) ) ;
    buf_clk new_AGEMA_reg_buffer_3090 ( .C (clk), .D (new_AGEMA_signal_4449), .Q (new_AGEMA_signal_4450) ) ;
    buf_clk new_AGEMA_reg_buffer_3092 ( .C (clk), .D (new_AGEMA_signal_4451), .Q (new_AGEMA_signal_4452) ) ;
    buf_clk new_AGEMA_reg_buffer_3094 ( .C (clk), .D (new_AGEMA_signal_4453), .Q (new_AGEMA_signal_4454) ) ;
    buf_clk new_AGEMA_reg_buffer_3098 ( .C (clk), .D (new_AGEMA_signal_4457), .Q (new_AGEMA_signal_4458) ) ;
    buf_clk new_AGEMA_reg_buffer_3102 ( .C (clk), .D (new_AGEMA_signal_4461), .Q (new_AGEMA_signal_4462) ) ;
    buf_clk new_AGEMA_reg_buffer_3104 ( .C (clk), .D (new_AGEMA_signal_4463), .Q (new_AGEMA_signal_4464) ) ;
    buf_clk new_AGEMA_reg_buffer_3106 ( .C (clk), .D (new_AGEMA_signal_4465), .Q (new_AGEMA_signal_4466) ) ;
    buf_clk new_AGEMA_reg_buffer_3110 ( .C (clk), .D (new_AGEMA_signal_4469), .Q (new_AGEMA_signal_4470) ) ;
    buf_clk new_AGEMA_reg_buffer_3114 ( .C (clk), .D (new_AGEMA_signal_4473), .Q (new_AGEMA_signal_4474) ) ;
    buf_clk new_AGEMA_reg_buffer_3116 ( .C (clk), .D (new_AGEMA_signal_4475), .Q (new_AGEMA_signal_4476) ) ;
    buf_clk new_AGEMA_reg_buffer_3118 ( .C (clk), .D (new_AGEMA_signal_4477), .Q (new_AGEMA_signal_4478) ) ;
    buf_clk new_AGEMA_reg_buffer_3122 ( .C (clk), .D (new_AGEMA_signal_4481), .Q (new_AGEMA_signal_4482) ) ;
    buf_clk new_AGEMA_reg_buffer_3126 ( .C (clk), .D (new_AGEMA_signal_4485), .Q (new_AGEMA_signal_4486) ) ;
    buf_clk new_AGEMA_reg_buffer_3128 ( .C (clk), .D (new_AGEMA_signal_4487), .Q (new_AGEMA_signal_4488) ) ;
    buf_clk new_AGEMA_reg_buffer_3130 ( .C (clk), .D (new_AGEMA_signal_4489), .Q (new_AGEMA_signal_4490) ) ;
    buf_clk new_AGEMA_reg_buffer_3134 ( .C (clk), .D (new_AGEMA_signal_4493), .Q (new_AGEMA_signal_4494) ) ;
    buf_clk new_AGEMA_reg_buffer_3138 ( .C (clk), .D (new_AGEMA_signal_4497), .Q (new_AGEMA_signal_4498) ) ;
    buf_clk new_AGEMA_reg_buffer_3140 ( .C (clk), .D (new_AGEMA_signal_4499), .Q (new_AGEMA_signal_4500) ) ;
    buf_clk new_AGEMA_reg_buffer_3142 ( .C (clk), .D (new_AGEMA_signal_4501), .Q (new_AGEMA_signal_4502) ) ;
    buf_clk new_AGEMA_reg_buffer_3146 ( .C (clk), .D (new_AGEMA_signal_4505), .Q (new_AGEMA_signal_4506) ) ;
    buf_clk new_AGEMA_reg_buffer_3150 ( .C (clk), .D (new_AGEMA_signal_4509), .Q (new_AGEMA_signal_4510) ) ;
    buf_clk new_AGEMA_reg_buffer_3152 ( .C (clk), .D (new_AGEMA_signal_4511), .Q (new_AGEMA_signal_4512) ) ;
    buf_clk new_AGEMA_reg_buffer_3154 ( .C (clk), .D (new_AGEMA_signal_4513), .Q (new_AGEMA_signal_4514) ) ;
    buf_clk new_AGEMA_reg_buffer_3158 ( .C (clk), .D (new_AGEMA_signal_4517), .Q (new_AGEMA_signal_4518) ) ;
    buf_clk new_AGEMA_reg_buffer_3162 ( .C (clk), .D (new_AGEMA_signal_4521), .Q (new_AGEMA_signal_4522) ) ;
    buf_clk new_AGEMA_reg_buffer_3164 ( .C (clk), .D (new_AGEMA_signal_4523), .Q (new_AGEMA_signal_4524) ) ;
    buf_clk new_AGEMA_reg_buffer_3166 ( .C (clk), .D (new_AGEMA_signal_4525), .Q (new_AGEMA_signal_4526) ) ;
    buf_clk new_AGEMA_reg_buffer_3170 ( .C (clk), .D (new_AGEMA_signal_4529), .Q (new_AGEMA_signal_4530) ) ;
    buf_clk new_AGEMA_reg_buffer_3174 ( .C (clk), .D (new_AGEMA_signal_4533), .Q (new_AGEMA_signal_4534) ) ;
    buf_clk new_AGEMA_reg_buffer_3176 ( .C (clk), .D (new_AGEMA_signal_4535), .Q (new_AGEMA_signal_4536) ) ;
    buf_clk new_AGEMA_reg_buffer_3178 ( .C (clk), .D (new_AGEMA_signal_4537), .Q (new_AGEMA_signal_4538) ) ;
    buf_clk new_AGEMA_reg_buffer_3182 ( .C (clk), .D (new_AGEMA_signal_4541), .Q (new_AGEMA_signal_4542) ) ;
    buf_clk new_AGEMA_reg_buffer_3186 ( .C (clk), .D (new_AGEMA_signal_4545), .Q (new_AGEMA_signal_4546) ) ;
    buf_clk new_AGEMA_reg_buffer_3188 ( .C (clk), .D (new_AGEMA_signal_4547), .Q (new_AGEMA_signal_4548) ) ;
    buf_clk new_AGEMA_reg_buffer_3190 ( .C (clk), .D (new_AGEMA_signal_4549), .Q (new_AGEMA_signal_4550) ) ;
    buf_clk new_AGEMA_reg_buffer_3194 ( .C (clk), .D (new_AGEMA_signal_4553), .Q (new_AGEMA_signal_4554) ) ;
    buf_clk new_AGEMA_reg_buffer_3198 ( .C (clk), .D (new_AGEMA_signal_4557), .Q (new_AGEMA_signal_4558) ) ;
    buf_clk new_AGEMA_reg_buffer_3200 ( .C (clk), .D (new_AGEMA_signal_4559), .Q (new_AGEMA_signal_4560) ) ;
    buf_clk new_AGEMA_reg_buffer_3202 ( .C (clk), .D (new_AGEMA_signal_4561), .Q (new_AGEMA_signal_4562) ) ;
    buf_clk new_AGEMA_reg_buffer_3206 ( .C (clk), .D (new_AGEMA_signal_4565), .Q (new_AGEMA_signal_4566) ) ;
    buf_clk new_AGEMA_reg_buffer_3210 ( .C (clk), .D (new_AGEMA_signal_4569), .Q (new_AGEMA_signal_4570) ) ;
    buf_clk new_AGEMA_reg_buffer_3212 ( .C (clk), .D (new_AGEMA_signal_4571), .Q (new_AGEMA_signal_4572) ) ;
    buf_clk new_AGEMA_reg_buffer_3214 ( .C (clk), .D (new_AGEMA_signal_4573), .Q (new_AGEMA_signal_4574) ) ;
    buf_clk new_AGEMA_reg_buffer_3218 ( .C (clk), .D (new_AGEMA_signal_4577), .Q (new_AGEMA_signal_4578) ) ;
    buf_clk new_AGEMA_reg_buffer_3222 ( .C (clk), .D (new_AGEMA_signal_4581), .Q (new_AGEMA_signal_4582) ) ;
    buf_clk new_AGEMA_reg_buffer_3224 ( .C (clk), .D (new_AGEMA_signal_4583), .Q (new_AGEMA_signal_4584) ) ;
    buf_clk new_AGEMA_reg_buffer_3226 ( .C (clk), .D (new_AGEMA_signal_4585), .Q (new_AGEMA_signal_4586) ) ;
    buf_clk new_AGEMA_reg_buffer_3230 ( .C (clk), .D (new_AGEMA_signal_4589), .Q (new_AGEMA_signal_4590) ) ;
    buf_clk new_AGEMA_reg_buffer_3234 ( .C (clk), .D (new_AGEMA_signal_4593), .Q (new_AGEMA_signal_4594) ) ;
    buf_clk new_AGEMA_reg_buffer_3236 ( .C (clk), .D (new_AGEMA_signal_4595), .Q (new_AGEMA_signal_4596) ) ;
    buf_clk new_AGEMA_reg_buffer_3238 ( .C (clk), .D (new_AGEMA_signal_4597), .Q (new_AGEMA_signal_4598) ) ;
    buf_clk new_AGEMA_reg_buffer_3242 ( .C (clk), .D (new_AGEMA_signal_4601), .Q (new_AGEMA_signal_4602) ) ;
    buf_clk new_AGEMA_reg_buffer_3246 ( .C (clk), .D (new_AGEMA_signal_4605), .Q (new_AGEMA_signal_4606) ) ;
    buf_clk new_AGEMA_reg_buffer_3248 ( .C (clk), .D (new_AGEMA_signal_4607), .Q (new_AGEMA_signal_4608) ) ;
    buf_clk new_AGEMA_reg_buffer_3250 ( .C (clk), .D (new_AGEMA_signal_4609), .Q (new_AGEMA_signal_4610) ) ;
    buf_clk new_AGEMA_reg_buffer_3254 ( .C (clk), .D (new_AGEMA_signal_4613), .Q (new_AGEMA_signal_4614) ) ;
    buf_clk new_AGEMA_reg_buffer_3258 ( .C (clk), .D (new_AGEMA_signal_4617), .Q (new_AGEMA_signal_4618) ) ;
    buf_clk new_AGEMA_reg_buffer_3392 ( .C (clk), .D (new_AGEMA_signal_4751), .Q (new_AGEMA_signal_4752) ) ;
    buf_clk new_AGEMA_reg_buffer_3400 ( .C (clk), .D (new_AGEMA_signal_4759), .Q (new_AGEMA_signal_4760) ) ;
    buf_clk new_AGEMA_reg_buffer_3408 ( .C (clk), .D (new_AGEMA_signal_4767), .Q (new_AGEMA_signal_4768) ) ;
    buf_clk new_AGEMA_reg_buffer_3416 ( .C (clk), .D (new_AGEMA_signal_4775), .Q (new_AGEMA_signal_4776) ) ;
    buf_clk new_AGEMA_reg_buffer_3424 ( .C (clk), .D (new_AGEMA_signal_4783), .Q (new_AGEMA_signal_4784) ) ;
    buf_clk new_AGEMA_reg_buffer_3432 ( .C (clk), .D (new_AGEMA_signal_4791), .Q (new_AGEMA_signal_4792) ) ;
    buf_clk new_AGEMA_reg_buffer_3440 ( .C (clk), .D (new_AGEMA_signal_4799), .Q (new_AGEMA_signal_4800) ) ;
    buf_clk new_AGEMA_reg_buffer_3448 ( .C (clk), .D (new_AGEMA_signal_4807), .Q (new_AGEMA_signal_4808) ) ;
    buf_clk new_AGEMA_reg_buffer_3456 ( .C (clk), .D (new_AGEMA_signal_4815), .Q (new_AGEMA_signal_4816) ) ;
    buf_clk new_AGEMA_reg_buffer_3464 ( .C (clk), .D (new_AGEMA_signal_4823), .Q (new_AGEMA_signal_4824) ) ;

    /* cells in depth 7 */
    buf_clk new_AGEMA_reg_buffer_2041 ( .C (clk), .D (new_AGEMA_signal_2440), .Q (new_AGEMA_signal_3401) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C (clk), .D (new_AGEMA_signal_3408), .Q (new_AGEMA_signal_3409) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C (clk), .D (new_AGEMA_signal_3416), .Q (new_AGEMA_signal_3417) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C (clk), .D (new_AGEMA_signal_3424), .Q (new_AGEMA_signal_3425) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C (clk), .D (new_AGEMA_signal_3432), .Q (new_AGEMA_signal_3433) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C (clk), .D (new_AGEMA_signal_3440), .Q (new_AGEMA_signal_3441) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C (clk), .D (new_AGEMA_signal_3448), .Q (new_AGEMA_signal_3449) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C (clk), .D (new_AGEMA_signal_3456), .Q (new_AGEMA_signal_3457) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C (clk), .D (new_AGEMA_signal_3464), .Q (new_AGEMA_signal_3465) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C (clk), .D (new_AGEMA_signal_3472), .Q (new_AGEMA_signal_3473) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C (clk), .D (new_AGEMA_signal_3480), .Q (new_AGEMA_signal_3481) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C (clk), .D (new_AGEMA_signal_3488), .Q (new_AGEMA_signal_3489) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C (clk), .D (new_AGEMA_signal_3496), .Q (new_AGEMA_signal_3497) ) ;
    buf_clk new_AGEMA_reg_buffer_2145 ( .C (clk), .D (new_AGEMA_signal_3504), .Q (new_AGEMA_signal_3505) ) ;
    buf_clk new_AGEMA_reg_buffer_2153 ( .C (clk), .D (new_AGEMA_signal_3512), .Q (new_AGEMA_signal_3513) ) ;
    buf_clk new_AGEMA_reg_buffer_2161 ( .C (clk), .D (new_AGEMA_signal_3520), .Q (new_AGEMA_signal_3521) ) ;
    buf_clk new_AGEMA_reg_buffer_2169 ( .C (clk), .D (new_AGEMA_signal_3528), .Q (new_AGEMA_signal_3529) ) ;
    buf_clk new_AGEMA_reg_buffer_2177 ( .C (clk), .D (new_AGEMA_signal_3536), .Q (new_AGEMA_signal_3537) ) ;
    buf_clk new_AGEMA_reg_buffer_2185 ( .C (clk), .D (new_AGEMA_signal_3544), .Q (new_AGEMA_signal_3545) ) ;
    buf_clk new_AGEMA_reg_buffer_2193 ( .C (clk), .D (new_AGEMA_signal_3552), .Q (new_AGEMA_signal_3553) ) ;
    buf_clk new_AGEMA_reg_buffer_2201 ( .C (clk), .D (new_AGEMA_signal_3560), .Q (new_AGEMA_signal_3561) ) ;
    buf_clk new_AGEMA_reg_buffer_2209 ( .C (clk), .D (new_AGEMA_signal_3568), .Q (new_AGEMA_signal_3569) ) ;
    buf_clk new_AGEMA_reg_buffer_2217 ( .C (clk), .D (new_AGEMA_signal_3576), .Q (new_AGEMA_signal_3577) ) ;
    buf_clk new_AGEMA_reg_buffer_2225 ( .C (clk), .D (new_AGEMA_signal_3584), .Q (new_AGEMA_signal_3585) ) ;
    buf_clk new_AGEMA_reg_buffer_2233 ( .C (clk), .D (new_AGEMA_signal_3592), .Q (new_AGEMA_signal_3593) ) ;
    buf_clk new_AGEMA_reg_buffer_2241 ( .C (clk), .D (new_AGEMA_signal_3600), .Q (new_AGEMA_signal_3601) ) ;
    buf_clk new_AGEMA_reg_buffer_2249 ( .C (clk), .D (new_AGEMA_signal_3608), .Q (new_AGEMA_signal_3609) ) ;
    buf_clk new_AGEMA_reg_buffer_2257 ( .C (clk), .D (new_AGEMA_signal_3616), .Q (new_AGEMA_signal_3617) ) ;
    buf_clk new_AGEMA_reg_buffer_2265 ( .C (clk), .D (new_AGEMA_signal_3624), .Q (new_AGEMA_signal_3625) ) ;
    buf_clk new_AGEMA_reg_buffer_2273 ( .C (clk), .D (new_AGEMA_signal_3632), .Q (new_AGEMA_signal_3633) ) ;
    buf_clk new_AGEMA_reg_buffer_2281 ( .C (clk), .D (new_AGEMA_signal_3640), .Q (new_AGEMA_signal_3641) ) ;
    buf_clk new_AGEMA_reg_buffer_2289 ( .C (clk), .D (new_AGEMA_signal_3648), .Q (new_AGEMA_signal_3649) ) ;
    buf_clk new_AGEMA_reg_buffer_2297 ( .C (clk), .D (new_AGEMA_signal_3656), .Q (new_AGEMA_signal_3657) ) ;
    buf_clk new_AGEMA_reg_buffer_2305 ( .C (clk), .D (new_AGEMA_signal_3664), .Q (new_AGEMA_signal_3665) ) ;
    buf_clk new_AGEMA_reg_buffer_2313 ( .C (clk), .D (new_AGEMA_signal_3672), .Q (new_AGEMA_signal_3673) ) ;
    buf_clk new_AGEMA_reg_buffer_2321 ( .C (clk), .D (new_AGEMA_signal_3680), .Q (new_AGEMA_signal_3681) ) ;
    buf_clk new_AGEMA_reg_buffer_2329 ( .C (clk), .D (new_AGEMA_signal_3688), .Q (new_AGEMA_signal_3689) ) ;
    buf_clk new_AGEMA_reg_buffer_2337 ( .C (clk), .D (new_AGEMA_signal_3696), .Q (new_AGEMA_signal_3697) ) ;
    buf_clk new_AGEMA_reg_buffer_2345 ( .C (clk), .D (new_AGEMA_signal_3704), .Q (new_AGEMA_signal_3705) ) ;
    buf_clk new_AGEMA_reg_buffer_2353 ( .C (clk), .D (new_AGEMA_signal_3712), .Q (new_AGEMA_signal_3713) ) ;
    buf_clk new_AGEMA_reg_buffer_2361 ( .C (clk), .D (new_AGEMA_signal_3720), .Q (new_AGEMA_signal_3721) ) ;
    buf_clk new_AGEMA_reg_buffer_2369 ( .C (clk), .D (new_AGEMA_signal_3728), .Q (new_AGEMA_signal_3729) ) ;
    buf_clk new_AGEMA_reg_buffer_2377 ( .C (clk), .D (new_AGEMA_signal_3736), .Q (new_AGEMA_signal_3737) ) ;
    buf_clk new_AGEMA_reg_buffer_2385 ( .C (clk), .D (new_AGEMA_signal_3744), .Q (new_AGEMA_signal_3745) ) ;
    buf_clk new_AGEMA_reg_buffer_2393 ( .C (clk), .D (new_AGEMA_signal_3752), .Q (new_AGEMA_signal_3753) ) ;
    buf_clk new_AGEMA_reg_buffer_2401 ( .C (clk), .D (new_AGEMA_signal_3760), .Q (new_AGEMA_signal_3761) ) ;
    buf_clk new_AGEMA_reg_buffer_2409 ( .C (clk), .D (new_AGEMA_signal_3768), .Q (new_AGEMA_signal_3769) ) ;
    buf_clk new_AGEMA_reg_buffer_2417 ( .C (clk), .D (new_AGEMA_signal_3776), .Q (new_AGEMA_signal_3777) ) ;
    buf_clk new_AGEMA_reg_buffer_2425 ( .C (clk), .D (new_AGEMA_signal_3784), .Q (new_AGEMA_signal_3785) ) ;
    buf_clk new_AGEMA_reg_buffer_2433 ( .C (clk), .D (new_AGEMA_signal_3792), .Q (new_AGEMA_signal_3793) ) ;
    buf_clk new_AGEMA_reg_buffer_2441 ( .C (clk), .D (new_AGEMA_signal_3800), .Q (new_AGEMA_signal_3801) ) ;
    buf_clk new_AGEMA_reg_buffer_2449 ( .C (clk), .D (new_AGEMA_signal_3808), .Q (new_AGEMA_signal_3809) ) ;
    buf_clk new_AGEMA_reg_buffer_2457 ( .C (clk), .D (new_AGEMA_signal_3816), .Q (new_AGEMA_signal_3817) ) ;
    buf_clk new_AGEMA_reg_buffer_2465 ( .C (clk), .D (new_AGEMA_signal_3824), .Q (new_AGEMA_signal_3825) ) ;
    buf_clk new_AGEMA_reg_buffer_2473 ( .C (clk), .D (new_AGEMA_signal_3832), .Q (new_AGEMA_signal_3833) ) ;
    buf_clk new_AGEMA_reg_buffer_2481 ( .C (clk), .D (new_AGEMA_signal_3840), .Q (new_AGEMA_signal_3841) ) ;
    buf_clk new_AGEMA_reg_buffer_2489 ( .C (clk), .D (new_AGEMA_signal_3848), .Q (new_AGEMA_signal_3849) ) ;
    buf_clk new_AGEMA_reg_buffer_2497 ( .C (clk), .D (new_AGEMA_signal_3856), .Q (new_AGEMA_signal_3857) ) ;
    buf_clk new_AGEMA_reg_buffer_2505 ( .C (clk), .D (new_AGEMA_signal_3864), .Q (new_AGEMA_signal_3865) ) ;
    buf_clk new_AGEMA_reg_buffer_2513 ( .C (clk), .D (new_AGEMA_signal_3872), .Q (new_AGEMA_signal_3873) ) ;
    buf_clk new_AGEMA_reg_buffer_2521 ( .C (clk), .D (new_AGEMA_signal_3880), .Q (new_AGEMA_signal_3881) ) ;
    buf_clk new_AGEMA_reg_buffer_2529 ( .C (clk), .D (new_AGEMA_signal_3888), .Q (new_AGEMA_signal_3889) ) ;
    buf_clk new_AGEMA_reg_buffer_2537 ( .C (clk), .D (new_AGEMA_signal_3896), .Q (new_AGEMA_signal_3897) ) ;
    buf_clk new_AGEMA_reg_buffer_2545 ( .C (clk), .D (new_AGEMA_signal_3904), .Q (new_AGEMA_signal_3905) ) ;
    buf_clk new_AGEMA_reg_buffer_2553 ( .C (clk), .D (new_AGEMA_signal_3912), .Q (new_AGEMA_signal_3913) ) ;
    buf_clk new_AGEMA_reg_buffer_2561 ( .C (clk), .D (new_AGEMA_signal_3920), .Q (new_AGEMA_signal_3921) ) ;
    buf_clk new_AGEMA_reg_buffer_2569 ( .C (clk), .D (new_AGEMA_signal_3928), .Q (new_AGEMA_signal_3929) ) ;
    buf_clk new_AGEMA_reg_buffer_2577 ( .C (clk), .D (new_AGEMA_signal_3936), .Q (new_AGEMA_signal_3937) ) ;
    buf_clk new_AGEMA_reg_buffer_2585 ( .C (clk), .D (new_AGEMA_signal_3944), .Q (new_AGEMA_signal_3945) ) ;
    buf_clk new_AGEMA_reg_buffer_2593 ( .C (clk), .D (new_AGEMA_signal_3952), .Q (new_AGEMA_signal_3953) ) ;
    buf_clk new_AGEMA_reg_buffer_2601 ( .C (clk), .D (new_AGEMA_signal_3960), .Q (new_AGEMA_signal_3961) ) ;
    buf_clk new_AGEMA_reg_buffer_2609 ( .C (clk), .D (new_AGEMA_signal_3968), .Q (new_AGEMA_signal_3969) ) ;
    buf_clk new_AGEMA_reg_buffer_2617 ( .C (clk), .D (new_AGEMA_signal_3976), .Q (new_AGEMA_signal_3977) ) ;
    buf_clk new_AGEMA_reg_buffer_2625 ( .C (clk), .D (new_AGEMA_signal_3984), .Q (new_AGEMA_signal_3985) ) ;
    buf_clk new_AGEMA_reg_buffer_2633 ( .C (clk), .D (new_AGEMA_signal_3992), .Q (new_AGEMA_signal_3993) ) ;
    buf_clk new_AGEMA_reg_buffer_2641 ( .C (clk), .D (new_AGEMA_signal_4000), .Q (new_AGEMA_signal_4001) ) ;
    buf_clk new_AGEMA_reg_buffer_2649 ( .C (clk), .D (new_AGEMA_signal_4008), .Q (new_AGEMA_signal_4009) ) ;
    buf_clk new_AGEMA_reg_buffer_2657 ( .C (clk), .D (new_AGEMA_signal_4016), .Q (new_AGEMA_signal_4017) ) ;
    buf_clk new_AGEMA_reg_buffer_2665 ( .C (clk), .D (new_AGEMA_signal_4024), .Q (new_AGEMA_signal_4025) ) ;
    buf_clk new_AGEMA_reg_buffer_2673 ( .C (clk), .D (new_AGEMA_signal_4032), .Q (new_AGEMA_signal_4033) ) ;
    buf_clk new_AGEMA_reg_buffer_2681 ( .C (clk), .D (new_AGEMA_signal_4040), .Q (new_AGEMA_signal_4041) ) ;
    buf_clk new_AGEMA_reg_buffer_2689 ( .C (clk), .D (new_AGEMA_signal_4048), .Q (new_AGEMA_signal_4049) ) ;
    buf_clk new_AGEMA_reg_buffer_2697 ( .C (clk), .D (new_AGEMA_signal_4056), .Q (new_AGEMA_signal_4057) ) ;
    buf_clk new_AGEMA_reg_buffer_2705 ( .C (clk), .D (new_AGEMA_signal_4064), .Q (new_AGEMA_signal_4065) ) ;
    buf_clk new_AGEMA_reg_buffer_2713 ( .C (clk), .D (new_AGEMA_signal_4072), .Q (new_AGEMA_signal_4073) ) ;
    buf_clk new_AGEMA_reg_buffer_2721 ( .C (clk), .D (new_AGEMA_signal_4080), .Q (new_AGEMA_signal_4081) ) ;
    buf_clk new_AGEMA_reg_buffer_2729 ( .C (clk), .D (new_AGEMA_signal_4088), .Q (new_AGEMA_signal_4089) ) ;
    buf_clk new_AGEMA_reg_buffer_2737 ( .C (clk), .D (new_AGEMA_signal_4096), .Q (new_AGEMA_signal_4097) ) ;
    buf_clk new_AGEMA_reg_buffer_2745 ( .C (clk), .D (new_AGEMA_signal_4104), .Q (new_AGEMA_signal_4105) ) ;
    buf_clk new_AGEMA_reg_buffer_2753 ( .C (clk), .D (new_AGEMA_signal_4112), .Q (new_AGEMA_signal_4113) ) ;
    buf_clk new_AGEMA_reg_buffer_2761 ( .C (clk), .D (new_AGEMA_signal_4120), .Q (new_AGEMA_signal_4121) ) ;
    buf_clk new_AGEMA_reg_buffer_2769 ( .C (clk), .D (new_AGEMA_signal_4128), .Q (new_AGEMA_signal_4129) ) ;
    buf_clk new_AGEMA_reg_buffer_2777 ( .C (clk), .D (new_AGEMA_signal_4136), .Q (new_AGEMA_signal_4137) ) ;
    buf_clk new_AGEMA_reg_buffer_2785 ( .C (clk), .D (new_AGEMA_signal_4144), .Q (new_AGEMA_signal_4145) ) ;
    buf_clk new_AGEMA_reg_buffer_2793 ( .C (clk), .D (new_AGEMA_signal_4152), .Q (new_AGEMA_signal_4153) ) ;
    buf_clk new_AGEMA_reg_buffer_2801 ( .C (clk), .D (new_AGEMA_signal_4160), .Q (new_AGEMA_signal_4161) ) ;
    buf_clk new_AGEMA_reg_buffer_2809 ( .C (clk), .D (new_AGEMA_signal_4168), .Q (new_AGEMA_signal_4169) ) ;
    buf_clk new_AGEMA_reg_buffer_2817 ( .C (clk), .D (new_AGEMA_signal_4176), .Q (new_AGEMA_signal_4177) ) ;
    buf_clk new_AGEMA_reg_buffer_2825 ( .C (clk), .D (new_AGEMA_signal_4184), .Q (new_AGEMA_signal_4185) ) ;
    buf_clk new_AGEMA_reg_buffer_2833 ( .C (clk), .D (new_AGEMA_signal_4192), .Q (new_AGEMA_signal_4193) ) ;
    buf_clk new_AGEMA_reg_buffer_2841 ( .C (clk), .D (new_AGEMA_signal_4200), .Q (new_AGEMA_signal_4201) ) ;
    buf_clk new_AGEMA_reg_buffer_2849 ( .C (clk), .D (new_AGEMA_signal_4208), .Q (new_AGEMA_signal_4209) ) ;
    buf_clk new_AGEMA_reg_buffer_2857 ( .C (clk), .D (new_AGEMA_signal_4216), .Q (new_AGEMA_signal_4217) ) ;
    buf_clk new_AGEMA_reg_buffer_2865 ( .C (clk), .D (new_AGEMA_signal_4224), .Q (new_AGEMA_signal_4225) ) ;
    buf_clk new_AGEMA_reg_buffer_2873 ( .C (clk), .D (new_AGEMA_signal_4232), .Q (new_AGEMA_signal_4233) ) ;
    buf_clk new_AGEMA_reg_buffer_2881 ( .C (clk), .D (new_AGEMA_signal_4240), .Q (new_AGEMA_signal_4241) ) ;
    buf_clk new_AGEMA_reg_buffer_2889 ( .C (clk), .D (new_AGEMA_signal_4248), .Q (new_AGEMA_signal_4249) ) ;
    buf_clk new_AGEMA_reg_buffer_2897 ( .C (clk), .D (new_AGEMA_signal_4256), .Q (new_AGEMA_signal_4257) ) ;
    buf_clk new_AGEMA_reg_buffer_2905 ( .C (clk), .D (new_AGEMA_signal_4264), .Q (new_AGEMA_signal_4265) ) ;
    buf_clk new_AGEMA_reg_buffer_2913 ( .C (clk), .D (new_AGEMA_signal_4272), .Q (new_AGEMA_signal_4273) ) ;
    buf_clk new_AGEMA_reg_buffer_2921 ( .C (clk), .D (new_AGEMA_signal_4280), .Q (new_AGEMA_signal_4281) ) ;
    buf_clk new_AGEMA_reg_buffer_2929 ( .C (clk), .D (new_AGEMA_signal_4288), .Q (new_AGEMA_signal_4289) ) ;
    buf_clk new_AGEMA_reg_buffer_2937 ( .C (clk), .D (new_AGEMA_signal_4296), .Q (new_AGEMA_signal_4297) ) ;
    buf_clk new_AGEMA_reg_buffer_2945 ( .C (clk), .D (new_AGEMA_signal_4304), .Q (new_AGEMA_signal_4305) ) ;
    buf_clk new_AGEMA_reg_buffer_2953 ( .C (clk), .D (new_AGEMA_signal_4312), .Q (new_AGEMA_signal_4313) ) ;
    buf_clk new_AGEMA_reg_buffer_2961 ( .C (clk), .D (new_AGEMA_signal_4320), .Q (new_AGEMA_signal_4321) ) ;
    buf_clk new_AGEMA_reg_buffer_2969 ( .C (clk), .D (new_AGEMA_signal_4328), .Q (new_AGEMA_signal_4329) ) ;
    buf_clk new_AGEMA_reg_buffer_2977 ( .C (clk), .D (new_AGEMA_signal_4336), .Q (new_AGEMA_signal_4337) ) ;
    buf_clk new_AGEMA_reg_buffer_2985 ( .C (clk), .D (new_AGEMA_signal_4344), .Q (new_AGEMA_signal_4345) ) ;
    buf_clk new_AGEMA_reg_buffer_2993 ( .C (clk), .D (new_AGEMA_signal_4352), .Q (new_AGEMA_signal_4353) ) ;
    buf_clk new_AGEMA_reg_buffer_3001 ( .C (clk), .D (new_AGEMA_signal_4360), .Q (new_AGEMA_signal_4361) ) ;
    buf_clk new_AGEMA_reg_buffer_3009 ( .C (clk), .D (new_AGEMA_signal_4368), .Q (new_AGEMA_signal_4369) ) ;
    buf_clk new_AGEMA_reg_buffer_3017 ( .C (clk), .D (new_AGEMA_signal_4376), .Q (new_AGEMA_signal_4377) ) ;
    buf_clk new_AGEMA_reg_buffer_3025 ( .C (clk), .D (new_AGEMA_signal_4384), .Q (new_AGEMA_signal_4385) ) ;
    buf_clk new_AGEMA_reg_buffer_3033 ( .C (clk), .D (new_AGEMA_signal_4392), .Q (new_AGEMA_signal_4393) ) ;
    buf_clk new_AGEMA_reg_buffer_3041 ( .C (clk), .D (new_AGEMA_signal_4400), .Q (new_AGEMA_signal_4401) ) ;
    buf_clk new_AGEMA_reg_buffer_3049 ( .C (clk), .D (new_AGEMA_signal_4408), .Q (new_AGEMA_signal_4409) ) ;
    buf_clk new_AGEMA_reg_buffer_3057 ( .C (clk), .D (new_AGEMA_signal_4416), .Q (new_AGEMA_signal_4417) ) ;
    buf_clk new_AGEMA_reg_buffer_3065 ( .C (clk), .D (new_AGEMA_signal_4424), .Q (new_AGEMA_signal_4425) ) ;
    buf_clk new_AGEMA_reg_buffer_3259 ( .C (clk), .D (AddRoundKeyOutput[63]), .Q (new_AGEMA_signal_4619) ) ;
    buf_clk new_AGEMA_reg_buffer_3261 ( .C (clk), .D (new_AGEMA_signal_1906), .Q (new_AGEMA_signal_4621) ) ;
    buf_clk new_AGEMA_reg_buffer_3263 ( .C (clk), .D (AddRoundKeyOutput[61]), .Q (new_AGEMA_signal_4623) ) ;
    buf_clk new_AGEMA_reg_buffer_3265 ( .C (clk), .D (new_AGEMA_signal_1904), .Q (new_AGEMA_signal_4625) ) ;
    buf_clk new_AGEMA_reg_buffer_3267 ( .C (clk), .D (AddRoundKeyOutput[59]), .Q (new_AGEMA_signal_4627) ) ;
    buf_clk new_AGEMA_reg_buffer_3269 ( .C (clk), .D (new_AGEMA_signal_1902), .Q (new_AGEMA_signal_4629) ) ;
    buf_clk new_AGEMA_reg_buffer_3271 ( .C (clk), .D (AddRoundKeyOutput[57]), .Q (new_AGEMA_signal_4631) ) ;
    buf_clk new_AGEMA_reg_buffer_3273 ( .C (clk), .D (new_AGEMA_signal_1900), .Q (new_AGEMA_signal_4633) ) ;
    buf_clk new_AGEMA_reg_buffer_3275 ( .C (clk), .D (AddRoundKeyOutput[55]), .Q (new_AGEMA_signal_4635) ) ;
    buf_clk new_AGEMA_reg_buffer_3277 ( .C (clk), .D (new_AGEMA_signal_1898), .Q (new_AGEMA_signal_4637) ) ;
    buf_clk new_AGEMA_reg_buffer_3279 ( .C (clk), .D (AddRoundKeyOutput[53]), .Q (new_AGEMA_signal_4639) ) ;
    buf_clk new_AGEMA_reg_buffer_3281 ( .C (clk), .D (new_AGEMA_signal_1896), .Q (new_AGEMA_signal_4641) ) ;
    buf_clk new_AGEMA_reg_buffer_3283 ( .C (clk), .D (AddRoundKeyOutput[51]), .Q (new_AGEMA_signal_4643) ) ;
    buf_clk new_AGEMA_reg_buffer_3285 ( .C (clk), .D (new_AGEMA_signal_1894), .Q (new_AGEMA_signal_4645) ) ;
    buf_clk new_AGEMA_reg_buffer_3287 ( .C (clk), .D (AddRoundKeyOutput[49]), .Q (new_AGEMA_signal_4647) ) ;
    buf_clk new_AGEMA_reg_buffer_3289 ( .C (clk), .D (new_AGEMA_signal_1892), .Q (new_AGEMA_signal_4649) ) ;
    buf_clk new_AGEMA_reg_buffer_3291 ( .C (clk), .D (AddRoundKeyOutput[47]), .Q (new_AGEMA_signal_4651) ) ;
    buf_clk new_AGEMA_reg_buffer_3293 ( .C (clk), .D (new_AGEMA_signal_1914), .Q (new_AGEMA_signal_4653) ) ;
    buf_clk new_AGEMA_reg_buffer_3295 ( .C (clk), .D (AddRoundKeyOutput[45]), .Q (new_AGEMA_signal_4655) ) ;
    buf_clk new_AGEMA_reg_buffer_3297 ( .C (clk), .D (new_AGEMA_signal_1912), .Q (new_AGEMA_signal_4657) ) ;
    buf_clk new_AGEMA_reg_buffer_3299 ( .C (clk), .D (AddRoundKeyOutput[43]), .Q (new_AGEMA_signal_4659) ) ;
    buf_clk new_AGEMA_reg_buffer_3301 ( .C (clk), .D (new_AGEMA_signal_1910), .Q (new_AGEMA_signal_4661) ) ;
    buf_clk new_AGEMA_reg_buffer_3303 ( .C (clk), .D (AddRoundKeyOutput[41]), .Q (new_AGEMA_signal_4663) ) ;
    buf_clk new_AGEMA_reg_buffer_3305 ( .C (clk), .D (new_AGEMA_signal_1908), .Q (new_AGEMA_signal_4665) ) ;
    buf_clk new_AGEMA_reg_buffer_3307 ( .C (clk), .D (AddRoundKeyOutput[39]), .Q (new_AGEMA_signal_4667) ) ;
    buf_clk new_AGEMA_reg_buffer_3309 ( .C (clk), .D (new_AGEMA_signal_1922), .Q (new_AGEMA_signal_4669) ) ;
    buf_clk new_AGEMA_reg_buffer_3311 ( .C (clk), .D (AddRoundKeyOutput[37]), .Q (new_AGEMA_signal_4671) ) ;
    buf_clk new_AGEMA_reg_buffer_3313 ( .C (clk), .D (new_AGEMA_signal_1920), .Q (new_AGEMA_signal_4673) ) ;
    buf_clk new_AGEMA_reg_buffer_3315 ( .C (clk), .D (AddRoundKeyOutput[35]), .Q (new_AGEMA_signal_4675) ) ;
    buf_clk new_AGEMA_reg_buffer_3317 ( .C (clk), .D (new_AGEMA_signal_1918), .Q (new_AGEMA_signal_4677) ) ;
    buf_clk new_AGEMA_reg_buffer_3319 ( .C (clk), .D (AddRoundKeyOutput[33]), .Q (new_AGEMA_signal_4679) ) ;
    buf_clk new_AGEMA_reg_buffer_3321 ( .C (clk), .D (new_AGEMA_signal_1916), .Q (new_AGEMA_signal_4681) ) ;
    buf_clk new_AGEMA_reg_buffer_3323 ( .C (clk), .D (AddRoundKeyOutput[31]), .Q (new_AGEMA_signal_4683) ) ;
    buf_clk new_AGEMA_reg_buffer_3325 ( .C (clk), .D (new_AGEMA_signal_1858), .Q (new_AGEMA_signal_4685) ) ;
    buf_clk new_AGEMA_reg_buffer_3327 ( .C (clk), .D (AddRoundKeyOutput[29]), .Q (new_AGEMA_signal_4687) ) ;
    buf_clk new_AGEMA_reg_buffer_3329 ( .C (clk), .D (new_AGEMA_signal_1856), .Q (new_AGEMA_signal_4689) ) ;
    buf_clk new_AGEMA_reg_buffer_3331 ( .C (clk), .D (AddRoundKeyOutput[27]), .Q (new_AGEMA_signal_4691) ) ;
    buf_clk new_AGEMA_reg_buffer_3333 ( .C (clk), .D (new_AGEMA_signal_1854), .Q (new_AGEMA_signal_4693) ) ;
    buf_clk new_AGEMA_reg_buffer_3335 ( .C (clk), .D (AddRoundKeyOutput[25]), .Q (new_AGEMA_signal_4695) ) ;
    buf_clk new_AGEMA_reg_buffer_3337 ( .C (clk), .D (new_AGEMA_signal_1852), .Q (new_AGEMA_signal_4697) ) ;
    buf_clk new_AGEMA_reg_buffer_3339 ( .C (clk), .D (AddRoundKeyOutput[23]), .Q (new_AGEMA_signal_4699) ) ;
    buf_clk new_AGEMA_reg_buffer_3341 ( .C (clk), .D (new_AGEMA_signal_1850), .Q (new_AGEMA_signal_4701) ) ;
    buf_clk new_AGEMA_reg_buffer_3343 ( .C (clk), .D (AddRoundKeyOutput[21]), .Q (new_AGEMA_signal_4703) ) ;
    buf_clk new_AGEMA_reg_buffer_3345 ( .C (clk), .D (new_AGEMA_signal_1848), .Q (new_AGEMA_signal_4705) ) ;
    buf_clk new_AGEMA_reg_buffer_3347 ( .C (clk), .D (AddRoundKeyOutput[19]), .Q (new_AGEMA_signal_4707) ) ;
    buf_clk new_AGEMA_reg_buffer_3349 ( .C (clk), .D (new_AGEMA_signal_1846), .Q (new_AGEMA_signal_4709) ) ;
    buf_clk new_AGEMA_reg_buffer_3351 ( .C (clk), .D (AddRoundKeyOutput[17]), .Q (new_AGEMA_signal_4711) ) ;
    buf_clk new_AGEMA_reg_buffer_3353 ( .C (clk), .D (new_AGEMA_signal_1844), .Q (new_AGEMA_signal_4713) ) ;
    buf_clk new_AGEMA_reg_buffer_3355 ( .C (clk), .D (AddRoundKeyOutput[15]), .Q (new_AGEMA_signal_4715) ) ;
    buf_clk new_AGEMA_reg_buffer_3357 ( .C (clk), .D (new_AGEMA_signal_1842), .Q (new_AGEMA_signal_4717) ) ;
    buf_clk new_AGEMA_reg_buffer_3359 ( .C (clk), .D (AddRoundKeyOutput[13]), .Q (new_AGEMA_signal_4719) ) ;
    buf_clk new_AGEMA_reg_buffer_3361 ( .C (clk), .D (new_AGEMA_signal_1840), .Q (new_AGEMA_signal_4721) ) ;
    buf_clk new_AGEMA_reg_buffer_3363 ( .C (clk), .D (AddRoundKeyOutput[11]), .Q (new_AGEMA_signal_4723) ) ;
    buf_clk new_AGEMA_reg_buffer_3365 ( .C (clk), .D (new_AGEMA_signal_1838), .Q (new_AGEMA_signal_4725) ) ;
    buf_clk new_AGEMA_reg_buffer_3367 ( .C (clk), .D (AddRoundKeyOutput[9]), .Q (new_AGEMA_signal_4727) ) ;
    buf_clk new_AGEMA_reg_buffer_3369 ( .C (clk), .D (new_AGEMA_signal_1836), .Q (new_AGEMA_signal_4729) ) ;
    buf_clk new_AGEMA_reg_buffer_3371 ( .C (clk), .D (AddRoundKeyOutput[7]), .Q (new_AGEMA_signal_4731) ) ;
    buf_clk new_AGEMA_reg_buffer_3373 ( .C (clk), .D (new_AGEMA_signal_1834), .Q (new_AGEMA_signal_4733) ) ;
    buf_clk new_AGEMA_reg_buffer_3375 ( .C (clk), .D (AddRoundKeyOutput[5]), .Q (new_AGEMA_signal_4735) ) ;
    buf_clk new_AGEMA_reg_buffer_3377 ( .C (clk), .D (new_AGEMA_signal_1832), .Q (new_AGEMA_signal_4737) ) ;
    buf_clk new_AGEMA_reg_buffer_3379 ( .C (clk), .D (AddRoundKeyOutput[3]), .Q (new_AGEMA_signal_4739) ) ;
    buf_clk new_AGEMA_reg_buffer_3381 ( .C (clk), .D (new_AGEMA_signal_1830), .Q (new_AGEMA_signal_4741) ) ;
    buf_clk new_AGEMA_reg_buffer_3383 ( .C (clk), .D (AddRoundKeyOutput[1]), .Q (new_AGEMA_signal_4743) ) ;
    buf_clk new_AGEMA_reg_buffer_3385 ( .C (clk), .D (new_AGEMA_signal_1828), .Q (new_AGEMA_signal_4745) ) ;
    buf_clk new_AGEMA_reg_buffer_3393 ( .C (clk), .D (new_AGEMA_signal_4752), .Q (new_AGEMA_signal_4753) ) ;
    buf_clk new_AGEMA_reg_buffer_3401 ( .C (clk), .D (new_AGEMA_signal_4760), .Q (new_AGEMA_signal_4761) ) ;
    buf_clk new_AGEMA_reg_buffer_3409 ( .C (clk), .D (new_AGEMA_signal_4768), .Q (new_AGEMA_signal_4769) ) ;
    buf_clk new_AGEMA_reg_buffer_3417 ( .C (clk), .D (new_AGEMA_signal_4776), .Q (new_AGEMA_signal_4777) ) ;
    buf_clk new_AGEMA_reg_buffer_3425 ( .C (clk), .D (new_AGEMA_signal_4784), .Q (new_AGEMA_signal_4785) ) ;
    buf_clk new_AGEMA_reg_buffer_3433 ( .C (clk), .D (new_AGEMA_signal_4792), .Q (new_AGEMA_signal_4793) ) ;
    buf_clk new_AGEMA_reg_buffer_3441 ( .C (clk), .D (new_AGEMA_signal_4800), .Q (new_AGEMA_signal_4801) ) ;
    buf_clk new_AGEMA_reg_buffer_3449 ( .C (clk), .D (new_AGEMA_signal_4808), .Q (new_AGEMA_signal_4809) ) ;
    buf_clk new_AGEMA_reg_buffer_3457 ( .C (clk), .D (new_AGEMA_signal_4816), .Q (new_AGEMA_signal_4817) ) ;
    buf_clk new_AGEMA_reg_buffer_3465 ( .C (clk), .D (new_AGEMA_signal_4824), .Q (new_AGEMA_signal_4825) ) ;

    /* cells in depth 8 */
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_0_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1374, Feedback[0]}), .a ({new_AGEMA_signal_3418, new_AGEMA_signal_3410}), .c ({new_AGEMA_signal_1580, MCOutput[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_2_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1372, Feedback[2]}), .a ({new_AGEMA_signal_3434, new_AGEMA_signal_3426}), .c ({new_AGEMA_signal_1584, MCOutput[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_4_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1378, Feedback[4]}), .a ({new_AGEMA_signal_3450, new_AGEMA_signal_3442}), .c ({new_AGEMA_signal_1588, MCOutput[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_6_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1376, Feedback[6]}), .a ({new_AGEMA_signal_3466, new_AGEMA_signal_3458}), .c ({new_AGEMA_signal_1592, MCOutput[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_8_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1382, Feedback[8]}), .a ({new_AGEMA_signal_3482, new_AGEMA_signal_3474}), .c ({new_AGEMA_signal_1596, MCOutput[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_10_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1380, Feedback[10]}), .a ({new_AGEMA_signal_3498, new_AGEMA_signal_3490}), .c ({new_AGEMA_signal_1600, MCOutput[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_12_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1386, Feedback[12]}), .a ({new_AGEMA_signal_3514, new_AGEMA_signal_3506}), .c ({new_AGEMA_signal_1604, MCOutput[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_14_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1384, Feedback[14]}), .a ({new_AGEMA_signal_3530, new_AGEMA_signal_3522}), .c ({new_AGEMA_signal_1608, MCOutput[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_16_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1390, Feedback[16]}), .a ({new_AGEMA_signal_3546, new_AGEMA_signal_3538}), .c ({new_AGEMA_signal_1612, MCOutput[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_18_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1388, Feedback[18]}), .a ({new_AGEMA_signal_3562, new_AGEMA_signal_3554}), .c ({new_AGEMA_signal_1616, MCOutput[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_20_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1394, Feedback[20]}), .a ({new_AGEMA_signal_3578, new_AGEMA_signal_3570}), .c ({new_AGEMA_signal_1620, MCOutput[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_22_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1392, Feedback[22]}), .a ({new_AGEMA_signal_3594, new_AGEMA_signal_3586}), .c ({new_AGEMA_signal_1624, MCOutput[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_24_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1398, Feedback[24]}), .a ({new_AGEMA_signal_3610, new_AGEMA_signal_3602}), .c ({new_AGEMA_signal_1628, MCOutput[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_26_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1396, Feedback[26]}), .a ({new_AGEMA_signal_3626, new_AGEMA_signal_3618}), .c ({new_AGEMA_signal_1632, MCOutput[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_28_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1402, Feedback[28]}), .a ({new_AGEMA_signal_3642, new_AGEMA_signal_3634}), .c ({new_AGEMA_signal_1636, MCOutput[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_30_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1400, Feedback[30]}), .a ({new_AGEMA_signal_3658, new_AGEMA_signal_3650}), .c ({new_AGEMA_signal_1640, MCOutput[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_32_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1406, Feedback[32]}), .a ({new_AGEMA_signal_3674, new_AGEMA_signal_3666}), .c ({new_AGEMA_signal_1644, MCInput[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_34_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1404, Feedback[34]}), .a ({new_AGEMA_signal_3690, new_AGEMA_signal_3682}), .c ({new_AGEMA_signal_1648, MCInput[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_36_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1410, Feedback[36]}), .a ({new_AGEMA_signal_3706, new_AGEMA_signal_3698}), .c ({new_AGEMA_signal_1652, MCInput[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_38_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1408, Feedback[38]}), .a ({new_AGEMA_signal_3722, new_AGEMA_signal_3714}), .c ({new_AGEMA_signal_1656, MCInput[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_40_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1414, Feedback[40]}), .a ({new_AGEMA_signal_3738, new_AGEMA_signal_3730}), .c ({new_AGEMA_signal_1660, MCInput[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_42_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1412, Feedback[42]}), .a ({new_AGEMA_signal_3754, new_AGEMA_signal_3746}), .c ({new_AGEMA_signal_1664, MCInput[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_44_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1418, Feedback[44]}), .a ({new_AGEMA_signal_3770, new_AGEMA_signal_3762}), .c ({new_AGEMA_signal_1668, MCInput[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_46_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1416, Feedback[46]}), .a ({new_AGEMA_signal_3786, new_AGEMA_signal_3778}), .c ({new_AGEMA_signal_1672, MCInput[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_48_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1422, Feedback[48]}), .a ({new_AGEMA_signal_3802, new_AGEMA_signal_3794}), .c ({new_AGEMA_signal_1676, MCInput[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_50_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1420, Feedback[50]}), .a ({new_AGEMA_signal_3818, new_AGEMA_signal_3810}), .c ({new_AGEMA_signal_1680, MCInput[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_52_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1426, Feedback[52]}), .a ({new_AGEMA_signal_3834, new_AGEMA_signal_3826}), .c ({new_AGEMA_signal_1684, MCInput[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_54_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1424, Feedback[54]}), .a ({new_AGEMA_signal_3850, new_AGEMA_signal_3842}), .c ({new_AGEMA_signal_1688, MCInput[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_56_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1430, Feedback[56]}), .a ({new_AGEMA_signal_3866, new_AGEMA_signal_3858}), .c ({new_AGEMA_signal_1692, MCInput[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_58_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1428, Feedback[58]}), .a ({new_AGEMA_signal_3882, new_AGEMA_signal_3874}), .c ({new_AGEMA_signal_1696, MCInput[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_60_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1434, Feedback[60]}), .a ({new_AGEMA_signal_3898, new_AGEMA_signal_3890}), .c ({new_AGEMA_signal_1700, MCInput[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) InputMUX_MUXInst_62_U1 ( .s (new_AGEMA_signal_3402), .b ({new_AGEMA_signal_1432, Feedback[62]}), .a ({new_AGEMA_signal_3914, new_AGEMA_signal_3906}), .c ({new_AGEMA_signal_1704, MCInput[62]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_0_U3 ( .a ({new_AGEMA_signal_1716, MCInst_XOR_r0_Inst_0_n2}), .b ({new_AGEMA_signal_1715, MCInst_XOR_r0_Inst_0_n1}), .c ({new_AGEMA_signal_1795, MCOutput[48]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_0_U2 ( .a ({new_AGEMA_signal_1612, MCOutput[16]}), .b ({new_AGEMA_signal_1580, MCOutput[0]}), .c ({new_AGEMA_signal_1715, MCInst_XOR_r0_Inst_0_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1676, MCInput[48]}), .c ({new_AGEMA_signal_1716, MCInst_XOR_r0_Inst_0_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_0_U2 ( .a ({new_AGEMA_signal_1717, MCInst_XOR_r1_Inst_0_n1}), .b ({new_AGEMA_signal_1580, MCOutput[0]}), .c ({new_AGEMA_signal_1796, MCOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1644, MCInput[32]}), .c ({new_AGEMA_signal_1717, MCInst_XOR_r1_Inst_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_2_U3 ( .a ({new_AGEMA_signal_1722, MCInst_XOR_r0_Inst_2_n2}), .b ({new_AGEMA_signal_1721, MCInst_XOR_r0_Inst_2_n1}), .c ({new_AGEMA_signal_1799, MCOutput[50]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_2_U2 ( .a ({new_AGEMA_signal_1616, MCOutput[18]}), .b ({new_AGEMA_signal_1584, MCOutput[2]}), .c ({new_AGEMA_signal_1721, MCInst_XOR_r0_Inst_2_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1680, MCInput[50]}), .c ({new_AGEMA_signal_1722, MCInst_XOR_r0_Inst_2_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_2_U2 ( .a ({new_AGEMA_signal_1723, MCInst_XOR_r1_Inst_2_n1}), .b ({new_AGEMA_signal_1584, MCOutput[2]}), .c ({new_AGEMA_signal_1800, MCOutput[34]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1648, MCInput[34]}), .c ({new_AGEMA_signal_1723, MCInst_XOR_r1_Inst_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_4_U3 ( .a ({new_AGEMA_signal_1728, MCInst_XOR_r0_Inst_4_n2}), .b ({new_AGEMA_signal_1727, MCInst_XOR_r0_Inst_4_n1}), .c ({new_AGEMA_signal_1803, MCOutput[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_4_U2 ( .a ({new_AGEMA_signal_1620, MCOutput[20]}), .b ({new_AGEMA_signal_1588, MCOutput[4]}), .c ({new_AGEMA_signal_1727, MCInst_XOR_r0_Inst_4_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_4_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1684, MCInput[52]}), .c ({new_AGEMA_signal_1728, MCInst_XOR_r0_Inst_4_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_4_U2 ( .a ({new_AGEMA_signal_1729, MCInst_XOR_r1_Inst_4_n1}), .b ({new_AGEMA_signal_1588, MCOutput[4]}), .c ({new_AGEMA_signal_1804, MCOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_4_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1652, MCInput[36]}), .c ({new_AGEMA_signal_1729, MCInst_XOR_r1_Inst_4_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_6_U3 ( .a ({new_AGEMA_signal_1734, MCInst_XOR_r0_Inst_6_n2}), .b ({new_AGEMA_signal_1733, MCInst_XOR_r0_Inst_6_n1}), .c ({new_AGEMA_signal_1807, MCOutput[54]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_6_U2 ( .a ({new_AGEMA_signal_1624, MCOutput[22]}), .b ({new_AGEMA_signal_1592, MCOutput[6]}), .c ({new_AGEMA_signal_1733, MCInst_XOR_r0_Inst_6_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_6_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1688, MCInput[54]}), .c ({new_AGEMA_signal_1734, MCInst_XOR_r0_Inst_6_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_6_U2 ( .a ({new_AGEMA_signal_1735, MCInst_XOR_r1_Inst_6_n1}), .b ({new_AGEMA_signal_1592, MCOutput[6]}), .c ({new_AGEMA_signal_1808, MCOutput[38]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_6_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1656, MCInput[38]}), .c ({new_AGEMA_signal_1735, MCInst_XOR_r1_Inst_6_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_8_U3 ( .a ({new_AGEMA_signal_1740, MCInst_XOR_r0_Inst_8_n2}), .b ({new_AGEMA_signal_1739, MCInst_XOR_r0_Inst_8_n1}), .c ({new_AGEMA_signal_1811, MCOutput[56]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_8_U2 ( .a ({new_AGEMA_signal_1628, MCOutput[24]}), .b ({new_AGEMA_signal_1596, MCOutput[8]}), .c ({new_AGEMA_signal_1739, MCInst_XOR_r0_Inst_8_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_8_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1692, MCInput[56]}), .c ({new_AGEMA_signal_1740, MCInst_XOR_r0_Inst_8_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_8_U2 ( .a ({new_AGEMA_signal_1741, MCInst_XOR_r1_Inst_8_n1}), .b ({new_AGEMA_signal_1596, MCOutput[8]}), .c ({new_AGEMA_signal_1812, MCOutput[40]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_8_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1660, MCInput[40]}), .c ({new_AGEMA_signal_1741, MCInst_XOR_r1_Inst_8_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_10_U3 ( .a ({new_AGEMA_signal_1746, MCInst_XOR_r0_Inst_10_n2}), .b ({new_AGEMA_signal_1745, MCInst_XOR_r0_Inst_10_n1}), .c ({new_AGEMA_signal_1815, MCOutput[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_10_U2 ( .a ({new_AGEMA_signal_1632, MCOutput[26]}), .b ({new_AGEMA_signal_1600, MCOutput[10]}), .c ({new_AGEMA_signal_1745, MCInst_XOR_r0_Inst_10_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_10_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1696, MCInput[58]}), .c ({new_AGEMA_signal_1746, MCInst_XOR_r0_Inst_10_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_10_U2 ( .a ({new_AGEMA_signal_1747, MCInst_XOR_r1_Inst_10_n1}), .b ({new_AGEMA_signal_1600, MCOutput[10]}), .c ({new_AGEMA_signal_1816, MCOutput[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_10_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1664, MCInput[42]}), .c ({new_AGEMA_signal_1747, MCInst_XOR_r1_Inst_10_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_12_U3 ( .a ({new_AGEMA_signal_1752, MCInst_XOR_r0_Inst_12_n2}), .b ({new_AGEMA_signal_1751, MCInst_XOR_r0_Inst_12_n1}), .c ({new_AGEMA_signal_1819, MCOutput[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_12_U2 ( .a ({new_AGEMA_signal_1636, MCOutput[28]}), .b ({new_AGEMA_signal_1604, MCOutput[12]}), .c ({new_AGEMA_signal_1751, MCInst_XOR_r0_Inst_12_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_12_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1700, MCInput[60]}), .c ({new_AGEMA_signal_1752, MCInst_XOR_r0_Inst_12_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_12_U2 ( .a ({new_AGEMA_signal_1753, MCInst_XOR_r1_Inst_12_n1}), .b ({new_AGEMA_signal_1604, MCOutput[12]}), .c ({new_AGEMA_signal_1820, MCOutput[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_12_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1668, MCInput[44]}), .c ({new_AGEMA_signal_1753, MCInst_XOR_r1_Inst_12_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_14_U3 ( .a ({new_AGEMA_signal_1758, MCInst_XOR_r0_Inst_14_n2}), .b ({new_AGEMA_signal_1757, MCInst_XOR_r0_Inst_14_n1}), .c ({new_AGEMA_signal_1823, MCOutput[62]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_14_U2 ( .a ({new_AGEMA_signal_1640, MCOutput[30]}), .b ({new_AGEMA_signal_1608, MCOutput[14]}), .c ({new_AGEMA_signal_1757, MCInst_XOR_r0_Inst_14_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r0_Inst_14_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1704, MCInput[62]}), .c ({new_AGEMA_signal_1758, MCInst_XOR_r0_Inst_14_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_14_U2 ( .a ({new_AGEMA_signal_1759, MCInst_XOR_r1_Inst_14_n1}), .b ({new_AGEMA_signal_1608, MCOutput[14]}), .c ({new_AGEMA_signal_1824, MCOutput[46]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) MCInst_XOR_r1_Inst_14_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1672, MCInput[46]}), .c ({new_AGEMA_signal_1759, MCInst_XOR_r1_Inst_14_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_1859, AddKeyXOR1_XORInst_0_0_n1}), .b ({new_AGEMA_signal_3930, new_AGEMA_signal_3922}), .c ({new_AGEMA_signal_1891, AddRoundKeyOutput[48]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_0_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1795, MCOutput[48]}), .c ({new_AGEMA_signal_1859, AddKeyXOR1_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_1861, AddKeyXOR1_XORInst_0_2_n1}), .b ({new_AGEMA_signal_3946, new_AGEMA_signal_3938}), .c ({new_AGEMA_signal_1893, AddRoundKeyOutput[50]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_0_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1799, MCOutput[50]}), .c ({new_AGEMA_signal_1861, AddKeyXOR1_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_1863, AddKeyXOR1_XORInst_1_0_n1}), .b ({new_AGEMA_signal_3962, new_AGEMA_signal_3954}), .c ({new_AGEMA_signal_1895, AddRoundKeyOutput[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_1_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1803, MCOutput[52]}), .c ({new_AGEMA_signal_1863, AddKeyXOR1_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_1865, AddKeyXOR1_XORInst_1_2_n1}), .b ({new_AGEMA_signal_3978, new_AGEMA_signal_3970}), .c ({new_AGEMA_signal_1897, AddRoundKeyOutput[54]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_1_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1807, MCOutput[54]}), .c ({new_AGEMA_signal_1865, AddKeyXOR1_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_1867, AddKeyXOR1_XORInst_2_0_n1}), .b ({new_AGEMA_signal_3994, new_AGEMA_signal_3986}), .c ({new_AGEMA_signal_1899, AddRoundKeyOutput[56]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_2_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1811, MCOutput[56]}), .c ({new_AGEMA_signal_1867, AddKeyXOR1_XORInst_2_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_1869, AddKeyXOR1_XORInst_2_2_n1}), .b ({new_AGEMA_signal_4010, new_AGEMA_signal_4002}), .c ({new_AGEMA_signal_1901, AddRoundKeyOutput[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_2_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1815, MCOutput[58]}), .c ({new_AGEMA_signal_1869, AddKeyXOR1_XORInst_2_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_1871, AddKeyXOR1_XORInst_3_0_n1}), .b ({new_AGEMA_signal_4026, new_AGEMA_signal_4018}), .c ({new_AGEMA_signal_1903, AddRoundKeyOutput[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_3_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1819, MCOutput[60]}), .c ({new_AGEMA_signal_1871, AddKeyXOR1_XORInst_3_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_1873, AddKeyXOR1_XORInst_3_2_n1}), .b ({new_AGEMA_signal_4042, new_AGEMA_signal_4034}), .c ({new_AGEMA_signal_1905, AddRoundKeyOutput[62]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR1_XORInst_3_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1823, MCOutput[62]}), .c ({new_AGEMA_signal_1873, AddKeyXOR1_XORInst_3_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_0_U3 ( .a ({new_AGEMA_signal_1875, AddKeyConstXOR_XORInst_0_0_n2}), .b ({new_AGEMA_signal_4058, new_AGEMA_signal_4050}), .c ({new_AGEMA_signal_1907, AddRoundKeyOutput[40]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1812, MCOutput[40]}), .c ({new_AGEMA_signal_1875, AddKeyConstXOR_XORInst_0_0_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_2_U3 ( .a ({new_AGEMA_signal_1877, AddKeyConstXOR_XORInst_0_2_n2}), .b ({new_AGEMA_signal_4074, new_AGEMA_signal_4066}), .c ({new_AGEMA_signal_1909, AddRoundKeyOutput[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_0_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1816, MCOutput[42]}), .c ({new_AGEMA_signal_1877, AddKeyConstXOR_XORInst_0_2_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_0_U3 ( .a ({new_AGEMA_signal_1879, AddKeyConstXOR_XORInst_1_0_n2}), .b ({new_AGEMA_signal_4090, new_AGEMA_signal_4082}), .c ({new_AGEMA_signal_1911, AddRoundKeyOutput[44]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1820, MCOutput[44]}), .c ({new_AGEMA_signal_1879, AddKeyConstXOR_XORInst_1_0_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_2_U3 ( .a ({new_AGEMA_signal_1881, AddKeyConstXOR_XORInst_1_2_n2}), .b ({new_AGEMA_signal_4106, new_AGEMA_signal_4098}), .c ({new_AGEMA_signal_1913, AddRoundKeyOutput[46]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyConstXOR_XORInst_1_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1824, MCOutput[46]}), .c ({new_AGEMA_signal_1881, AddKeyConstXOR_XORInst_1_2_n2}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_1763, AddKeyXOR2_XORInst_0_0_n1}), .b ({new_AGEMA_signal_4122, new_AGEMA_signal_4114}), .c ({new_AGEMA_signal_1827, AddRoundKeyOutput[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_0_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1580, MCOutput[0]}), .c ({new_AGEMA_signal_1763, AddKeyXOR2_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_1765, AddKeyXOR2_XORInst_0_2_n1}), .b ({new_AGEMA_signal_4138, new_AGEMA_signal_4130}), .c ({new_AGEMA_signal_1829, AddRoundKeyOutput[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_0_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1584, MCOutput[2]}), .c ({new_AGEMA_signal_1765, AddKeyXOR2_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_1767, AddKeyXOR2_XORInst_1_0_n1}), .b ({new_AGEMA_signal_4154, new_AGEMA_signal_4146}), .c ({new_AGEMA_signal_1831, AddRoundKeyOutput[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_1_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1588, MCOutput[4]}), .c ({new_AGEMA_signal_1767, AddKeyXOR2_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_1769, AddKeyXOR2_XORInst_1_2_n1}), .b ({new_AGEMA_signal_4170, new_AGEMA_signal_4162}), .c ({new_AGEMA_signal_1833, AddRoundKeyOutput[6]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_1_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1592, MCOutput[6]}), .c ({new_AGEMA_signal_1769, AddKeyXOR2_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_1771, AddKeyXOR2_XORInst_2_0_n1}), .b ({new_AGEMA_signal_4186, new_AGEMA_signal_4178}), .c ({new_AGEMA_signal_1835, AddRoundKeyOutput[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_2_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1596, MCOutput[8]}), .c ({new_AGEMA_signal_1771, AddKeyXOR2_XORInst_2_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_1773, AddKeyXOR2_XORInst_2_2_n1}), .b ({new_AGEMA_signal_4202, new_AGEMA_signal_4194}), .c ({new_AGEMA_signal_1837, AddRoundKeyOutput[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_2_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1600, MCOutput[10]}), .c ({new_AGEMA_signal_1773, AddKeyXOR2_XORInst_2_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_1775, AddKeyXOR2_XORInst_3_0_n1}), .b ({new_AGEMA_signal_4218, new_AGEMA_signal_4210}), .c ({new_AGEMA_signal_1839, AddRoundKeyOutput[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_3_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1604, MCOutput[12]}), .c ({new_AGEMA_signal_1775, AddKeyXOR2_XORInst_3_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_1777, AddKeyXOR2_XORInst_3_2_n1}), .b ({new_AGEMA_signal_4234, new_AGEMA_signal_4226}), .c ({new_AGEMA_signal_1841, AddRoundKeyOutput[14]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_3_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1608, MCOutput[14]}), .c ({new_AGEMA_signal_1777, AddKeyXOR2_XORInst_3_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_4_0_U2 ( .a ({new_AGEMA_signal_1779, AddKeyXOR2_XORInst_4_0_n1}), .b ({new_AGEMA_signal_4250, new_AGEMA_signal_4242}), .c ({new_AGEMA_signal_1843, AddRoundKeyOutput[16]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_4_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1612, MCOutput[16]}), .c ({new_AGEMA_signal_1779, AddKeyXOR2_XORInst_4_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_4_2_U2 ( .a ({new_AGEMA_signal_1781, AddKeyXOR2_XORInst_4_2_n1}), .b ({new_AGEMA_signal_4266, new_AGEMA_signal_4258}), .c ({new_AGEMA_signal_1845, AddRoundKeyOutput[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_4_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1616, MCOutput[18]}), .c ({new_AGEMA_signal_1781, AddKeyXOR2_XORInst_4_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_5_0_U2 ( .a ({new_AGEMA_signal_1783, AddKeyXOR2_XORInst_5_0_n1}), .b ({new_AGEMA_signal_4282, new_AGEMA_signal_4274}), .c ({new_AGEMA_signal_1847, AddRoundKeyOutput[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_5_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1620, MCOutput[20]}), .c ({new_AGEMA_signal_1783, AddKeyXOR2_XORInst_5_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_5_2_U2 ( .a ({new_AGEMA_signal_1785, AddKeyXOR2_XORInst_5_2_n1}), .b ({new_AGEMA_signal_4298, new_AGEMA_signal_4290}), .c ({new_AGEMA_signal_1849, AddRoundKeyOutput[22]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_5_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1624, MCOutput[22]}), .c ({new_AGEMA_signal_1785, AddKeyXOR2_XORInst_5_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_6_0_U2 ( .a ({new_AGEMA_signal_1787, AddKeyXOR2_XORInst_6_0_n1}), .b ({new_AGEMA_signal_4314, new_AGEMA_signal_4306}), .c ({new_AGEMA_signal_1851, AddRoundKeyOutput[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_6_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1628, MCOutput[24]}), .c ({new_AGEMA_signal_1787, AddKeyXOR2_XORInst_6_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_6_2_U2 ( .a ({new_AGEMA_signal_1789, AddKeyXOR2_XORInst_6_2_n1}), .b ({new_AGEMA_signal_4330, new_AGEMA_signal_4322}), .c ({new_AGEMA_signal_1853, AddRoundKeyOutput[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_6_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1632, MCOutput[26]}), .c ({new_AGEMA_signal_1789, AddKeyXOR2_XORInst_6_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_7_0_U2 ( .a ({new_AGEMA_signal_1791, AddKeyXOR2_XORInst_7_0_n1}), .b ({new_AGEMA_signal_4346, new_AGEMA_signal_4338}), .c ({new_AGEMA_signal_1855, AddRoundKeyOutput[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_7_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1636, MCOutput[28]}), .c ({new_AGEMA_signal_1791, AddKeyXOR2_XORInst_7_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_7_2_U2 ( .a ({new_AGEMA_signal_1793, AddKeyXOR2_XORInst_7_2_n1}), .b ({new_AGEMA_signal_4362, new_AGEMA_signal_4354}), .c ({new_AGEMA_signal_1857, AddRoundKeyOutput[30]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_7_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1640, MCOutput[30]}), .c ({new_AGEMA_signal_1793, AddKeyXOR2_XORInst_7_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_8_0_U2 ( .a ({new_AGEMA_signal_1883, AddKeyXOR2_XORInst_8_0_n1}), .b ({new_AGEMA_signal_4378, new_AGEMA_signal_4370}), .c ({new_AGEMA_signal_1915, AddRoundKeyOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_8_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1796, MCOutput[32]}), .c ({new_AGEMA_signal_1883, AddKeyXOR2_XORInst_8_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_8_2_U2 ( .a ({new_AGEMA_signal_1885, AddKeyXOR2_XORInst_8_2_n1}), .b ({new_AGEMA_signal_4394, new_AGEMA_signal_4386}), .c ({new_AGEMA_signal_1917, AddRoundKeyOutput[34]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_8_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1800, MCOutput[34]}), .c ({new_AGEMA_signal_1885, AddKeyXOR2_XORInst_8_2_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_9_0_U2 ( .a ({new_AGEMA_signal_1887, AddKeyXOR2_XORInst_9_0_n1}), .b ({new_AGEMA_signal_4410, new_AGEMA_signal_4402}), .c ({new_AGEMA_signal_1919, AddRoundKeyOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_9_0_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1804, MCOutput[36]}), .c ({new_AGEMA_signal_1887, AddKeyXOR2_XORInst_9_0_n1}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_9_2_U2 ( .a ({new_AGEMA_signal_1889, AddKeyXOR2_XORInst_9_2_n1}), .b ({new_AGEMA_signal_4426, new_AGEMA_signal_4418}), .c ({new_AGEMA_signal_1921, AddRoundKeyOutput[38]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) AddKeyXOR2_XORInst_9_2_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1808, MCOutput[38]}), .c ({new_AGEMA_signal_1889, AddKeyXOR2_XORInst_9_2_n1}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U17 ( .a ({new_AGEMA_signal_4430, new_AGEMA_signal_4428}), .b ({new_AGEMA_signal_1293, SubCellInst_SboxInst_0_n12}), .clk (clk), .r (Fresh[224]), .c ({new_AGEMA_signal_1372, Feedback[2]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_0_U8 ( .a ({new_AGEMA_signal_4438, new_AGEMA_signal_4434}), .b ({new_AGEMA_signal_1295, SubCellInst_SboxInst_0_n3}), .clk (clk), .r (Fresh[225]), .c ({new_AGEMA_signal_1374, Feedback[0]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U17 ( .a ({new_AGEMA_signal_4442, new_AGEMA_signal_4440}), .b ({new_AGEMA_signal_1298, SubCellInst_SboxInst_1_n12}), .clk (clk), .r (Fresh[226]), .c ({new_AGEMA_signal_1376, Feedback[6]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_1_U8 ( .a ({new_AGEMA_signal_4450, new_AGEMA_signal_4446}), .b ({new_AGEMA_signal_1300, SubCellInst_SboxInst_1_n3}), .clk (clk), .r (Fresh[227]), .c ({new_AGEMA_signal_1378, Feedback[4]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U17 ( .a ({new_AGEMA_signal_4454, new_AGEMA_signal_4452}), .b ({new_AGEMA_signal_1303, SubCellInst_SboxInst_2_n12}), .clk (clk), .r (Fresh[228]), .c ({new_AGEMA_signal_1380, Feedback[10]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_2_U8 ( .a ({new_AGEMA_signal_4462, new_AGEMA_signal_4458}), .b ({new_AGEMA_signal_1305, SubCellInst_SboxInst_2_n3}), .clk (clk), .r (Fresh[229]), .c ({new_AGEMA_signal_1382, Feedback[8]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U17 ( .a ({new_AGEMA_signal_4466, new_AGEMA_signal_4464}), .b ({new_AGEMA_signal_1308, SubCellInst_SboxInst_3_n12}), .clk (clk), .r (Fresh[230]), .c ({new_AGEMA_signal_1384, Feedback[14]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_3_U8 ( .a ({new_AGEMA_signal_4474, new_AGEMA_signal_4470}), .b ({new_AGEMA_signal_1310, SubCellInst_SboxInst_3_n3}), .clk (clk), .r (Fresh[231]), .c ({new_AGEMA_signal_1386, Feedback[12]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U17 ( .a ({new_AGEMA_signal_4478, new_AGEMA_signal_4476}), .b ({new_AGEMA_signal_1313, SubCellInst_SboxInst_4_n12}), .clk (clk), .r (Fresh[232]), .c ({new_AGEMA_signal_1388, Feedback[18]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_4_U8 ( .a ({new_AGEMA_signal_4486, new_AGEMA_signal_4482}), .b ({new_AGEMA_signal_1315, SubCellInst_SboxInst_4_n3}), .clk (clk), .r (Fresh[233]), .c ({new_AGEMA_signal_1390, Feedback[16]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U17 ( .a ({new_AGEMA_signal_4490, new_AGEMA_signal_4488}), .b ({new_AGEMA_signal_1318, SubCellInst_SboxInst_5_n12}), .clk (clk), .r (Fresh[234]), .c ({new_AGEMA_signal_1392, Feedback[22]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_5_U8 ( .a ({new_AGEMA_signal_4498, new_AGEMA_signal_4494}), .b ({new_AGEMA_signal_1320, SubCellInst_SboxInst_5_n3}), .clk (clk), .r (Fresh[235]), .c ({new_AGEMA_signal_1394, Feedback[20]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U17 ( .a ({new_AGEMA_signal_4502, new_AGEMA_signal_4500}), .b ({new_AGEMA_signal_1323, SubCellInst_SboxInst_6_n12}), .clk (clk), .r (Fresh[236]), .c ({new_AGEMA_signal_1396, Feedback[26]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_6_U8 ( .a ({new_AGEMA_signal_4510, new_AGEMA_signal_4506}), .b ({new_AGEMA_signal_1325, SubCellInst_SboxInst_6_n3}), .clk (clk), .r (Fresh[237]), .c ({new_AGEMA_signal_1398, Feedback[24]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U17 ( .a ({new_AGEMA_signal_4514, new_AGEMA_signal_4512}), .b ({new_AGEMA_signal_1328, SubCellInst_SboxInst_7_n12}), .clk (clk), .r (Fresh[238]), .c ({new_AGEMA_signal_1400, Feedback[30]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_7_U8 ( .a ({new_AGEMA_signal_4522, new_AGEMA_signal_4518}), .b ({new_AGEMA_signal_1330, SubCellInst_SboxInst_7_n3}), .clk (clk), .r (Fresh[239]), .c ({new_AGEMA_signal_1402, Feedback[28]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U17 ( .a ({new_AGEMA_signal_4526, new_AGEMA_signal_4524}), .b ({new_AGEMA_signal_1333, SubCellInst_SboxInst_8_n12}), .clk (clk), .r (Fresh[240]), .c ({new_AGEMA_signal_1404, Feedback[34]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_8_U8 ( .a ({new_AGEMA_signal_4534, new_AGEMA_signal_4530}), .b ({new_AGEMA_signal_1335, SubCellInst_SboxInst_8_n3}), .clk (clk), .r (Fresh[241]), .c ({new_AGEMA_signal_1406, Feedback[32]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U17 ( .a ({new_AGEMA_signal_4538, new_AGEMA_signal_4536}), .b ({new_AGEMA_signal_1338, SubCellInst_SboxInst_9_n12}), .clk (clk), .r (Fresh[242]), .c ({new_AGEMA_signal_1408, Feedback[38]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_9_U8 ( .a ({new_AGEMA_signal_4546, new_AGEMA_signal_4542}), .b ({new_AGEMA_signal_1340, SubCellInst_SboxInst_9_n3}), .clk (clk), .r (Fresh[243]), .c ({new_AGEMA_signal_1410, Feedback[36]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U17 ( .a ({new_AGEMA_signal_4550, new_AGEMA_signal_4548}), .b ({new_AGEMA_signal_1343, SubCellInst_SboxInst_10_n12}), .clk (clk), .r (Fresh[244]), .c ({new_AGEMA_signal_1412, Feedback[42]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_10_U8 ( .a ({new_AGEMA_signal_4558, new_AGEMA_signal_4554}), .b ({new_AGEMA_signal_1345, SubCellInst_SboxInst_10_n3}), .clk (clk), .r (Fresh[245]), .c ({new_AGEMA_signal_1414, Feedback[40]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U17 ( .a ({new_AGEMA_signal_4562, new_AGEMA_signal_4560}), .b ({new_AGEMA_signal_1348, SubCellInst_SboxInst_11_n12}), .clk (clk), .r (Fresh[246]), .c ({new_AGEMA_signal_1416, Feedback[46]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_11_U8 ( .a ({new_AGEMA_signal_4570, new_AGEMA_signal_4566}), .b ({new_AGEMA_signal_1350, SubCellInst_SboxInst_11_n3}), .clk (clk), .r (Fresh[247]), .c ({new_AGEMA_signal_1418, Feedback[44]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U17 ( .a ({new_AGEMA_signal_4574, new_AGEMA_signal_4572}), .b ({new_AGEMA_signal_1353, SubCellInst_SboxInst_12_n12}), .clk (clk), .r (Fresh[248]), .c ({new_AGEMA_signal_1420, Feedback[50]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_12_U8 ( .a ({new_AGEMA_signal_4582, new_AGEMA_signal_4578}), .b ({new_AGEMA_signal_1355, SubCellInst_SboxInst_12_n3}), .clk (clk), .r (Fresh[249]), .c ({new_AGEMA_signal_1422, Feedback[48]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U17 ( .a ({new_AGEMA_signal_4586, new_AGEMA_signal_4584}), .b ({new_AGEMA_signal_1358, SubCellInst_SboxInst_13_n12}), .clk (clk), .r (Fresh[250]), .c ({new_AGEMA_signal_1424, Feedback[54]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_13_U8 ( .a ({new_AGEMA_signal_4594, new_AGEMA_signal_4590}), .b ({new_AGEMA_signal_1360, SubCellInst_SboxInst_13_n3}), .clk (clk), .r (Fresh[251]), .c ({new_AGEMA_signal_1426, Feedback[52]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U17 ( .a ({new_AGEMA_signal_4598, new_AGEMA_signal_4596}), .b ({new_AGEMA_signal_1363, SubCellInst_SboxInst_14_n12}), .clk (clk), .r (Fresh[252]), .c ({new_AGEMA_signal_1428, Feedback[58]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_14_U8 ( .a ({new_AGEMA_signal_4606, new_AGEMA_signal_4602}), .b ({new_AGEMA_signal_1365, SubCellInst_SboxInst_14_n3}), .clk (clk), .r (Fresh[253]), .c ({new_AGEMA_signal_1430, Feedback[56]}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U17 ( .a ({new_AGEMA_signal_4610, new_AGEMA_signal_4608}), .b ({new_AGEMA_signal_1368, SubCellInst_SboxInst_15_n12}), .clk (clk), .r (Fresh[254]), .c ({new_AGEMA_signal_1432, Feedback[62]}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) SubCellInst_SboxInst_15_U8 ( .a ({new_AGEMA_signal_4618, new_AGEMA_signal_4614}), .b ({new_AGEMA_signal_1370, SubCellInst_SboxInst_15_n3}), .clk (clk), .r (Fresh[255]), .c ({new_AGEMA_signal_1434, Feedback[60]}) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C (clk), .D (new_AGEMA_signal_3401), .Q (new_AGEMA_signal_3402) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C (clk), .D (new_AGEMA_signal_3409), .Q (new_AGEMA_signal_3410) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C (clk), .D (new_AGEMA_signal_3417), .Q (new_AGEMA_signal_3418) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C (clk), .D (new_AGEMA_signal_3425), .Q (new_AGEMA_signal_3426) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C (clk), .D (new_AGEMA_signal_3433), .Q (new_AGEMA_signal_3434) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C (clk), .D (new_AGEMA_signal_3441), .Q (new_AGEMA_signal_3442) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C (clk), .D (new_AGEMA_signal_3449), .Q (new_AGEMA_signal_3450) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C (clk), .D (new_AGEMA_signal_3457), .Q (new_AGEMA_signal_3458) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C (clk), .D (new_AGEMA_signal_3465), .Q (new_AGEMA_signal_3466) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C (clk), .D (new_AGEMA_signal_3473), .Q (new_AGEMA_signal_3474) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C (clk), .D (new_AGEMA_signal_3481), .Q (new_AGEMA_signal_3482) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C (clk), .D (new_AGEMA_signal_3489), .Q (new_AGEMA_signal_3490) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C (clk), .D (new_AGEMA_signal_3497), .Q (new_AGEMA_signal_3498) ) ;
    buf_clk new_AGEMA_reg_buffer_2146 ( .C (clk), .D (new_AGEMA_signal_3505), .Q (new_AGEMA_signal_3506) ) ;
    buf_clk new_AGEMA_reg_buffer_2154 ( .C (clk), .D (new_AGEMA_signal_3513), .Q (new_AGEMA_signal_3514) ) ;
    buf_clk new_AGEMA_reg_buffer_2162 ( .C (clk), .D (new_AGEMA_signal_3521), .Q (new_AGEMA_signal_3522) ) ;
    buf_clk new_AGEMA_reg_buffer_2170 ( .C (clk), .D (new_AGEMA_signal_3529), .Q (new_AGEMA_signal_3530) ) ;
    buf_clk new_AGEMA_reg_buffer_2178 ( .C (clk), .D (new_AGEMA_signal_3537), .Q (new_AGEMA_signal_3538) ) ;
    buf_clk new_AGEMA_reg_buffer_2186 ( .C (clk), .D (new_AGEMA_signal_3545), .Q (new_AGEMA_signal_3546) ) ;
    buf_clk new_AGEMA_reg_buffer_2194 ( .C (clk), .D (new_AGEMA_signal_3553), .Q (new_AGEMA_signal_3554) ) ;
    buf_clk new_AGEMA_reg_buffer_2202 ( .C (clk), .D (new_AGEMA_signal_3561), .Q (new_AGEMA_signal_3562) ) ;
    buf_clk new_AGEMA_reg_buffer_2210 ( .C (clk), .D (new_AGEMA_signal_3569), .Q (new_AGEMA_signal_3570) ) ;
    buf_clk new_AGEMA_reg_buffer_2218 ( .C (clk), .D (new_AGEMA_signal_3577), .Q (new_AGEMA_signal_3578) ) ;
    buf_clk new_AGEMA_reg_buffer_2226 ( .C (clk), .D (new_AGEMA_signal_3585), .Q (new_AGEMA_signal_3586) ) ;
    buf_clk new_AGEMA_reg_buffer_2234 ( .C (clk), .D (new_AGEMA_signal_3593), .Q (new_AGEMA_signal_3594) ) ;
    buf_clk new_AGEMA_reg_buffer_2242 ( .C (clk), .D (new_AGEMA_signal_3601), .Q (new_AGEMA_signal_3602) ) ;
    buf_clk new_AGEMA_reg_buffer_2250 ( .C (clk), .D (new_AGEMA_signal_3609), .Q (new_AGEMA_signal_3610) ) ;
    buf_clk new_AGEMA_reg_buffer_2258 ( .C (clk), .D (new_AGEMA_signal_3617), .Q (new_AGEMA_signal_3618) ) ;
    buf_clk new_AGEMA_reg_buffer_2266 ( .C (clk), .D (new_AGEMA_signal_3625), .Q (new_AGEMA_signal_3626) ) ;
    buf_clk new_AGEMA_reg_buffer_2274 ( .C (clk), .D (new_AGEMA_signal_3633), .Q (new_AGEMA_signal_3634) ) ;
    buf_clk new_AGEMA_reg_buffer_2282 ( .C (clk), .D (new_AGEMA_signal_3641), .Q (new_AGEMA_signal_3642) ) ;
    buf_clk new_AGEMA_reg_buffer_2290 ( .C (clk), .D (new_AGEMA_signal_3649), .Q (new_AGEMA_signal_3650) ) ;
    buf_clk new_AGEMA_reg_buffer_2298 ( .C (clk), .D (new_AGEMA_signal_3657), .Q (new_AGEMA_signal_3658) ) ;
    buf_clk new_AGEMA_reg_buffer_2306 ( .C (clk), .D (new_AGEMA_signal_3665), .Q (new_AGEMA_signal_3666) ) ;
    buf_clk new_AGEMA_reg_buffer_2314 ( .C (clk), .D (new_AGEMA_signal_3673), .Q (new_AGEMA_signal_3674) ) ;
    buf_clk new_AGEMA_reg_buffer_2322 ( .C (clk), .D (new_AGEMA_signal_3681), .Q (new_AGEMA_signal_3682) ) ;
    buf_clk new_AGEMA_reg_buffer_2330 ( .C (clk), .D (new_AGEMA_signal_3689), .Q (new_AGEMA_signal_3690) ) ;
    buf_clk new_AGEMA_reg_buffer_2338 ( .C (clk), .D (new_AGEMA_signal_3697), .Q (new_AGEMA_signal_3698) ) ;
    buf_clk new_AGEMA_reg_buffer_2346 ( .C (clk), .D (new_AGEMA_signal_3705), .Q (new_AGEMA_signal_3706) ) ;
    buf_clk new_AGEMA_reg_buffer_2354 ( .C (clk), .D (new_AGEMA_signal_3713), .Q (new_AGEMA_signal_3714) ) ;
    buf_clk new_AGEMA_reg_buffer_2362 ( .C (clk), .D (new_AGEMA_signal_3721), .Q (new_AGEMA_signal_3722) ) ;
    buf_clk new_AGEMA_reg_buffer_2370 ( .C (clk), .D (new_AGEMA_signal_3729), .Q (new_AGEMA_signal_3730) ) ;
    buf_clk new_AGEMA_reg_buffer_2378 ( .C (clk), .D (new_AGEMA_signal_3737), .Q (new_AGEMA_signal_3738) ) ;
    buf_clk new_AGEMA_reg_buffer_2386 ( .C (clk), .D (new_AGEMA_signal_3745), .Q (new_AGEMA_signal_3746) ) ;
    buf_clk new_AGEMA_reg_buffer_2394 ( .C (clk), .D (new_AGEMA_signal_3753), .Q (new_AGEMA_signal_3754) ) ;
    buf_clk new_AGEMA_reg_buffer_2402 ( .C (clk), .D (new_AGEMA_signal_3761), .Q (new_AGEMA_signal_3762) ) ;
    buf_clk new_AGEMA_reg_buffer_2410 ( .C (clk), .D (new_AGEMA_signal_3769), .Q (new_AGEMA_signal_3770) ) ;
    buf_clk new_AGEMA_reg_buffer_2418 ( .C (clk), .D (new_AGEMA_signal_3777), .Q (new_AGEMA_signal_3778) ) ;
    buf_clk new_AGEMA_reg_buffer_2426 ( .C (clk), .D (new_AGEMA_signal_3785), .Q (new_AGEMA_signal_3786) ) ;
    buf_clk new_AGEMA_reg_buffer_2434 ( .C (clk), .D (new_AGEMA_signal_3793), .Q (new_AGEMA_signal_3794) ) ;
    buf_clk new_AGEMA_reg_buffer_2442 ( .C (clk), .D (new_AGEMA_signal_3801), .Q (new_AGEMA_signal_3802) ) ;
    buf_clk new_AGEMA_reg_buffer_2450 ( .C (clk), .D (new_AGEMA_signal_3809), .Q (new_AGEMA_signal_3810) ) ;
    buf_clk new_AGEMA_reg_buffer_2458 ( .C (clk), .D (new_AGEMA_signal_3817), .Q (new_AGEMA_signal_3818) ) ;
    buf_clk new_AGEMA_reg_buffer_2466 ( .C (clk), .D (new_AGEMA_signal_3825), .Q (new_AGEMA_signal_3826) ) ;
    buf_clk new_AGEMA_reg_buffer_2474 ( .C (clk), .D (new_AGEMA_signal_3833), .Q (new_AGEMA_signal_3834) ) ;
    buf_clk new_AGEMA_reg_buffer_2482 ( .C (clk), .D (new_AGEMA_signal_3841), .Q (new_AGEMA_signal_3842) ) ;
    buf_clk new_AGEMA_reg_buffer_2490 ( .C (clk), .D (new_AGEMA_signal_3849), .Q (new_AGEMA_signal_3850) ) ;
    buf_clk new_AGEMA_reg_buffer_2498 ( .C (clk), .D (new_AGEMA_signal_3857), .Q (new_AGEMA_signal_3858) ) ;
    buf_clk new_AGEMA_reg_buffer_2506 ( .C (clk), .D (new_AGEMA_signal_3865), .Q (new_AGEMA_signal_3866) ) ;
    buf_clk new_AGEMA_reg_buffer_2514 ( .C (clk), .D (new_AGEMA_signal_3873), .Q (new_AGEMA_signal_3874) ) ;
    buf_clk new_AGEMA_reg_buffer_2522 ( .C (clk), .D (new_AGEMA_signal_3881), .Q (new_AGEMA_signal_3882) ) ;
    buf_clk new_AGEMA_reg_buffer_2530 ( .C (clk), .D (new_AGEMA_signal_3889), .Q (new_AGEMA_signal_3890) ) ;
    buf_clk new_AGEMA_reg_buffer_2538 ( .C (clk), .D (new_AGEMA_signal_3897), .Q (new_AGEMA_signal_3898) ) ;
    buf_clk new_AGEMA_reg_buffer_2546 ( .C (clk), .D (new_AGEMA_signal_3905), .Q (new_AGEMA_signal_3906) ) ;
    buf_clk new_AGEMA_reg_buffer_2554 ( .C (clk), .D (new_AGEMA_signal_3913), .Q (new_AGEMA_signal_3914) ) ;
    buf_clk new_AGEMA_reg_buffer_2562 ( .C (clk), .D (new_AGEMA_signal_3921), .Q (new_AGEMA_signal_3922) ) ;
    buf_clk new_AGEMA_reg_buffer_2570 ( .C (clk), .D (new_AGEMA_signal_3929), .Q (new_AGEMA_signal_3930) ) ;
    buf_clk new_AGEMA_reg_buffer_2578 ( .C (clk), .D (new_AGEMA_signal_3937), .Q (new_AGEMA_signal_3938) ) ;
    buf_clk new_AGEMA_reg_buffer_2586 ( .C (clk), .D (new_AGEMA_signal_3945), .Q (new_AGEMA_signal_3946) ) ;
    buf_clk new_AGEMA_reg_buffer_2594 ( .C (clk), .D (new_AGEMA_signal_3953), .Q (new_AGEMA_signal_3954) ) ;
    buf_clk new_AGEMA_reg_buffer_2602 ( .C (clk), .D (new_AGEMA_signal_3961), .Q (new_AGEMA_signal_3962) ) ;
    buf_clk new_AGEMA_reg_buffer_2610 ( .C (clk), .D (new_AGEMA_signal_3969), .Q (new_AGEMA_signal_3970) ) ;
    buf_clk new_AGEMA_reg_buffer_2618 ( .C (clk), .D (new_AGEMA_signal_3977), .Q (new_AGEMA_signal_3978) ) ;
    buf_clk new_AGEMA_reg_buffer_2626 ( .C (clk), .D (new_AGEMA_signal_3985), .Q (new_AGEMA_signal_3986) ) ;
    buf_clk new_AGEMA_reg_buffer_2634 ( .C (clk), .D (new_AGEMA_signal_3993), .Q (new_AGEMA_signal_3994) ) ;
    buf_clk new_AGEMA_reg_buffer_2642 ( .C (clk), .D (new_AGEMA_signal_4001), .Q (new_AGEMA_signal_4002) ) ;
    buf_clk new_AGEMA_reg_buffer_2650 ( .C (clk), .D (new_AGEMA_signal_4009), .Q (new_AGEMA_signal_4010) ) ;
    buf_clk new_AGEMA_reg_buffer_2658 ( .C (clk), .D (new_AGEMA_signal_4017), .Q (new_AGEMA_signal_4018) ) ;
    buf_clk new_AGEMA_reg_buffer_2666 ( .C (clk), .D (new_AGEMA_signal_4025), .Q (new_AGEMA_signal_4026) ) ;
    buf_clk new_AGEMA_reg_buffer_2674 ( .C (clk), .D (new_AGEMA_signal_4033), .Q (new_AGEMA_signal_4034) ) ;
    buf_clk new_AGEMA_reg_buffer_2682 ( .C (clk), .D (new_AGEMA_signal_4041), .Q (new_AGEMA_signal_4042) ) ;
    buf_clk new_AGEMA_reg_buffer_2690 ( .C (clk), .D (new_AGEMA_signal_4049), .Q (new_AGEMA_signal_4050) ) ;
    buf_clk new_AGEMA_reg_buffer_2698 ( .C (clk), .D (new_AGEMA_signal_4057), .Q (new_AGEMA_signal_4058) ) ;
    buf_clk new_AGEMA_reg_buffer_2706 ( .C (clk), .D (new_AGEMA_signal_4065), .Q (new_AGEMA_signal_4066) ) ;
    buf_clk new_AGEMA_reg_buffer_2714 ( .C (clk), .D (new_AGEMA_signal_4073), .Q (new_AGEMA_signal_4074) ) ;
    buf_clk new_AGEMA_reg_buffer_2722 ( .C (clk), .D (new_AGEMA_signal_4081), .Q (new_AGEMA_signal_4082) ) ;
    buf_clk new_AGEMA_reg_buffer_2730 ( .C (clk), .D (new_AGEMA_signal_4089), .Q (new_AGEMA_signal_4090) ) ;
    buf_clk new_AGEMA_reg_buffer_2738 ( .C (clk), .D (new_AGEMA_signal_4097), .Q (new_AGEMA_signal_4098) ) ;
    buf_clk new_AGEMA_reg_buffer_2746 ( .C (clk), .D (new_AGEMA_signal_4105), .Q (new_AGEMA_signal_4106) ) ;
    buf_clk new_AGEMA_reg_buffer_2754 ( .C (clk), .D (new_AGEMA_signal_4113), .Q (new_AGEMA_signal_4114) ) ;
    buf_clk new_AGEMA_reg_buffer_2762 ( .C (clk), .D (new_AGEMA_signal_4121), .Q (new_AGEMA_signal_4122) ) ;
    buf_clk new_AGEMA_reg_buffer_2770 ( .C (clk), .D (new_AGEMA_signal_4129), .Q (new_AGEMA_signal_4130) ) ;
    buf_clk new_AGEMA_reg_buffer_2778 ( .C (clk), .D (new_AGEMA_signal_4137), .Q (new_AGEMA_signal_4138) ) ;
    buf_clk new_AGEMA_reg_buffer_2786 ( .C (clk), .D (new_AGEMA_signal_4145), .Q (new_AGEMA_signal_4146) ) ;
    buf_clk new_AGEMA_reg_buffer_2794 ( .C (clk), .D (new_AGEMA_signal_4153), .Q (new_AGEMA_signal_4154) ) ;
    buf_clk new_AGEMA_reg_buffer_2802 ( .C (clk), .D (new_AGEMA_signal_4161), .Q (new_AGEMA_signal_4162) ) ;
    buf_clk new_AGEMA_reg_buffer_2810 ( .C (clk), .D (new_AGEMA_signal_4169), .Q (new_AGEMA_signal_4170) ) ;
    buf_clk new_AGEMA_reg_buffer_2818 ( .C (clk), .D (new_AGEMA_signal_4177), .Q (new_AGEMA_signal_4178) ) ;
    buf_clk new_AGEMA_reg_buffer_2826 ( .C (clk), .D (new_AGEMA_signal_4185), .Q (new_AGEMA_signal_4186) ) ;
    buf_clk new_AGEMA_reg_buffer_2834 ( .C (clk), .D (new_AGEMA_signal_4193), .Q (new_AGEMA_signal_4194) ) ;
    buf_clk new_AGEMA_reg_buffer_2842 ( .C (clk), .D (new_AGEMA_signal_4201), .Q (new_AGEMA_signal_4202) ) ;
    buf_clk new_AGEMA_reg_buffer_2850 ( .C (clk), .D (new_AGEMA_signal_4209), .Q (new_AGEMA_signal_4210) ) ;
    buf_clk new_AGEMA_reg_buffer_2858 ( .C (clk), .D (new_AGEMA_signal_4217), .Q (new_AGEMA_signal_4218) ) ;
    buf_clk new_AGEMA_reg_buffer_2866 ( .C (clk), .D (new_AGEMA_signal_4225), .Q (new_AGEMA_signal_4226) ) ;
    buf_clk new_AGEMA_reg_buffer_2874 ( .C (clk), .D (new_AGEMA_signal_4233), .Q (new_AGEMA_signal_4234) ) ;
    buf_clk new_AGEMA_reg_buffer_2882 ( .C (clk), .D (new_AGEMA_signal_4241), .Q (new_AGEMA_signal_4242) ) ;
    buf_clk new_AGEMA_reg_buffer_2890 ( .C (clk), .D (new_AGEMA_signal_4249), .Q (new_AGEMA_signal_4250) ) ;
    buf_clk new_AGEMA_reg_buffer_2898 ( .C (clk), .D (new_AGEMA_signal_4257), .Q (new_AGEMA_signal_4258) ) ;
    buf_clk new_AGEMA_reg_buffer_2906 ( .C (clk), .D (new_AGEMA_signal_4265), .Q (new_AGEMA_signal_4266) ) ;
    buf_clk new_AGEMA_reg_buffer_2914 ( .C (clk), .D (new_AGEMA_signal_4273), .Q (new_AGEMA_signal_4274) ) ;
    buf_clk new_AGEMA_reg_buffer_2922 ( .C (clk), .D (new_AGEMA_signal_4281), .Q (new_AGEMA_signal_4282) ) ;
    buf_clk new_AGEMA_reg_buffer_2930 ( .C (clk), .D (new_AGEMA_signal_4289), .Q (new_AGEMA_signal_4290) ) ;
    buf_clk new_AGEMA_reg_buffer_2938 ( .C (clk), .D (new_AGEMA_signal_4297), .Q (new_AGEMA_signal_4298) ) ;
    buf_clk new_AGEMA_reg_buffer_2946 ( .C (clk), .D (new_AGEMA_signal_4305), .Q (new_AGEMA_signal_4306) ) ;
    buf_clk new_AGEMA_reg_buffer_2954 ( .C (clk), .D (new_AGEMA_signal_4313), .Q (new_AGEMA_signal_4314) ) ;
    buf_clk new_AGEMA_reg_buffer_2962 ( .C (clk), .D (new_AGEMA_signal_4321), .Q (new_AGEMA_signal_4322) ) ;
    buf_clk new_AGEMA_reg_buffer_2970 ( .C (clk), .D (new_AGEMA_signal_4329), .Q (new_AGEMA_signal_4330) ) ;
    buf_clk new_AGEMA_reg_buffer_2978 ( .C (clk), .D (new_AGEMA_signal_4337), .Q (new_AGEMA_signal_4338) ) ;
    buf_clk new_AGEMA_reg_buffer_2986 ( .C (clk), .D (new_AGEMA_signal_4345), .Q (new_AGEMA_signal_4346) ) ;
    buf_clk new_AGEMA_reg_buffer_2994 ( .C (clk), .D (new_AGEMA_signal_4353), .Q (new_AGEMA_signal_4354) ) ;
    buf_clk new_AGEMA_reg_buffer_3002 ( .C (clk), .D (new_AGEMA_signal_4361), .Q (new_AGEMA_signal_4362) ) ;
    buf_clk new_AGEMA_reg_buffer_3010 ( .C (clk), .D (new_AGEMA_signal_4369), .Q (new_AGEMA_signal_4370) ) ;
    buf_clk new_AGEMA_reg_buffer_3018 ( .C (clk), .D (new_AGEMA_signal_4377), .Q (new_AGEMA_signal_4378) ) ;
    buf_clk new_AGEMA_reg_buffer_3026 ( .C (clk), .D (new_AGEMA_signal_4385), .Q (new_AGEMA_signal_4386) ) ;
    buf_clk new_AGEMA_reg_buffer_3034 ( .C (clk), .D (new_AGEMA_signal_4393), .Q (new_AGEMA_signal_4394) ) ;
    buf_clk new_AGEMA_reg_buffer_3042 ( .C (clk), .D (new_AGEMA_signal_4401), .Q (new_AGEMA_signal_4402) ) ;
    buf_clk new_AGEMA_reg_buffer_3050 ( .C (clk), .D (new_AGEMA_signal_4409), .Q (new_AGEMA_signal_4410) ) ;
    buf_clk new_AGEMA_reg_buffer_3058 ( .C (clk), .D (new_AGEMA_signal_4417), .Q (new_AGEMA_signal_4418) ) ;
    buf_clk new_AGEMA_reg_buffer_3066 ( .C (clk), .D (new_AGEMA_signal_4425), .Q (new_AGEMA_signal_4426) ) ;
    buf_clk new_AGEMA_reg_buffer_3260 ( .C (clk), .D (new_AGEMA_signal_4619), .Q (new_AGEMA_signal_4620) ) ;
    buf_clk new_AGEMA_reg_buffer_3262 ( .C (clk), .D (new_AGEMA_signal_4621), .Q (new_AGEMA_signal_4622) ) ;
    buf_clk new_AGEMA_reg_buffer_3264 ( .C (clk), .D (new_AGEMA_signal_4623), .Q (new_AGEMA_signal_4624) ) ;
    buf_clk new_AGEMA_reg_buffer_3266 ( .C (clk), .D (new_AGEMA_signal_4625), .Q (new_AGEMA_signal_4626) ) ;
    buf_clk new_AGEMA_reg_buffer_3268 ( .C (clk), .D (new_AGEMA_signal_4627), .Q (new_AGEMA_signal_4628) ) ;
    buf_clk new_AGEMA_reg_buffer_3270 ( .C (clk), .D (new_AGEMA_signal_4629), .Q (new_AGEMA_signal_4630) ) ;
    buf_clk new_AGEMA_reg_buffer_3272 ( .C (clk), .D (new_AGEMA_signal_4631), .Q (new_AGEMA_signal_4632) ) ;
    buf_clk new_AGEMA_reg_buffer_3274 ( .C (clk), .D (new_AGEMA_signal_4633), .Q (new_AGEMA_signal_4634) ) ;
    buf_clk new_AGEMA_reg_buffer_3276 ( .C (clk), .D (new_AGEMA_signal_4635), .Q (new_AGEMA_signal_4636) ) ;
    buf_clk new_AGEMA_reg_buffer_3278 ( .C (clk), .D (new_AGEMA_signal_4637), .Q (new_AGEMA_signal_4638) ) ;
    buf_clk new_AGEMA_reg_buffer_3280 ( .C (clk), .D (new_AGEMA_signal_4639), .Q (new_AGEMA_signal_4640) ) ;
    buf_clk new_AGEMA_reg_buffer_3282 ( .C (clk), .D (new_AGEMA_signal_4641), .Q (new_AGEMA_signal_4642) ) ;
    buf_clk new_AGEMA_reg_buffer_3284 ( .C (clk), .D (new_AGEMA_signal_4643), .Q (new_AGEMA_signal_4644) ) ;
    buf_clk new_AGEMA_reg_buffer_3286 ( .C (clk), .D (new_AGEMA_signal_4645), .Q (new_AGEMA_signal_4646) ) ;
    buf_clk new_AGEMA_reg_buffer_3288 ( .C (clk), .D (new_AGEMA_signal_4647), .Q (new_AGEMA_signal_4648) ) ;
    buf_clk new_AGEMA_reg_buffer_3290 ( .C (clk), .D (new_AGEMA_signal_4649), .Q (new_AGEMA_signal_4650) ) ;
    buf_clk new_AGEMA_reg_buffer_3292 ( .C (clk), .D (new_AGEMA_signal_4651), .Q (new_AGEMA_signal_4652) ) ;
    buf_clk new_AGEMA_reg_buffer_3294 ( .C (clk), .D (new_AGEMA_signal_4653), .Q (new_AGEMA_signal_4654) ) ;
    buf_clk new_AGEMA_reg_buffer_3296 ( .C (clk), .D (new_AGEMA_signal_4655), .Q (new_AGEMA_signal_4656) ) ;
    buf_clk new_AGEMA_reg_buffer_3298 ( .C (clk), .D (new_AGEMA_signal_4657), .Q (new_AGEMA_signal_4658) ) ;
    buf_clk new_AGEMA_reg_buffer_3300 ( .C (clk), .D (new_AGEMA_signal_4659), .Q (new_AGEMA_signal_4660) ) ;
    buf_clk new_AGEMA_reg_buffer_3302 ( .C (clk), .D (new_AGEMA_signal_4661), .Q (new_AGEMA_signal_4662) ) ;
    buf_clk new_AGEMA_reg_buffer_3304 ( .C (clk), .D (new_AGEMA_signal_4663), .Q (new_AGEMA_signal_4664) ) ;
    buf_clk new_AGEMA_reg_buffer_3306 ( .C (clk), .D (new_AGEMA_signal_4665), .Q (new_AGEMA_signal_4666) ) ;
    buf_clk new_AGEMA_reg_buffer_3308 ( .C (clk), .D (new_AGEMA_signal_4667), .Q (new_AGEMA_signal_4668) ) ;
    buf_clk new_AGEMA_reg_buffer_3310 ( .C (clk), .D (new_AGEMA_signal_4669), .Q (new_AGEMA_signal_4670) ) ;
    buf_clk new_AGEMA_reg_buffer_3312 ( .C (clk), .D (new_AGEMA_signal_4671), .Q (new_AGEMA_signal_4672) ) ;
    buf_clk new_AGEMA_reg_buffer_3314 ( .C (clk), .D (new_AGEMA_signal_4673), .Q (new_AGEMA_signal_4674) ) ;
    buf_clk new_AGEMA_reg_buffer_3316 ( .C (clk), .D (new_AGEMA_signal_4675), .Q (new_AGEMA_signal_4676) ) ;
    buf_clk new_AGEMA_reg_buffer_3318 ( .C (clk), .D (new_AGEMA_signal_4677), .Q (new_AGEMA_signal_4678) ) ;
    buf_clk new_AGEMA_reg_buffer_3320 ( .C (clk), .D (new_AGEMA_signal_4679), .Q (new_AGEMA_signal_4680) ) ;
    buf_clk new_AGEMA_reg_buffer_3322 ( .C (clk), .D (new_AGEMA_signal_4681), .Q (new_AGEMA_signal_4682) ) ;
    buf_clk new_AGEMA_reg_buffer_3324 ( .C (clk), .D (new_AGEMA_signal_4683), .Q (new_AGEMA_signal_4684) ) ;
    buf_clk new_AGEMA_reg_buffer_3326 ( .C (clk), .D (new_AGEMA_signal_4685), .Q (new_AGEMA_signal_4686) ) ;
    buf_clk new_AGEMA_reg_buffer_3328 ( .C (clk), .D (new_AGEMA_signal_4687), .Q (new_AGEMA_signal_4688) ) ;
    buf_clk new_AGEMA_reg_buffer_3330 ( .C (clk), .D (new_AGEMA_signal_4689), .Q (new_AGEMA_signal_4690) ) ;
    buf_clk new_AGEMA_reg_buffer_3332 ( .C (clk), .D (new_AGEMA_signal_4691), .Q (new_AGEMA_signal_4692) ) ;
    buf_clk new_AGEMA_reg_buffer_3334 ( .C (clk), .D (new_AGEMA_signal_4693), .Q (new_AGEMA_signal_4694) ) ;
    buf_clk new_AGEMA_reg_buffer_3336 ( .C (clk), .D (new_AGEMA_signal_4695), .Q (new_AGEMA_signal_4696) ) ;
    buf_clk new_AGEMA_reg_buffer_3338 ( .C (clk), .D (new_AGEMA_signal_4697), .Q (new_AGEMA_signal_4698) ) ;
    buf_clk new_AGEMA_reg_buffer_3340 ( .C (clk), .D (new_AGEMA_signal_4699), .Q (new_AGEMA_signal_4700) ) ;
    buf_clk new_AGEMA_reg_buffer_3342 ( .C (clk), .D (new_AGEMA_signal_4701), .Q (new_AGEMA_signal_4702) ) ;
    buf_clk new_AGEMA_reg_buffer_3344 ( .C (clk), .D (new_AGEMA_signal_4703), .Q (new_AGEMA_signal_4704) ) ;
    buf_clk new_AGEMA_reg_buffer_3346 ( .C (clk), .D (new_AGEMA_signal_4705), .Q (new_AGEMA_signal_4706) ) ;
    buf_clk new_AGEMA_reg_buffer_3348 ( .C (clk), .D (new_AGEMA_signal_4707), .Q (new_AGEMA_signal_4708) ) ;
    buf_clk new_AGEMA_reg_buffer_3350 ( .C (clk), .D (new_AGEMA_signal_4709), .Q (new_AGEMA_signal_4710) ) ;
    buf_clk new_AGEMA_reg_buffer_3352 ( .C (clk), .D (new_AGEMA_signal_4711), .Q (new_AGEMA_signal_4712) ) ;
    buf_clk new_AGEMA_reg_buffer_3354 ( .C (clk), .D (new_AGEMA_signal_4713), .Q (new_AGEMA_signal_4714) ) ;
    buf_clk new_AGEMA_reg_buffer_3356 ( .C (clk), .D (new_AGEMA_signal_4715), .Q (new_AGEMA_signal_4716) ) ;
    buf_clk new_AGEMA_reg_buffer_3358 ( .C (clk), .D (new_AGEMA_signal_4717), .Q (new_AGEMA_signal_4718) ) ;
    buf_clk new_AGEMA_reg_buffer_3360 ( .C (clk), .D (new_AGEMA_signal_4719), .Q (new_AGEMA_signal_4720) ) ;
    buf_clk new_AGEMA_reg_buffer_3362 ( .C (clk), .D (new_AGEMA_signal_4721), .Q (new_AGEMA_signal_4722) ) ;
    buf_clk new_AGEMA_reg_buffer_3364 ( .C (clk), .D (new_AGEMA_signal_4723), .Q (new_AGEMA_signal_4724) ) ;
    buf_clk new_AGEMA_reg_buffer_3366 ( .C (clk), .D (new_AGEMA_signal_4725), .Q (new_AGEMA_signal_4726) ) ;
    buf_clk new_AGEMA_reg_buffer_3368 ( .C (clk), .D (new_AGEMA_signal_4727), .Q (new_AGEMA_signal_4728) ) ;
    buf_clk new_AGEMA_reg_buffer_3370 ( .C (clk), .D (new_AGEMA_signal_4729), .Q (new_AGEMA_signal_4730) ) ;
    buf_clk new_AGEMA_reg_buffer_3372 ( .C (clk), .D (new_AGEMA_signal_4731), .Q (new_AGEMA_signal_4732) ) ;
    buf_clk new_AGEMA_reg_buffer_3374 ( .C (clk), .D (new_AGEMA_signal_4733), .Q (new_AGEMA_signal_4734) ) ;
    buf_clk new_AGEMA_reg_buffer_3376 ( .C (clk), .D (new_AGEMA_signal_4735), .Q (new_AGEMA_signal_4736) ) ;
    buf_clk new_AGEMA_reg_buffer_3378 ( .C (clk), .D (new_AGEMA_signal_4737), .Q (new_AGEMA_signal_4738) ) ;
    buf_clk new_AGEMA_reg_buffer_3380 ( .C (clk), .D (new_AGEMA_signal_4739), .Q (new_AGEMA_signal_4740) ) ;
    buf_clk new_AGEMA_reg_buffer_3382 ( .C (clk), .D (new_AGEMA_signal_4741), .Q (new_AGEMA_signal_4742) ) ;
    buf_clk new_AGEMA_reg_buffer_3384 ( .C (clk), .D (new_AGEMA_signal_4743), .Q (new_AGEMA_signal_4744) ) ;
    buf_clk new_AGEMA_reg_buffer_3386 ( .C (clk), .D (new_AGEMA_signal_4745), .Q (new_AGEMA_signal_4746) ) ;
    buf_clk new_AGEMA_reg_buffer_3394 ( .C (clk), .D (new_AGEMA_signal_4753), .Q (new_AGEMA_signal_4754) ) ;
    buf_clk new_AGEMA_reg_buffer_3402 ( .C (clk), .D (new_AGEMA_signal_4761), .Q (new_AGEMA_signal_4762) ) ;
    buf_clk new_AGEMA_reg_buffer_3410 ( .C (clk), .D (new_AGEMA_signal_4769), .Q (new_AGEMA_signal_4770) ) ;
    buf_clk new_AGEMA_reg_buffer_3418 ( .C (clk), .D (new_AGEMA_signal_4777), .Q (new_AGEMA_signal_4778) ) ;
    buf_clk new_AGEMA_reg_buffer_3426 ( .C (clk), .D (new_AGEMA_signal_4785), .Q (new_AGEMA_signal_4786) ) ;
    buf_clk new_AGEMA_reg_buffer_3434 ( .C (clk), .D (new_AGEMA_signal_4793), .Q (new_AGEMA_signal_4794) ) ;
    buf_clk new_AGEMA_reg_buffer_3442 ( .C (clk), .D (new_AGEMA_signal_4801), .Q (new_AGEMA_signal_4802) ) ;
    buf_clk new_AGEMA_reg_buffer_3450 ( .C (clk), .D (new_AGEMA_signal_4809), .Q (new_AGEMA_signal_4810) ) ;
    buf_clk new_AGEMA_reg_buffer_3458 ( .C (clk), .D (new_AGEMA_signal_4817), .Q (new_AGEMA_signal_4818) ) ;
    buf_clk new_AGEMA_reg_buffer_3466 ( .C (clk), .D (new_AGEMA_signal_4825), .Q (new_AGEMA_signal_4826) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_63__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4622, new_AGEMA_signal_4620}), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_62__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1905, AddRoundKeyOutput[62]}), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_61__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4626, new_AGEMA_signal_4624}), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_60__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1903, AddRoundKeyOutput[60]}), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_59__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4630, new_AGEMA_signal_4628}), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_58__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1901, AddRoundKeyOutput[58]}), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_57__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4634, new_AGEMA_signal_4632}), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_56__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1899, AddRoundKeyOutput[56]}), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_55__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4638, new_AGEMA_signal_4636}), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_54__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1897, AddRoundKeyOutput[54]}), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_53__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4642, new_AGEMA_signal_4640}), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_52__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1895, AddRoundKeyOutput[52]}), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_51__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4646, new_AGEMA_signal_4644}), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_50__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1893, AddRoundKeyOutput[50]}), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_49__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4650, new_AGEMA_signal_4648}), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_48__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1891, AddRoundKeyOutput[48]}), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_47__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4654, new_AGEMA_signal_4652}), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_46__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1913, AddRoundKeyOutput[46]}), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_45__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4658, new_AGEMA_signal_4656}), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_44__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1911, AddRoundKeyOutput[44]}), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_43__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4662, new_AGEMA_signal_4660}), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_42__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1909, AddRoundKeyOutput[42]}), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_41__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4666, new_AGEMA_signal_4664}), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_40__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1907, AddRoundKeyOutput[40]}), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_39__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4670, new_AGEMA_signal_4668}), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_38__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1921, AddRoundKeyOutput[38]}), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_37__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4674, new_AGEMA_signal_4672}), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_36__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1919, AddRoundKeyOutput[36]}), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_35__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4678, new_AGEMA_signal_4676}), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_34__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1917, AddRoundKeyOutput[34]}), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_33__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4682, new_AGEMA_signal_4680}), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_32__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1915, AddRoundKeyOutput[32]}), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_31__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4686, new_AGEMA_signal_4684}), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_30__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1857, AddRoundKeyOutput[30]}), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_29__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4690, new_AGEMA_signal_4688}), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_28__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1855, AddRoundKeyOutput[28]}), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_27__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4694, new_AGEMA_signal_4692}), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_26__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1853, AddRoundKeyOutput[26]}), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_25__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4698, new_AGEMA_signal_4696}), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_24__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1851, AddRoundKeyOutput[24]}), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_23__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4702, new_AGEMA_signal_4700}), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_22__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1849, AddRoundKeyOutput[22]}), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_21__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4706, new_AGEMA_signal_4704}), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_20__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1847, AddRoundKeyOutput[20]}), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_19__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4710, new_AGEMA_signal_4708}), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_18__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1845, AddRoundKeyOutput[18]}), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_17__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4714, new_AGEMA_signal_4712}), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_16__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1843, AddRoundKeyOutput[16]}), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_15__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4718, new_AGEMA_signal_4716}), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_14__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1841, AddRoundKeyOutput[14]}), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_13__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4722, new_AGEMA_signal_4720}), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_12__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1839, AddRoundKeyOutput[12]}), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_11__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4726, new_AGEMA_signal_4724}), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_10__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1837, AddRoundKeyOutput[10]}), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_9__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4730, new_AGEMA_signal_4728}), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_8__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1835, AddRoundKeyOutput[8]}), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_7__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4734, new_AGEMA_signal_4732}), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_6__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1833, AddRoundKeyOutput[6]}), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_5__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4738, new_AGEMA_signal_4736}), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_4__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1831, AddRoundKeyOutput[4]}), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4742, new_AGEMA_signal_4740}), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1829, AddRoundKeyOutput[2]}), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_4746, new_AGEMA_signal_4744}), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) StateReg_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1827, AddRoundKeyOutput[0]}), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_6__FF_FF ( .CK (clk), .D (new_AGEMA_signal_4754), .Q (FSMReg[6]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_5__FF_FF ( .CK (clk), .D (new_AGEMA_signal_4762), .Q (FSMReg[5]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_4__FF_FF ( .CK (clk), .D (new_AGEMA_signal_4770), .Q (FSMReg[4]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_3__FF_FF ( .CK (clk), .D (new_AGEMA_signal_4778), .Q (FSMReg[3]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_2__FF_FF ( .CK (clk), .D (new_AGEMA_signal_4786), .Q (FSMReg[2]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_4794), .Q (FSMReg[1]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_4802), .Q (FSMReg[0]), .QN () ) ;
    DFF_X1 selectsRegInst_s_current_state_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_4810), .Q (selectsReg[1]), .QN () ) ;
    DFF_X1 selectsRegInst_s_current_state_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_4818), .Q (selectsReg[0]), .QN () ) ;
    DFF_X1 done_reg_FF_FF ( .CK (clk), .D (new_AGEMA_signal_4826), .Q (done), .QN () ) ;
endmodule
